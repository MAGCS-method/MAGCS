module top
#( parameter param538 = {((-{((8'hb3) << (8'hac)), ((8'hbb) && (8'hac))}) ? (7'h42) : (((~(8'ha3)) | {(8'ha2), (8'ha0)}) ? (^~(~(8'hbc))) : ((~^(8'h9d)) ? ((8'hbf) ? (8'ha1) : (8'hac)) : ((8'hb3) ? (8'h9f) : (8'hb4)))))} )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h2c1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire0;
  input wire signed [(5'h11):(1'h0)] wire1;
  input wire [(5'h16):(1'h0)] wire2;
  input wire signed [(4'hc):(1'h0)] wire3;
  input wire [(5'h14):(1'h0)] wire4;
  wire [(2'h2):(1'h0)] wire537;
  wire [(4'hb):(1'h0)] wire536;
  reg signed [(3'h5):(1'h0)] reg535 = (1'h0);
  reg [(4'ha):(1'h0)] reg534 = (1'h0);
  reg [(3'h6):(1'h0)] reg533 = (1'h0);
  reg [(4'h8):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg531 = (1'h0);
  reg [(3'h4):(1'h0)] reg530 = (1'h0);
  reg [(4'ha):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg528 = (1'h0);
  reg [(3'h7):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg525 = (1'h0);
  reg [(5'h11):(1'h0)] reg524 = (1'h0);
  reg [(2'h3):(1'h0)] reg523 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar522 = (1'h0);
  reg [(4'h9):(1'h0)] reg522 = (1'h0);
  reg [(4'hf):(1'h0)] reg521 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg520 = (1'h0);
  reg [(4'ha):(1'h0)] forvar519 = (1'h0);
  wire [(2'h2):(1'h0)] wire518;
  reg signed [(5'h12):(1'h0)] reg517 = (1'h0);
  reg [(4'hc):(1'h0)] reg516 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar514 = (1'h0);
  reg [(3'h6):(1'h0)] reg513 = (1'h0);
  reg [(5'h10):(1'h0)] reg512 = (1'h0);
  reg [(2'h3):(1'h0)] reg511 = (1'h0);
  reg [(5'h16):(1'h0)] forvar510 = (1'h0);
  reg signed [(4'he):(1'h0)] reg509 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire5;
  wire signed [(3'h7):(1'h0)] wire58;
  reg [(4'h8):(1'h0)] forvar60 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar61 = (1'h0);
  reg [(2'h3):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg63 = (1'h0);
  reg [(4'hd):(1'h0)] reg64 = (1'h0);
  reg [(4'hf):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg66 = (1'h0);
  wire [(4'hd):(1'h0)] wire67;
  reg signed [(4'hd):(1'h0)] reg68 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg69 = (1'h0);
  reg [(3'h5):(1'h0)] reg70 = (1'h0);
  reg [(3'h7):(1'h0)] forvar71 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg72 = (1'h0);
  reg [(4'h9):(1'h0)] reg73 = (1'h0);
  reg [(5'h13):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg75 = (1'h0);
  reg signed [(4'he):(1'h0)] reg76 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg77 = (1'h0);
  reg [(3'h4):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar79 = (1'h0);
  reg [(4'ha):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg81 = (1'h0);
  reg [(5'h13):(1'h0)] reg82 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg83 = (1'h0);
  reg [(5'h11):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg85 = (1'h0);
  wire [(4'he):(1'h0)] wire86;
  wire [(4'ha):(1'h0)] wire87;
  wire [(5'h13):(1'h0)] wire88;
  wire [(5'h16):(1'h0)] wire507;
  assign y = {wire537,
                 wire536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 forvar522,
                 reg522,
                 reg521,
                 reg520,
                 forvar519,
                 wire518,
                 reg517,
                 reg516,
                 reg515,
                 forvar514,
                 reg513,
                 reg512,
                 reg511,
                 forvar510,
                 reg509,
                 wire5,
                 wire58,
                 forvar60,
                 forvar61,
                 reg62,
                 reg63,
                 reg64,
                 reg65,
                 reg66,
                 wire67,
                 reg68,
                 reg69,
                 reg70,
                 forvar71,
                 reg72,
                 reg73,
                 reg74,
                 reg75,
                 reg76,
                 reg77,
                 reg78,
                 forvar79,
                 reg80,
                 reg81,
                 reg82,
                 reg83,
                 reg84,
                 reg85,
                 wire86,
                 wire87,
                 wire88,
                 wire507,
                 (1'h0)};
  assign wire5 = {wire2[(5'h14):(5'h13)]};
  module6 modinst59 (.wire9(wire1), .clk(clk), .wire7(wire3), .wire10(wire4), .y(wire58), .wire8(wire2));
  always
    @(posedge clk) begin
      for (forvar60 = (1'h0); (forvar60 < (1'h1)); forvar60 = (forvar60 + (1'h1)))
        begin
          for (forvar61 = (1'h0); (forvar61 < (2'h2)); forvar61 = (forvar61 + (1'h1)))
            begin
              reg62 = ((wire5 ?
                      (($unsigned(forvar61) != wire3[(1'h1):(1'h0)]) ~^ wire58[(1'h1):(1'h0)]) : wire5[(4'h8):(3'h4)]) ?
                  $unsigned({$signed(wire1),
                      $unsigned({wire3, (8'ha2)})}) : wire3);
              reg63 <= (((((forvar61 != (8'hbe)) ?
                      (wire2 ?
                          wire2 : reg62) : reg62[(2'h3):(2'h2)]) << (~|(wire5 ?
                      forvar60 : (8'hb7)))) + (+(&reg62[(2'h3):(1'h1)]))) ?
                  $signed({$unsigned(wire58)}) : (wire1[(4'ha):(4'ha)] ?
                      $signed($signed($unsigned(wire2))) : ($signed((8'ha6)) ?
                          ((wire4 && wire2) ?
                              (forvar60 ?
                                  wire0 : reg62) : (&wire1)) : ($unsigned(wire0) ^~ (+wire1)))));
              reg64 <= ($signed({wire3,
                  reg62}) <<< ($signed((|reg62[(2'h3):(2'h3)])) >>> wire1));
              reg65 <= forvar60[(3'h5):(3'h5)];
            end
        end
      reg66 = $signed((wire1 || wire1[(2'h3):(1'h1)]));
    end
  assign wire67 = wire2;
  always
    @(posedge clk) begin
      reg68 <= wire3[(3'h6):(1'h1)];
      reg69 = reg63;
      reg70 <= $unsigned($unsigned((reg63 >>> $unsigned((wire1 ?
          reg64 : (8'hb5))))));
    end
  always
    @(posedge clk) begin
      for (forvar71 = (1'h0); (forvar71 < (2'h2)); forvar71 = (forvar71 + (1'h1)))
        begin
          if ($unsigned(forvar71))
            begin
              reg72 = ($signed((+{{reg63}})) ?
                  $signed(((&(wire0 ? (8'hac) : (7'h40))) ?
                      reg70[(2'h3):(1'h1)] : ((reg65 <<< reg63) ?
                          (!wire5) : $unsigned(reg62)))) : $unsigned($unsigned((((7'h42) <= reg69) ?
                      (|(8'h9c)) : (~(7'h42))))));
              reg73 = $unsigned((~|$signed(((wire5 ?
                  wire3 : wire3) ^~ (|reg65)))));
              reg74 = {(|wire5[(1'h0):(1'h0)]),
                  ({wire5[(4'h9):(3'h4)],
                      (wire58[(1'h0):(1'h0)] - $signed((8'hb9)))} - reg66)};
              reg75 = {reg70[(1'h1):(1'h1)]};
            end
          else
            begin
              reg72 <= $signed(wire0[(4'ha):(1'h1)]);
            end
          reg76 = $unsigned((reg64[(3'h4):(2'h3)] - reg66[(4'hf):(4'h9)]));
          if ({$unsigned((~|({wire5, reg64} ~^ $unsigned((8'ha1)))))})
            begin
              reg77 = (+forvar61);
              reg78 <= (+(~|(|$unsigned(reg70[(2'h3):(1'h0)]))));
            end
          else
            begin
              reg77 = (8'ha6);
              reg78 = $signed($unsigned(forvar61[(2'h2):(1'h1)]));
            end
          for (forvar79 = (1'h0); (forvar79 < (1'h0)); forvar79 = (forvar79 + (1'h1)))
            begin
              reg80 <= wire0;
              reg81 <= (reg74 != wire67);
              reg82 <= wire0;
              reg83 = reg70;
              reg84 = (wire2[(2'h3):(2'h3)] ?
                  (~(+reg63)) : ((!$signed((reg66 ? forvar79 : reg75))) ?
                      (($signed(reg72) ? $signed(wire2) : reg74) == (wire4 ?
                          (forvar60 + reg81) : wire5[(3'h4):(3'h4)])) : (reg68[(3'h5):(2'h3)] ?
                          reg72 : reg66[(4'h9):(3'h4)])));
            end
          reg85 <= (^~($signed($unsigned(forvar61[(1'h1):(1'h1)])) <<< reg77[(4'h9):(1'h0)]));
        end
    end
  assign wire86 = $unsigned((~&$unsigned(reg73)));
  assign wire87 = (!(~wire1));
  assign wire88 = reg80;
  module89 modinst508 (wire507, clk, reg82, reg77, reg81, wire2, reg74);
  always
    @(posedge clk) begin
      reg509 <= {$unsigned((|((-reg82) ? reg69 : $unsigned(reg83))))};
      for (forvar510 = (1'h0); (forvar510 < (2'h2)); forvar510 = (forvar510 + (1'h1)))
        begin
          reg511 = (reg85[(3'h5):(1'h1)] ? forvar79 : (8'hb6));
          reg512 <= $unsigned((8'hb1));
        end
      reg513 <= (-{$signed((~reg65[(4'hf):(3'h4)]))});
      for (forvar514 = (1'h0); (forvar514 < (2'h3)); forvar514 = (forvar514 + (1'h1)))
        begin
          if ((^$unsigned((~|((reg78 ^~ wire4) + wire0[(4'h8):(3'h7)])))))
            begin
              reg515 = (8'h9d);
              reg516 = ((^~(^~$unsigned((~^reg82)))) <<< $unsigned(reg511[(1'h1):(1'h1)]));
            end
          else
            begin
              reg515 = {(wire5[(4'ha):(2'h3)] || {$signed($unsigned(reg82)),
                      (reg509 + $signed(reg84))})};
              reg516 = reg76;
            end
          reg517 = $signed(reg516);
        end
    end
  assign wire518 = $unsigned($unsigned($signed((|{(8'h9d), wire58}))));
  always
    @(posedge clk) begin
      for (forvar519 = (1'h0); (forvar519 < (3'h4)); forvar519 = (forvar519 + (1'h1)))
        begin
          reg520 <= $unsigned($signed(reg69[(2'h2):(2'h2)]));
        end
      if ((~&(&(((reg66 ? forvar510 : reg66) * (reg512 ?
          reg513 : (7'h41))) * forvar514[(5'h12):(4'ha)]))))
        begin
          if (forvar519)
            begin
              reg521 = (~&reg515[(4'ha):(3'h5)]);
              reg522 <= $unsigned({reg80,
                  {$unsigned($unsigned(reg521)), $signed((reg63 + (7'h46)))}});
            end
          else
            begin
              reg521 <= ($unsigned(((wire518 >>> (+(8'ha4))) ?
                  {$unsigned(reg515),
                      (~wire507)} : {reg73[(2'h2):(2'h2)]})) && (^((reg81 - $unsigned(reg515)) > $unsigned($unsigned((8'ha6))))));
            end
        end
      else
        begin
          reg521 <= (~&reg70[(1'h0):(1'h0)]);
          for (forvar522 = (1'h0); (forvar522 < (2'h3)); forvar522 = (forvar522 + (1'h1)))
            begin
              reg523 = $unsigned($signed((~|reg83)));
              reg524 = {($signed($signed(forvar79[(1'h1):(1'h0)])) << (((~|reg74) ?
                      (^~(7'h41)) : (!reg62)) < $signed($signed(reg76)))),
                  reg66[(3'h4):(3'h4)]};
              reg525 <= reg523[(1'h0):(1'h0)];
              reg526 = ($unsigned((((reg525 <= reg77) ?
                          ((8'had) ? wire3 : (8'ha4)) : (forvar519 ?
                              reg517 : reg517)) ?
                      (!{forvar61}) : forvar71)) ?
                  (wire4 ?
                      (!(~^(forvar60 <= reg82))) : $signed((reg76 ?
                          $unsigned(reg520) : reg76[(4'hd):(4'ha)]))) : ($signed((!(forvar61 <<< wire58))) ?
                      $signed((wire1 ?
                          (reg523 << reg525) : $signed((8'hbe)))) : (^((^forvar79) != $unsigned(reg73)))));
              reg527 = reg525[(5'h12):(4'he)];
            end
          reg528 <= (|$signed((reg83 < $signed(wire0))));
          if ($unsigned((~&((reg517 ?
              (wire518 ? forvar522 : reg527) : (wire86 || forvar60)) | reg81))))
            begin
              reg529 <= {reg516[(4'ha):(1'h0)],
                  (|((reg528 && (7'h45)) ?
                      $unsigned($signed(forvar61)) : $unsigned({reg65})))};
            end
          else
            begin
              reg529 <= $signed($signed(($unsigned((~forvar71)) != ((reg515 ?
                  wire507 : reg68) == (reg62 <= forvar71)))));
              reg530 = reg74;
              reg531 <= (reg526 && (8'hb3));
              reg532 <= $signed(((((^~wire87) ?
                          $unsigned(wire507) : wire1[(4'hf):(4'h8)]) ?
                      reg527 : ($signed(forvar510) ?
                          reg80[(2'h3):(2'h3)] : $unsigned((7'h46)))) ?
                  $signed($signed((~|reg527))) : $signed(reg73[(4'h8):(2'h2)])));
              reg533 = (~$signed($unsigned($signed((|(8'hac))))));
            end
        end
      reg534 = {reg513, $unsigned((-wire87[(4'h8):(3'h6)]))};
      reg535 = ($signed($signed(reg70)) ?
          forvar61 : $signed($unsigned(reg78[(3'h4):(1'h1)])));
    end
  assign wire536 = (^~({(~^{(7'h42), forvar514})} ?
                       ((-$signed(reg532)) ?
                           {{wire87, reg83}} : (((8'hb3) ? wire67 : reg85) ?
                               wire507[(4'ha):(3'h4)] : wire518[(1'h1):(1'h0)])) : (($signed((8'hb4)) & reg84) ?
                           reg535[(2'h3):(1'h1)] : (~^$unsigned(wire1)))));
  assign wire537 = ($signed(($signed(reg534) - {(!reg520),
                       ((8'had) ? reg78 : reg70)})) * forvar510[(4'hc):(4'ha)]);
endmodule

module module89
#( parameter param505 = (^(((^((8'hb1) ? (8'hb5) : (8'hb2))) ? (7'h45) : (((7'h40) ? (8'ha8) : (8'ha6)) <= (^(8'hbd)))) & ((~^((8'hba) != (8'hb8))) ? ((8'ha9) & {(8'hbe)}) : (~^((8'hb0) * (8'hab))))))
, parameter param506 = {((param505 ? {(param505 ^ (8'hab))} : ((param505 ? param505 : param505) ? {param505} : (param505 ? param505 : param505))) + (param505 ? param505 : ((param505 || param505) ? (+param505) : (^param505)))), param505} )
(y, clk, wire90, wire91, wire92, wire93, wire94);
  output wire [(32'h6c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire90;
  input wire [(3'h7):(1'h0)] wire91;
  input wire [(5'h14):(1'h0)] wire92;
  input wire [(5'h16):(1'h0)] wire93;
  input wire [(5'h13):(1'h0)] wire94;
  wire signed [(5'h12):(1'h0)] wire95;
  wire [(3'h6):(1'h0)] wire96;
  wire signed [(5'h15):(1'h0)] wire198;
  wire signed [(5'h16):(1'h0)] wire200;
  reg signed [(5'h13):(1'h0)] reg201 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire202;
  wire [(3'h7):(1'h0)] wire269;
  wire [(4'ha):(1'h0)] wire503;
  assign y = {wire95,
                 wire96,
                 wire198,
                 wire200,
                 reg201,
                 wire202,
                 wire269,
                 wire503,
                 (1'h0)};
  assign wire95 = (^~wire92[(5'h13):(5'h12)]);
  assign wire96 = $signed($unsigned(wire94[(3'h5):(3'h4)]));
  module97 modinst199 (.clk(clk), .wire99(wire90), .wire100(wire93), .wire101(wire91), .y(wire198), .wire98(wire95));
  assign wire200 = {$unsigned((!((wire91 ? (8'hb2) : wire94) > wire94))),
                       $unsigned((((&wire95) ?
                               $unsigned(wire95) : wire90[(3'h4):(2'h3)]) ?
                           ($unsigned(wire93) ^~ $unsigned(wire198)) : wire93[(4'ha):(2'h2)]))};
  always
    @(posedge clk) begin
      reg201 <= (&(8'haf));
    end
  assign wire202 = wire200[(4'hb):(4'hb)];
  module203 modinst270 (wire269, clk, wire95, wire198, wire200, wire94);
  module271 modinst504 (.wire274(wire94), .wire273(wire198), .clk(clk), .wire275(wire202), .wire276(wire90), .wire272(reg201), .y(wire503));
endmodule

module module6
#( parameter param56 = (&(((~|{(8'ha7)}) && (((7'h41) >> (7'h42)) - ((7'h41) == (8'hbc)))) ? ({((8'hab) ~^ (8'hb9)), (-(7'h44))} ? (((8'hbb) ? (7'h42) : (8'h9d)) ^~ ((8'hb9) ? (8'ha2) : (8'ha8))) : (7'h46)) : (((8'hbb) & ((8'hb8) ? (7'h45) : (8'hb8))) ~^ (((8'ha5) ? (8'h9d) : (8'h9e)) - ((7'h41) > (8'h9c))))))
, parameter param57 = param56 )
(y, clk, wire10, wire9, wire8, wire7);
  output wire [(32'h1f9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire10;
  input wire [(2'h2):(1'h0)] wire9;
  input wire signed [(5'h16):(1'h0)] wire8;
  input wire signed [(4'hc):(1'h0)] wire7;
  reg [(4'ha):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg54 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg53 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire52;
  reg signed [(2'h3):(1'h0)] reg51 = (1'h0);
  reg [(2'h2):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg49 = (1'h0);
  reg [(5'h11):(1'h0)] reg48 = (1'h0);
  reg [(5'h11):(1'h0)] forvar47 = (1'h0);
  reg [(3'h7):(1'h0)] reg46 = (1'h0);
  reg [(4'ha):(1'h0)] reg45 = (1'h0);
  reg [(4'hb):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar43 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg40 = (1'h0);
  wire signed [(4'he):(1'h0)] wire39;
  reg [(3'h5):(1'h0)] reg38 = (1'h0);
  reg [(3'h5):(1'h0)] reg37 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg36 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg35 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar34 = (1'h0);
  reg [(2'h3):(1'h0)] reg33 = (1'h0);
  reg [(2'h2):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar31 = (1'h0);
  reg [(4'ha):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar25 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg29 = (1'h0);
  reg [(5'h15):(1'h0)] reg28 = (1'h0);
  reg [(5'h15):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg26 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg25 = (1'h0);
  reg [(3'h4):(1'h0)] reg24 = (1'h0);
  reg [(5'h10):(1'h0)] forvar23 = (1'h0);
  reg [(4'hf):(1'h0)] reg22 = (1'h0);
  reg [(3'h7):(1'h0)] forvar21 = (1'h0);
  reg [(3'h6):(1'h0)] reg20 = (1'h0);
  reg [(5'h10):(1'h0)] reg19 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg18 = (1'h0);
  reg signed [(4'he):(1'h0)] reg17 = (1'h0);
  reg [(4'hd):(1'h0)] reg16 = (1'h0);
  reg signed [(4'he):(1'h0)] reg15 = (1'h0);
  reg [(4'h8):(1'h0)] reg14 = (1'h0);
  reg [(4'ha):(1'h0)] forvar13 = (1'h0);
  reg [(3'h7):(1'h0)] reg12 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg11 = (1'h0);
  assign y = {reg55,
                 reg54,
                 reg53,
                 wire52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 forvar47,
                 reg46,
                 reg45,
                 reg44,
                 forvar43,
                 reg42,
                 reg41,
                 reg40,
                 wire39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 forvar34,
                 reg33,
                 reg32,
                 forvar31,
                 reg30,
                 forvar25,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 forvar23,
                 reg22,
                 forvar21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 forvar13,
                 reg12,
                 reg11,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg11 <= wire10;
      if (wire10)
        begin
          reg12 <= (~|$signed($unsigned(wire7)));
        end
      else
        begin
          reg12 = ($unsigned(reg12[(2'h2):(1'h1)]) ^ wire10);
          for (forvar13 = (1'h0); (forvar13 < (2'h3)); forvar13 = (forvar13 + (1'h1)))
            begin
              reg14 = (wire7[(3'h6):(3'h6)] ?
                  $unsigned($signed(({(8'ha6), reg12} ?
                      $signed(wire10) : (~^wire7)))) : (({$signed(wire8),
                      (forvar13 ? wire8 : wire9)} > ((~&wire7) ?
                      (reg11 | wire9) : forvar13)) && wire9[(2'h2):(1'h0)]));
            end
          reg15 = (((wire8[(4'hd):(2'h2)] <= {$unsigned(forvar13)}) && $unsigned(wire10[(3'h6):(2'h2)])) ?
              wire8 : $unsigned($signed((^~(reg14 > reg11)))));
          reg16 = wire10;
          if (wire8[(5'h14):(2'h3)])
            begin
              reg17 = $unsigned($signed((reg11[(2'h2):(2'h2)] ?
                  reg14 : wire10[(2'h2):(1'h0)])));
              reg18 <= (~^reg12[(1'h1):(1'h1)]);
              reg19 <= (+((~reg14) ?
                  ($signed($unsigned((8'h9d))) != (~|$unsigned(reg17))) : wire10));
              reg20 = (({reg16, (+$signed(reg14))} ?
                      reg18 : $signed(((!forvar13) >> reg12[(3'h5):(1'h1)]))) ?
                  reg14 : ((^~({reg15, reg15} ? (&reg15) : (reg14 + wire9))) ?
                      $signed($unsigned({reg18})) : reg16));
            end
          else
            begin
              reg17 <= forvar13;
              reg18 = (-reg17);
              reg19 <= $signed(reg16[(2'h3):(1'h0)]);
            end
        end
      for (forvar21 = (1'h0); (forvar21 < (3'h4)); forvar21 = (forvar21 + (1'h1)))
        begin
          reg22 = (|(reg11[(4'h8):(2'h3)] ^ reg12));
          for (forvar23 = (1'h0); (forvar23 < (2'h3)); forvar23 = (forvar23 + (1'h1)))
            begin
              reg24 = $unsigned($unsigned(reg17[(3'h5):(1'h0)]));
            end
        end
    end
  always
    @(posedge clk) begin
      if (($unsigned((+((~|reg12) ^~ $unsigned(wire10)))) ?
          (^forvar13[(3'h7):(1'h0)]) : {reg17, (~&{{(8'h9d)}, {reg11}})}))
        begin
          if (reg12)
            begin
              reg25 <= reg17[(4'hc):(2'h3)];
              reg26 = ((~|$signed(reg11[(4'hf):(4'hf)])) ?
                  ((~&(-forvar23[(4'h9):(4'h8)])) ?
                      (((reg11 >= reg20) ?
                              ((8'haa) ~^ reg20) : $signed(reg17)) ?
                          (-$unsigned(wire9)) : (^$signed(reg18))) : $signed(((|forvar23) ?
                          $unsigned(reg20) : (8'hbb)))) : {$unsigned($signed(reg16[(4'hb):(4'hb)]))});
              reg27 = (^$signed((((7'h41) > reg11[(3'h5):(3'h5)]) ~^ ((&wire8) ?
                  reg12[(2'h3):(2'h3)] : (8'ha8)))));
            end
          else
            begin
              reg25 <= ($signed({$signed((reg19 > wire7)),
                      ((reg12 && (8'hac)) > {reg17, wire9})}) ?
                  (^reg14) : $signed(($signed($signed(wire8)) ?
                      forvar23[(4'hc):(3'h4)] : (((8'hbb) ?
                          forvar21 : reg17) || $unsigned(forvar21)))));
              reg26 = (^~($signed(wire9[(2'h2):(2'h2)]) ?
                  $signed(reg19) : reg17[(4'ha):(3'h4)]));
              reg27 = (+wire8[(4'hf):(1'h0)]);
              reg28 = $unsigned((((^((8'hb6) ?
                  reg17 : reg11)) >>> $unsigned((-reg17))) ~^ reg12[(3'h7):(3'h7)]));
              reg29 <= $unsigned(reg12[(2'h2):(2'h2)]);
            end
        end
      else
        begin
          for (forvar25 = (1'h0); (forvar25 < (2'h2)); forvar25 = (forvar25 + (1'h1)))
            begin
              reg26 = (^wire9);
            end
          if ($unsigned({forvar21[(2'h2):(1'h1)],
              (reg25 ?
                  (reg25[(3'h4):(1'h1)] ~^ reg26[(3'h6):(2'h3)]) : $signed(reg29))}))
            begin
              reg27 = ($signed({((8'hbd) ? reg16 : (^reg18))}) ?
                  ($signed(($signed(reg28) ?
                      $signed(reg17) : (+reg19))) >= (reg17[(1'h1):(1'h0)] && (&$unsigned(forvar13)))) : ((wire10[(3'h5):(1'h1)] ?
                          $unsigned($signed((8'ha9))) : $unsigned((+(8'ha5)))) ?
                      reg26 : ($unsigned($signed(reg22)) + {(forvar23 - reg22)})));
              reg28 <= reg20;
              reg29 = (~^(!reg29[(1'h0):(1'h0)]));
              reg30 <= ((+{forvar13}) ?
                  (^~((8'hb2) ?
                      ((reg28 ?
                          (8'hb0) : wire7) && reg22) : reg14)) : $unsigned(forvar23[(4'he):(1'h0)]));
            end
          else
            begin
              reg27 <= $unsigned($unsigned(((&{reg18}) ^~ $unsigned((reg26 ?
                  reg11 : (8'had))))));
              reg28 = {$signed((forvar21 + (reg25 & {reg30}))),
                  $signed(((^(8'ha4)) ? forvar21[(2'h2):(1'h0)] : (!reg30)))};
              reg29 = (&(reg24 <<< ((wire8 <= reg12) ^~ ((forvar21 || wire10) ?
                  (|reg30) : reg24[(2'h3):(1'h1)]))));
              reg30 = $unsigned(reg12[(3'h7):(2'h2)]);
            end
        end
      for (forvar31 = (1'h0); (forvar31 < (2'h3)); forvar31 = (forvar31 + (1'h1)))
        begin
          reg32 <= $unsigned(($signed($signed((reg14 || wire7))) * reg24));
          reg33 = ((reg17 ?
              $unsigned(reg22[(1'h0):(1'h0)]) : reg27) >= $unsigned((!$signed(reg18))));
          for (forvar34 = (1'h0); (forvar34 < (1'h0)); forvar34 = (forvar34 + (1'h1)))
            begin
              reg35 <= reg26;
            end
        end
      reg36 <= $unsigned(wire8[(3'h5):(1'h0)]);
      reg37 <= {(reg11[(3'h6):(3'h5)] && reg29[(3'h6):(1'h1)]),
          ($signed($unsigned((reg29 ? wire10 : reg36))) + (8'hb4))};
      reg38 <= (wire7[(4'h8):(3'h4)] < (reg32[(1'h1):(1'h1)] ?
          ($unsigned(reg24[(2'h2):(1'h0)]) - forvar34[(2'h3):(1'h0)]) : $unsigned(forvar21)));
    end
  assign wire39 = (~&reg18[(4'ha):(1'h1)]);
  always
    @(posedge clk) begin
      reg40 <= wire9[(2'h2):(1'h1)];
      reg41 = ((($signed(reg20[(1'h0):(1'h0)]) || $signed($signed(reg12))) ?
              $unsigned(reg15) : ((&forvar21[(3'h5):(3'h4)]) || (~{(7'h40)}))) ?
          {reg33[(2'h3):(2'h2)],
              ($unsigned((-reg37)) ?
                  (reg40[(1'h0):(1'h0)] ?
                      {reg38,
                          reg16} : $unsigned(forvar25)) : (~&reg24[(1'h0):(1'h0)]))} : (((reg17[(4'ha):(3'h5)] && {forvar23}) ?
                  wire7 : reg22) ?
              (reg28[(3'h4):(3'h4)] ?
                  ((wire7 ? reg14 : reg15) ?
                      (reg35 ?
                          forvar21 : (8'hbf)) : (&reg22)) : $signed($unsigned(wire9))) : $signed(((reg32 & (8'hb8)) <= ((8'ha7) ?
                  wire7 : reg24)))));
      reg42 = (&{$signed($signed(reg11))});
      for (forvar43 = (1'h0); (forvar43 < (3'h4)); forvar43 = (forvar43 + (1'h1)))
        begin
          reg44 = $signed({(|(+$signed(forvar43))), (~^(+(reg25 >= reg33)))});
          reg45 = reg30;
          reg46 = ((reg19[(4'h9):(2'h3)] | ($signed($unsigned(reg40)) == $signed(reg45[(3'h7):(3'h7)]))) ?
              (~(-((reg45 & forvar43) > {(8'haf)}))) : ($unsigned(forvar25) ?
                  reg32 : $signed(((reg38 < reg16) - $unsigned(reg37)))));
          for (forvar47 = (1'h0); (forvar47 < (1'h0)); forvar47 = (forvar47 + (1'h1)))
            begin
              reg48 = ($signed($unsigned(wire8)) ? forvar47 : reg45);
              reg49 <= ((~^((wire9 ?
                          (reg25 << (8'h9e)) : wire10[(3'h5):(2'h2)]) ?
                      ((forvar13 ? reg40 : reg32) ?
                          $unsigned(reg30) : $signed(reg37)) : $signed((reg36 & reg11)))) ?
                  ({(~|(reg36 | reg41)),
                      (~&wire39[(4'he):(2'h2)])} && (+reg11[(4'he):(1'h1)])) : {reg46,
                      $unsigned(reg45[(2'h2):(1'h1)])});
              reg50 = (^$unsigned($unsigned((^(reg45 ? forvar34 : reg19)))));
              reg51 = $unsigned((-reg41));
            end
        end
    end
  assign wire52 = (8'hbc);
  always
    @(posedge clk) begin
      reg53 <= ($unsigned({(-reg37)}) ?
          $signed($unsigned(forvar47[(3'h7):(3'h5)])) : $signed(reg11[(4'hb):(4'hb)]));
      reg54 <= reg36;
      reg55 <= (+reg19);
    end
endmodule

module module271
#( parameter param502 = ((((+((8'haf) ^ (8'hb9))) - (|((8'ha6) ? (8'hb3) : (8'h9c)))) && {({(8'h9e)} & {(8'ha4), (8'haf)}), (~{(8'h9c)})}) ? (((^(-(7'h41))) - (((8'hbf) >>> (8'h9f)) ? (-(8'hac)) : ((8'ha2) ? (8'hb6) : (8'ha2)))) - (^(((8'h9e) ? (7'h45) : (8'hb6)) ? (+(7'h43)) : ((8'hbb) - (8'hb0))))) : ({((8'h9f) ? ((8'hbb) ? (8'ha1) : (8'h9e)) : (~^(8'ha7))), (((8'hbe) ? (7'h43) : (8'hb3)) ? {(8'ha6), (8'hb3)} : {(7'h45), (8'hbc)})} ? ({(+(8'hbd))} ? (((8'h9d) ? (8'hbd) : (7'h43)) || ((8'hb1) ? (8'hba) : (7'h44))) : (!((8'hb9) ? (8'hb8) : (8'hbc)))) : ((((8'hb0) ? (8'ha6) : (8'ha3)) ? ((8'haa) ^ (8'hb1)) : (^(8'hba))) != ((+(8'hb3)) ? {(8'ha6), (7'h44)} : ((7'h45) ? (8'haa) : (8'haf)))))) )
(y, clk, wire276, wire275, wire274, wire273, wire272);
  output wire [(32'h2ea):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire276;
  input wire [(3'h4):(1'h0)] wire275;
  input wire signed [(5'h13):(1'h0)] wire274;
  input wire signed [(5'h15):(1'h0)] wire273;
  input wire signed [(3'h7):(1'h0)] wire272;
  wire signed [(3'h7):(1'h0)] wire501;
  wire [(5'h13):(1'h0)] wire500;
  reg [(5'h11):(1'h0)] reg499 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg498 = (1'h0);
  reg [(4'hf):(1'h0)] reg489 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg497 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg496 = (1'h0);
  reg [(5'h14):(1'h0)] reg495 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg494 = (1'h0);
  reg [(4'hd):(1'h0)] reg493 = (1'h0);
  reg [(4'hd):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg491 = (1'h0);
  reg [(4'h9):(1'h0)] reg490 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar489 = (1'h0);
  reg [(4'he):(1'h0)] reg488 = (1'h0);
  reg [(2'h3):(1'h0)] reg487 = (1'h0);
  reg [(5'h12):(1'h0)] reg486 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg485 = (1'h0);
  wire [(3'h4):(1'h0)] wire484;
  wire signed [(4'h9):(1'h0)] wire483;
  wire [(5'h13):(1'h0)] wire482;
  reg signed [(3'h4):(1'h0)] reg481 = (1'h0);
  wire [(4'h9):(1'h0)] wire480;
  wire [(4'h8):(1'h0)] wire479;
  wire [(5'h16):(1'h0)] wire478;
  wire signed [(4'hd):(1'h0)] wire477;
  wire signed [(5'h11):(1'h0)] wire476;
  wire [(3'h4):(1'h0)] wire475;
  reg signed [(4'he):(1'h0)] reg474 = (1'h0);
  reg [(4'he):(1'h0)] reg473 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg472 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg471 = (1'h0);
  reg [(4'h9):(1'h0)] reg470 = (1'h0);
  reg [(5'h15):(1'h0)] reg469 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg468 = (1'h0);
  reg [(2'h2):(1'h0)] reg467 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg466 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg465 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg464 = (1'h0);
  reg [(4'ha):(1'h0)] reg463 = (1'h0);
  reg [(2'h3):(1'h0)] forvar462 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg461 = (1'h0);
  reg [(4'he):(1'h0)] reg460 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg459 = (1'h0);
  reg [(5'h16):(1'h0)] reg458 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg457 = (1'h0);
  reg [(4'hd):(1'h0)] reg456 = (1'h0);
  reg [(5'h13):(1'h0)] forvar455 = (1'h0);
  reg [(3'h6):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg453 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar452 = (1'h0);
  reg [(3'h6):(1'h0)] reg451 = (1'h0);
  reg [(5'h16):(1'h0)] reg450 = (1'h0);
  reg [(5'h10):(1'h0)] reg449 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar448 = (1'h0);
  reg [(5'h15):(1'h0)] reg447 = (1'h0);
  reg [(4'he):(1'h0)] forvar446 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire445;
  wire signed [(2'h2):(1'h0)] wire443;
  wire signed [(4'hc):(1'h0)] wire277;
  assign y = {wire501,
                 wire500,
                 reg499,
                 reg498,
                 reg489,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 forvar489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 wire484,
                 wire483,
                 wire482,
                 reg481,
                 wire480,
                 wire479,
                 wire478,
                 wire477,
                 wire476,
                 wire475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 forvar462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 forvar455,
                 reg454,
                 reg453,
                 forvar452,
                 reg451,
                 reg450,
                 reg449,
                 forvar448,
                 reg447,
                 forvar446,
                 wire445,
                 wire443,
                 wire277,
                 (1'h0)};
  assign wire277 = {((-$unsigned((+wire275))) > $signed((wire275[(2'h2):(1'h0)] ?
                           $signed(wire276) : (wire272 >= wire275)))),
                       wire274[(3'h7):(1'h1)]};
  module278 modinst444 (wire443, clk, wire276, wire272, wire274, wire277);
  assign wire445 = {wire274};
  always
    @(posedge clk) begin
      for (forvar446 = (1'h0); (forvar446 < (1'h1)); forvar446 = (forvar446 + (1'h1)))
        begin
          reg447 <= ((~$unsigned(forvar446)) < (wire272 ~^ wire276[(4'h8):(1'h0)]));
          for (forvar448 = (1'h0); (forvar448 < (3'h4)); forvar448 = (forvar448 + (1'h1)))
            begin
              reg449 <= (+wire445);
            end
          reg450 = reg449;
          reg451 <= ({forvar448,
              ((forvar448 ?
                      reg449[(4'hf):(3'h6)] : (wire277 ? (8'ha5) : reg447)) ?
                  wire277[(4'ha):(3'h7)] : $unsigned((~&wire277)))} >>> reg449[(4'ha):(3'h5)]);
        end
      for (forvar452 = (1'h0); (forvar452 < (1'h1)); forvar452 = (forvar452 + (1'h1)))
        begin
          reg453 <= wire274[(5'h13):(3'h6)];
          reg454 = wire445;
          for (forvar455 = (1'h0); (forvar455 < (2'h2)); forvar455 = (forvar455 + (1'h1)))
            begin
              reg456 <= $signed((!(+((wire273 >> wire274) * (wire277 ?
                  reg450 : reg450)))));
              reg457 <= ((^$signed($signed($unsigned((7'h44))))) ?
                  ($signed((^$unsigned(reg454))) > $signed({wire445[(1'h1):(1'h0)]})) : reg453);
              reg458 <= wire277;
            end
        end
      reg459 = reg457;
      reg460 = wire274[(1'h0):(1'h0)];
      reg461 = {wire443[(2'h2):(2'h2)]};
    end
  always
    @(posedge clk) begin
      for (forvar462 = (1'h0); (forvar462 < (2'h2)); forvar462 = (forvar462 + (1'h1)))
        begin
          reg463 = reg454[(1'h0):(1'h0)];
          reg464 <= wire445[(2'h2):(2'h2)];
          if ({{forvar446}})
            begin
              reg465 <= ((-$unsigned((+(~|reg457)))) & (reg454 > ($unsigned((-forvar446)) ~^ reg454[(2'h3):(1'h0)])));
              reg466 <= (^~wire275);
              reg467 = forvar462;
              reg468 <= forvar452;
              reg469 <= {$unsigned((reg460[(2'h3):(2'h2)] ?
                      $unsigned($unsigned(forvar455)) : $unsigned((~&reg464))))};
            end
          else
            begin
              reg465 = (|$signed((((reg456 ? reg459 : forvar448) ?
                  forvar446[(3'h4):(2'h2)] : (reg451 && reg450)) >= (reg449[(2'h3):(1'h0)] ?
                  wire273[(2'h2):(2'h2)] : (forvar452 >= reg461)))));
            end
          if (forvar452)
            begin
              reg470 <= (reg457[(2'h2):(1'h1)] ?
                  ({((~forvar452) >= $signed((8'h9f))),
                      reg465} > $signed(($unsigned(wire443) ?
                      $unsigned(forvar448) : reg454[(2'h2):(1'h0)]))) : $signed((^((reg459 + reg464) ^~ (8'ha3)))));
              reg471 <= ((wire275[(1'h1):(1'h1)] | (^$signed($unsigned((8'hac))))) ?
                  {(reg449 ?
                          $unsigned(reg460[(4'hc):(4'ha)]) : reg464[(5'h15):(4'hd)]),
                      $unsigned(reg451)} : ((($signed((7'h42)) >= forvar446) ?
                      $signed((^~(8'ha5))) : $signed($signed(reg463))) + (wire277[(4'hb):(4'h9)] >= reg447)));
            end
          else
            begin
              reg470 = wire276[(3'h5):(1'h0)];
              reg471 <= wire272;
              reg472 = reg447[(5'h15):(4'h8)];
              reg473 = reg472[(5'h10):(4'hd)];
              reg474 <= forvar462[(1'h1):(1'h0)];
            end
        end
    end
  assign wire475 = (8'hb2);
  assign wire476 = {$signed($signed((reg466[(3'h4):(2'h2)] > reg453))),
                       (reg450 ?
                           ({$unsigned((7'h43)), (wire276 < wire272)} ?
                               {$signed(reg461)} : reg463[(4'ha):(4'h9)]) : forvar448)};
  assign wire477 = wire274;
  assign wire478 = $signed(($unsigned(wire477[(4'h8):(3'h6)]) >= $unsigned($signed((reg449 >>> reg466)))));
  assign wire479 = ((($signed($signed(reg466)) != {(!reg469),
                       $unsigned(reg449)}) << wire274[(4'h8):(3'h4)]) <<< $signed((&wire445)));
  assign wire480 = {wire273[(1'h1):(1'h0)], reg460};
  always
    @(posedge clk) begin
      reg481 = $unsigned($signed(wire479));
    end
  assign wire482 = (((~wire479[(2'h2):(1'h1)]) ?
                           $signed({$signed((8'h9f))}) : reg474) ?
                       wire277[(1'h0):(1'h0)] : {reg447, (&$unsigned(reg466))});
  assign wire483 = (($signed(reg465[(3'h5):(1'h0)]) && wire477) ~^ ((&(^(~&forvar452))) ?
                       (-(~&wire478[(4'he):(2'h2)])) : reg472));
  assign wire484 = ((forvar455 ^~ ({{wire475, (8'had)}} ?
                       $unsigned((|forvar448)) : $signed(forvar455[(3'h5):(1'h1)]))) ~^ $signed($signed(wire272)));
  always
    @(posedge clk) begin
      if ($unsigned({{$unsigned(((8'haf) < reg453)), reg467}}))
        begin
          if (($unsigned($unsigned(($unsigned((7'h43)) ?
              $signed((8'hb0)) : $signed(forvar448)))) + ($unsigned($signed((reg465 >>> wire443))) ?
              wire277[(4'h9):(3'h4)] : (~|$signed(forvar448[(4'hf):(3'h5)])))))
            begin
              reg485 = reg470[(2'h3):(1'h0)];
              reg486 = (~&$signed((reg450 >= ((reg485 | wire476) & (reg468 >= reg474)))));
              reg487 <= (wire272[(1'h1):(1'h0)] ~^ ((|$unsigned((reg450 ?
                  reg449 : forvar455))) + (wire484[(2'h2):(1'h1)] ?
                  (wire478[(4'h9):(3'h4)] ?
                      (wire274 <= reg464) : $unsigned(reg456)) : ($unsigned(wire443) ?
                      reg463[(1'h0):(1'h0)] : (wire273 ? reg468 : wire277)))));
              reg488 <= (($signed((~(wire276 <= wire477))) ^~ (^~$signed((wire478 ^ wire476)))) ?
                  forvar455 : (^~(|((8'hb6) > $signed(reg472)))));
            end
          else
            begin
              reg485 = $signed(forvar446);
            end
          for (forvar489 = (1'h0); (forvar489 < (2'h2)); forvar489 = (forvar489 + (1'h1)))
            begin
              reg490 <= ({$unsigned($signed((!forvar452))), $signed(reg456)} ?
                  (|(|((wire475 ? reg473 : wire482) ?
                      (8'hb0) : $unsigned(reg488)))) : $signed($signed(reg473)));
              reg491 <= (reg460 ?
                  wire479[(4'h8):(3'h7)] : wire479[(3'h4):(1'h1)]);
              reg492 <= $signed(($signed($unsigned((~^reg471))) ?
                  forvar462 : $signed(reg459)));
              reg493 <= {wire275[(2'h3):(2'h3)],
                  ($unsigned(wire274[(3'h5):(3'h4)]) <<< reg461[(5'h13):(4'hc)])};
              reg494 = $signed(wire479[(4'h8):(3'h6)]);
            end
          if (reg470)
            begin
              reg495 = (!reg469[(5'h14):(1'h0)]);
            end
          else
            begin
              reg495 = forvar455[(3'h7):(2'h2)];
            end
          reg496 <= wire272[(3'h6):(1'h1)];
          reg497 <= (|{forvar455[(3'h4):(3'h4)],
              (forvar489[(3'h4):(3'h4)] ?
                  ((reg481 ? wire475 : (8'h9e)) ?
                      reg487[(1'h0):(1'h0)] : ((8'ha1) && reg459)) : $unsigned($unsigned((8'hb5))))});
        end
      else
        begin
          reg485 <= ($signed((wire276 ^~ (((8'ha1) + wire277) * forvar446))) ^ $signed(reg457[(1'h0):(1'h0)]));
          if (reg463)
            begin
              reg486 = (+$signed(wire273[(5'h15):(2'h2)]));
              reg487 = $unsigned(wire274);
              reg488 = $unsigned($signed((wire443[(1'h0):(1'h0)] ?
                  reg470 : ((&forvar452) ?
                      (+(8'ha9)) : reg468[(1'h1):(1'h1)]))));
            end
          else
            begin
              reg486 = forvar448;
              reg487 <= $signed(wire483[(4'h8):(3'h6)]);
              reg488 = reg454;
            end
          if ((wire475 + {((|(wire484 ?
                  reg497 : wire445)) <<< $signed($unsigned(wire277))),
              {$signed($signed(reg486))}}))
            begin
              reg489 = (|$unsigned($unsigned(($unsigned(forvar452) ?
                  (reg472 ? reg453 : (7'h40)) : $unsigned(reg456)))));
            end
          else
            begin
              reg489 = (reg496 || {$signed((reg463 == $signed(reg491)))});
            end
          reg490 <= {{reg463[(4'h9):(3'h7)]}};
        end
      reg498 = (reg490[(1'h1):(1'h0)] != wire477);
      reg499 <= reg449[(4'hc):(1'h1)];
    end
  assign wire500 = (&($unsigned(reg493) ?
                       ($unsigned((reg486 ? reg449 : wire476)) ?
                           (((8'ha9) == reg473) > wire480) : (-$signed(reg495))) : (wire476[(4'hc):(4'h9)] ?
                           reg453 : reg447[(3'h5):(2'h3)])));
  assign wire501 = reg465;
endmodule

module module203
#( parameter param267 = (~&({((8'hb4) + ((8'h9d) != (8'hb3))), (((8'h9e) ? (8'hac) : (8'hac)) & (~(8'hb0)))} ? ((((8'ha3) - (8'hbd)) ? ((8'h9e) ? (7'h46) : (7'h43)) : (7'h40)) >= {((8'h9c) & (8'ha5)), ((7'h45) ? (8'hbe) : (7'h41))}) : (({(7'h43), (8'ha3)} > ((8'had) ? (7'h40) : (7'h42))) ? (((8'hb2) ? (8'h9d) : (8'hb5)) ? ((8'hb2) + (8'hb8)) : ((8'had) != (8'ha6))) : ((-(8'hb8)) ? (~&(8'h9e)) : ((7'h41) <= (8'ha4))))))
, parameter param268 = (((+param267) ? (param267 == (+{param267})) : ({(~|param267), {(8'hbc)}} && {((7'h42) ? (8'hb7) : param267)})) ^~ param267) )
(y, clk, wire207, wire206, wire205, wire204);
  output wire [(32'h304):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire207;
  input wire signed [(4'h8):(1'h0)] wire206;
  input wire [(5'h16):(1'h0)] wire205;
  input wire signed [(3'h5):(1'h0)] wire204;
  wire [(5'h12):(1'h0)] wire266;
  reg signed [(5'h14):(1'h0)] reg265 = (1'h0);
  reg [(4'ha):(1'h0)] reg264 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg260 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar259 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg263 = (1'h0);
  reg [(5'h14):(1'h0)] reg262 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg261 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar260 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg259 = (1'h0);
  reg [(4'hb):(1'h0)] reg258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg257 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg256 = (1'h0);
  reg [(5'h13):(1'h0)] reg255 = (1'h0);
  reg [(4'hd):(1'h0)] reg254 = (1'h0);
  reg [(5'h13):(1'h0)] forvar253 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg251 = (1'h0);
  reg [(4'hc):(1'h0)] reg250 = (1'h0);
  reg [(5'h12):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg248 = (1'h0);
  reg [(4'hc):(1'h0)] reg247 = (1'h0);
  reg [(3'h5):(1'h0)] forvar246 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar245 = (1'h0);
  reg [(2'h2):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg243 = (1'h0);
  reg signed [(4'he):(1'h0)] reg242 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg241 = (1'h0);
  reg [(5'h12):(1'h0)] forvar240 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg239 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg237 = (1'h0);
  reg [(5'h11):(1'h0)] forvar236 = (1'h0);
  reg [(5'h12):(1'h0)] forvar235 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg234 = (1'h0);
  wire [(5'h11):(1'h0)] wire233;
  wire signed [(4'he):(1'h0)] wire232;
  wire signed [(2'h2):(1'h0)] wire231;
  reg [(3'h6):(1'h0)] reg230 = (1'h0);
  reg [(4'h9):(1'h0)] reg229 = (1'h0);
  reg [(4'hd):(1'h0)] reg228 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg227 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg226 = (1'h0);
  reg [(4'h8):(1'h0)] forvar225 = (1'h0);
  reg [(5'h13):(1'h0)] forvar224 = (1'h0);
  reg [(3'h5):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg223 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg222 = (1'h0);
  reg [(4'hb):(1'h0)] reg221 = (1'h0);
  reg [(4'hc):(1'h0)] reg220 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg219 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar218 = (1'h0);
  reg [(3'h4):(1'h0)] reg217 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg216 = (1'h0);
  reg [(5'h13):(1'h0)] reg215 = (1'h0);
  reg [(3'h4):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg212 = (1'h0);
  reg [(5'h11):(1'h0)] reg211 = (1'h0);
  wire [(5'h11):(1'h0)] wire210;
  wire [(5'h12):(1'h0)] wire209;
  wire signed [(4'hc):(1'h0)] wire208;
  assign y = {wire266,
                 reg265,
                 reg264,
                 reg260,
                 forvar259,
                 reg263,
                 reg262,
                 reg261,
                 forvar260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 forvar253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 forvar246,
                 forvar245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 forvar240,
                 reg239,
                 reg238,
                 reg237,
                 forvar236,
                 forvar235,
                 reg234,
                 wire233,
                 wire232,
                 wire231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 forvar225,
                 forvar224,
                 reg218,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 forvar218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 wire210,
                 wire209,
                 wire208,
                 (1'h0)};
  assign wire208 = ({$unsigned($unsigned(wire204)), {wire204[(3'h5):(1'h0)]}} ?
                       $unsigned($signed((wire205 - wire206))) : ((8'h9f) ?
                           (($unsigned(wire207) << {wire204}) || wire206[(2'h3):(1'h1)]) : (~&$unsigned((wire206 ?
                               (8'hae) : wire204)))));
  assign wire209 = wire206;
  assign wire210 = (8'hbf);
  always
    @(posedge clk) begin
      if ((-((((^~wire207) - (+wire204)) != $unsigned(wire207)) >>> ((^wire209) ?
          (~wire210[(4'hd):(2'h2)]) : wire209[(4'hd):(2'h3)]))))
        begin
          reg211 = ((8'ha2) ?
              {(^$signed(wire204)),
                  ($unsigned(wire209) ~^ wire204)} : $unsigned((8'hb0)));
          if (($signed((~wire209[(5'h11):(3'h4)])) ?
              ($signed(((&wire205) ? wire206[(4'h8):(1'h0)] : wire204)) ?
                  ((&reg211[(4'hf):(3'h5)]) ?
                      ((wire209 >> wire208) ?
                          $unsigned(wire205) : wire208) : (wire204 & wire206[(3'h6):(3'h6)])) : (&((!wire207) >>> {reg211}))) : (wire210[(3'h7):(3'h7)] ?
                  reg211 : wire210[(3'h6):(2'h3)])))
            begin
              reg212 <= (~wire206[(1'h0):(1'h0)]);
              reg213 <= (((!reg211[(4'hc):(1'h0)]) ?
                      ((~&wire210[(1'h0):(1'h0)]) << $unsigned(wire208)) : (-{(+wire204),
                          (wire209 ? wire207 : wire208)})) ?
                  $unsigned($signed(((wire204 ? reg212 : wire204) - (reg212 ?
                      reg212 : reg212)))) : ((|wire208) - wire207));
              reg214 = ($signed((($signed(wire209) ?
                      (+reg212) : (wire205 ? wire206 : (8'hbc))) ?
                  (wire207 ?
                      (wire204 ?
                          reg212 : (8'hb8)) : (8'ha1)) : $signed((reg211 ?
                      wire206 : reg212)))) < ($unsigned($signed(wire206)) <<< $signed(wire205[(1'h0):(1'h0)])));
              reg215 = $signed(((~|(reg212[(4'hd):(4'h8)] ^~ (reg213 & wire210))) ?
                  (~&wire206[(3'h6):(3'h6)]) : wire205));
            end
          else
            begin
              reg212 <= (~(-wire204[(2'h3):(2'h2)]));
              reg213 = $signed(wire210);
              reg214 = wire207[(3'h5):(2'h3)];
              reg215 = reg213[(3'h4):(1'h0)];
            end
        end
      else
        begin
          if (((wire209 ?
                  ({$unsigned(wire206)} << $unsigned($signed(reg212))) : wire207[(4'hd):(2'h3)]) ?
              (wire205[(3'h5):(2'h2)] ?
                  (8'hbd) : {wire210[(3'h7):(3'h6)]}) : (wire208[(3'h5):(2'h2)] ?
                  wire209 : (reg211[(3'h5):(3'h4)] ? reg214 : (~|wire208)))))
            begin
              reg211 = reg213;
              reg212 <= (reg212[(3'h4):(1'h0)] + $signed((!reg215[(2'h2):(1'h1)])));
              reg213 <= $unsigned((8'hae));
              reg214 = reg213;
            end
          else
            begin
              reg211 <= reg213[(4'hf):(4'h9)];
            end
          reg215 = (|reg214[(2'h3):(2'h2)]);
        end
      if ((8'hbe))
        begin
          reg216 <= $unsigned({wire204[(3'h4):(2'h3)], reg213});
          reg217 <= $signed({((reg211[(4'hb):(4'ha)] << reg216[(3'h7):(3'h5)]) && $signed(wire209[(4'hb):(3'h6)]))});
          for (forvar218 = (1'h0); (forvar218 < (1'h0)); forvar218 = (forvar218 + (1'h1)))
            begin
              reg219 <= (({$unsigned((+wire209)),
                          ((wire205 - reg211) ?
                              $unsigned(wire206) : reg214[(3'h4):(2'h2)])} ?
                      ($unsigned($unsigned(reg217)) <= reg214[(1'h0):(1'h0)]) : $signed((((7'h45) ?
                              reg211 : wire204) ?
                          wire204 : wire207[(4'hd):(3'h7)]))) ?
                  (~|reg213[(3'h7):(1'h0)]) : ($unsigned((reg215[(4'ha):(2'h2)] != (forvar218 || reg214))) && {$unsigned({reg212,
                          (8'hbd)}),
                      reg214[(1'h1):(1'h0)]}));
              reg220 <= reg215[(5'h10):(4'hf)];
              reg221 = reg214[(1'h0):(1'h0)];
              reg222 <= {((wire210 ?
                      ($signed(wire208) * wire210[(3'h6):(3'h5)]) : {(~reg217),
                          (reg221 ?
                              wire204 : wire210)}) ~^ $signed($unsigned((wire206 <= forvar218)))),
                  (reg217[(1'h1):(1'h0)] ?
                      (!$signed(reg216)) : wire209[(2'h3):(1'h0)])};
              reg223 <= reg212;
            end
        end
      else
        begin
          reg216 <= reg214[(2'h3):(1'h1)];
          reg217 = $signed((^~{reg215}));
          reg218 = ($unsigned($unsigned({(wire205 ? reg222 : reg215)})) ?
              (~^wire206[(3'h5):(1'h1)]) : ({wire209[(1'h0):(1'h0)]} ?
                  (~&{$unsigned(reg222)}) : (!(8'hb3))));
        end
      for (forvar224 = (1'h0); (forvar224 < (2'h2)); forvar224 = (forvar224 + (1'h1)))
        begin
          for (forvar225 = (1'h0); (forvar225 < (2'h3)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 <= (-reg213);
              reg227 = (($signed(reg216) << (reg222[(3'h7):(2'h2)] ?
                  wire205 : ($unsigned(wire210) ?
                      wire210 : (|reg211)))) < (~&$signed(reg213)));
              reg228 <= reg213[(3'h5):(2'h2)];
              reg229 <= $signed((8'ha0));
              reg230 = $signed((reg226 ~^ ($signed(reg223) >= $signed((reg217 ^~ wire209)))));
            end
        end
    end
  assign wire231 = reg212[(4'hd):(4'ha)];
  assign wire232 = reg214[(1'h1):(1'h1)];
  assign wire233 = (^((forvar225[(3'h4):(3'h4)] ?
                           $signed(reg227[(4'hc):(3'h5)]) : (^$signed(reg218))) ?
                       wire231[(1'h1):(1'h0)] : reg220[(4'hc):(4'h9)]));
  always
    @(posedge clk) begin
      reg234 <= (-$unsigned(wire233[(1'h1):(1'h1)]));
      for (forvar235 = (1'h0); (forvar235 < (2'h2)); forvar235 = (forvar235 + (1'h1)))
        begin
          for (forvar236 = (1'h0); (forvar236 < (1'h0)); forvar236 = (forvar236 + (1'h1)))
            begin
              reg237 = wire208;
              reg238 <= (~^reg219[(4'he):(4'hb)]);
              reg239 = {forvar236[(4'h8):(3'h4)],
                  ({$unsigned(reg226[(3'h5):(3'h4)])} ?
                      (reg238[(4'hd):(4'h8)] ?
                          {forvar236[(5'h10):(4'hf)]} : {(reg234 ?
                                  reg229 : wire207),
                              reg221[(4'h8):(2'h2)]}) : {$unsigned((wire210 * (8'ha6))),
                          $unsigned($unsigned(forvar236))})};
            end
          for (forvar240 = (1'h0); (forvar240 < (2'h3)); forvar240 = (forvar240 + (1'h1)))
            begin
              reg241 <= ((reg218 & $unsigned($signed(reg219[(1'h0):(1'h0)]))) * ((wire208[(1'h1):(1'h1)] ?
                  forvar218 : reg214[(1'h1):(1'h1)]) ^ {(~^(~&reg218)),
                  {(reg238 - (8'hb6)), $signed(forvar225)}}));
              reg242 <= (wire206 ?
                  (~$unsigned(((wire207 ?
                      forvar218 : reg229) <= reg241))) : forvar235[(4'h9):(4'h9)]);
              reg243 = (((reg234 + $signed((-reg230))) ?
                  reg228[(1'h1):(1'h0)] : $unsigned(reg223[(5'h11):(3'h5)])) + $signed((wire204[(1'h0):(1'h0)] <= reg230[(3'h6):(2'h2)])));
            end
          reg244 <= (($signed({(reg218 ~^ (8'hb3)),
                  (^~reg238)}) ~^ (^$signed(forvar235))) ?
              reg239 : ({$signed(reg211),
                      ((8'ha5) ? $signed(reg237) : $unsigned((8'h9e)))} ?
                  (^$unsigned({reg229})) : reg223[(3'h4):(2'h2)]));
        end
      for (forvar245 = (1'h0); (forvar245 < (3'h4)); forvar245 = (forvar245 + (1'h1)))
        begin
          for (forvar246 = (1'h0); (forvar246 < (2'h2)); forvar246 = (forvar246 + (1'h1)))
            begin
              reg247 <= ({(reg214[(1'h0):(1'h0)] ^ ((8'hb3) ^~ reg242[(4'h9):(4'h9)]))} ?
                  $signed({(~(^reg234)),
                      (~^(|wire205))}) : {$unsigned(reg244[(2'h2):(2'h2)])});
              reg248 = reg243[(3'h7):(2'h2)];
              reg249 = $unsigned($unsigned({$signed(wire208)}));
              reg250 = (7'h42);
            end
          if (wire209[(3'h6):(1'h0)])
            begin
              reg251 <= reg212;
              reg252 <= (^$unsigned(($signed($signed(reg249)) ?
                  (-$unsigned(reg229)) : (8'hb1))));
            end
          else
            begin
              reg251 <= reg213;
            end
          for (forvar253 = (1'h0); (forvar253 < (2'h3)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 <= {((7'h44) ^ (&((8'haf) != reg227[(4'he):(4'h8)]))),
                  forvar218};
              reg255 = $signed((~^$unsigned($signed(wire205))));
              reg256 <= forvar236[(3'h6):(3'h4)];
            end
        end
      reg257 <= ($unsigned($unsigned(((reg229 ?
              reg221 : reg212) <= (~|reg241)))) ?
          forvar235 : ({(!$signed(forvar245))} >>> $signed($unsigned(forvar225[(3'h7):(3'h7)]))));
      reg258 <= (reg254[(2'h2):(2'h2)] ?
          $unsigned((~|(forvar246 <<< (reg249 ?
              reg241 : wire208)))) : ($signed((&(+(8'hba)))) ?
              $unsigned(reg227[(4'hf):(1'h0)]) : $signed(reg220)));
    end
  always
    @(posedge clk) begin
      if ((^~((reg214[(2'h2):(1'h0)] <= (~|$unsigned(reg258))) <= $unsigned($unsigned(((8'hae) ^ reg212))))))
        begin
          reg259 = (&(8'h9d));
          for (forvar260 = (1'h0); (forvar260 < (1'h0)); forvar260 = (forvar260 + (1'h1)))
            begin
              reg261 = ((~^((^~(reg234 ?
                  forvar235 : reg218)) - (~^reg239[(3'h4):(1'h1)]))) >= $signed((($unsigned(reg221) ^~ $unsigned(forvar235)) ^ (8'h9c))));
              reg262 <= $unsigned(reg258);
              reg263 = ((reg239[(2'h3):(1'h0)] || $signed(($unsigned(reg250) == wire232))) ?
                  $signed($signed(reg256)) : $unsigned((($unsigned(reg247) << forvar260) ?
                      (reg241[(1'h1):(1'h1)] | (wire204 + reg220)) : $unsigned({reg257,
                          forvar245}))));
            end
        end
      else
        begin
          for (forvar259 = (1'h0); (forvar259 < (1'h1)); forvar259 = (forvar259 + (1'h1)))
            begin
              reg260 <= reg255[(4'h8):(3'h4)];
            end
        end
      reg264 = reg257[(1'h0):(1'h0)];
      reg265 <= (forvar245 >>> reg215);
    end
  assign wire266 = reg238;
endmodule

module module97  (y, clk, wire101, wire100, wire99, wire98);
  output wire [(32'h4ca):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire101;
  input wire signed [(5'h16):(1'h0)] wire100;
  input wire [(3'h7):(1'h0)] wire99;
  input wire signed [(3'h5):(1'h0)] wire98;
  wire signed [(5'h12):(1'h0)] wire197;
  wire [(4'hd):(1'h0)] wire196;
  wire [(3'h5):(1'h0)] wire195;
  wire signed [(5'h15):(1'h0)] wire194;
  reg [(4'hf):(1'h0)] reg193 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg192 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar190 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg189 = (1'h0);
  reg [(5'h11):(1'h0)] reg188 = (1'h0);
  reg [(5'h14):(1'h0)] reg187 = (1'h0);
  reg [(5'h12):(1'h0)] forvar186 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg184 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg183 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar182 = (1'h0);
  reg [(5'h13):(1'h0)] forvar181 = (1'h0);
  reg [(2'h3):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar171 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg180 = (1'h0);
  reg [(3'h4):(1'h0)] reg179 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg178 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar177 = (1'h0);
  reg [(5'h12):(1'h0)] reg176 = (1'h0);
  reg [(5'h10):(1'h0)] reg175 = (1'h0);
  reg [(2'h3):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg172 = (1'h0);
  reg [(5'h13):(1'h0)] reg171 = (1'h0);
  reg [(4'h8):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg169 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg168 = (1'h0);
  reg [(5'h13):(1'h0)] reg167 = (1'h0);
  reg [(2'h2):(1'h0)] reg166 = (1'h0);
  reg [(2'h3):(1'h0)] forvar165 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg164 = (1'h0);
  reg [(5'h12):(1'h0)] reg163 = (1'h0);
  reg [(4'he):(1'h0)] reg162 = (1'h0);
  reg [(5'h13):(1'h0)] reg161 = (1'h0);
  reg [(5'h16):(1'h0)] reg160 = (1'h0);
  reg [(4'hb):(1'h0)] forvar159 = (1'h0);
  reg [(5'h13):(1'h0)] forvar158 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg157 = (1'h0);
  reg [(2'h2):(1'h0)] reg156 = (1'h0);
  reg [(4'hd):(1'h0)] reg155 = (1'h0);
  reg [(5'h15):(1'h0)] forvar154 = (1'h0);
  reg [(5'h16):(1'h0)] reg153 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg150 = (1'h0);
  reg [(4'ha):(1'h0)] reg149 = (1'h0);
  reg [(5'h16):(1'h0)] reg148 = (1'h0);
  reg [(3'h5):(1'h0)] forvar147 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar146 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire145;
  wire signed [(4'he):(1'h0)] wire144;
  reg [(4'h8):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar135 = (1'h0);
  reg [(2'h2):(1'h0)] reg132 = (1'h0);
  reg [(4'hc):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg143 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg142 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg141 = (1'h0);
  reg [(3'h6):(1'h0)] reg140 = (1'h0);
  reg signed [(4'he):(1'h0)] reg139 = (1'h0);
  reg [(5'h11):(1'h0)] forvar138 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg137 = (1'h0);
  reg [(5'h11):(1'h0)] reg136 = (1'h0);
  reg [(4'hf):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg134 = (1'h0);
  reg [(4'h8):(1'h0)] reg133 = (1'h0);
  reg [(4'hf):(1'h0)] forvar132 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg131 = (1'h0);
  reg [(4'hc):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg129 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg128 = (1'h0);
  reg [(3'h4):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar126 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg125 = (1'h0);
  reg [(5'h15):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg123 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg122 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar121 = (1'h0);
  reg [(2'h3):(1'h0)] forvar120 = (1'h0);
  reg [(4'hd):(1'h0)] reg119 = (1'h0);
  reg [(2'h3):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg117 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg116 = (1'h0);
  reg signed [(4'he):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg114 = (1'h0);
  reg [(4'h9):(1'h0)] reg113 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar112 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg111 = (1'h0);
  reg [(4'h9):(1'h0)] reg110 = (1'h0);
  reg [(4'hc):(1'h0)] reg109 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg108 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg106 = (1'h0);
  reg [(5'h10):(1'h0)] reg105 = (1'h0);
  reg [(5'h12):(1'h0)] forvar103 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg104 = (1'h0);
  reg [(2'h2):(1'h0)] reg103 = (1'h0);
  reg [(4'h8):(1'h0)] reg102 = (1'h0);
  assign y = {wire197,
                 wire196,
                 wire195,
                 wire194,
                 reg193,
                 reg192,
                 reg191,
                 forvar190,
                 reg189,
                 reg188,
                 reg187,
                 forvar186,
                 reg185,
                 reg184,
                 reg183,
                 forvar182,
                 forvar181,
                 reg177,
                 forvar171,
                 reg180,
                 reg179,
                 reg178,
                 forvar177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 forvar165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 forvar159,
                 forvar158,
                 reg157,
                 reg156,
                 reg155,
                 forvar154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 forvar147,
                 forvar146,
                 wire145,
                 wire144,
                 reg138,
                 forvar135,
                 reg132,
                 reg126,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 forvar138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 forvar132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 forvar126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 forvar121,
                 forvar120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 forvar112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 forvar103,
                 reg104,
                 reg103,
                 reg102,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (($signed((~&$unsigned(((8'ha1) + wire98)))) << $unsigned((wire100[(5'h15):(5'h15)] >>> wire101[(2'h2):(1'h0)]))))
        begin
          reg102 <= $signed($signed((!(wire98[(2'h2):(1'h0)] ?
              ((8'hb7) ? wire101 : (8'hb4)) : (wire98 ? (8'ha4) : (8'hb2))))));
          reg103 = wire98[(1'h0):(1'h0)];
          reg104 = wire101[(1'h1):(1'h0)];
        end
      else
        begin
          reg102 <= (((-$unsigned((reg102 ? reg104 : wire100))) ?
              wire100[(3'h7):(3'h5)] : (~({reg104} > (&wire100)))) - ({((!wire101) ^~ wire100),
                  (-(reg104 ? reg104 : wire101))} ?
              ({{reg104, wire101}} ?
                  ((8'ha2) ?
                      (wire100 ^~ reg104) : $unsigned(reg103)) : ($unsigned(reg104) <= reg102)) : (8'hbf)));
          for (forvar103 = (1'h0); (forvar103 < (1'h0)); forvar103 = (forvar103 + (1'h1)))
            begin
              reg104 = wire98[(3'h4):(2'h2)];
              reg105 <= reg102[(4'h8):(2'h3)];
              reg106 <= reg102[(2'h3):(1'h0)];
            end
          if ((^reg106[(3'h6):(3'h4)]))
            begin
              reg107 = ($unsigned(reg106[(1'h0):(1'h0)]) != $signed($unsigned(((8'hb3) ?
                  wire101 : $signed(forvar103)))));
              reg108 <= reg105[(4'h8):(1'h0)];
              reg109 <= $unsigned({{wire98[(3'h4):(2'h3)]}});
              reg110 = ((wire99 + $unsigned($signed(reg104))) ?
                  (reg107 ?
                      (&{(~reg105),
                          wire100}) : wire101[(1'h0):(1'h0)]) : $signed(reg107));
            end
          else
            begin
              reg107 = forvar103[(5'h11):(1'h0)];
              reg108 = (+(^$signed({((8'ha6) ? reg107 : reg108)})));
              reg109 = wire98[(1'h0):(1'h0)];
            end
        end
      reg111 = (8'ha3);
      for (forvar112 = (1'h0); (forvar112 < (2'h3)); forvar112 = (forvar112 + (1'h1)))
        begin
          if ({(&{$signed(((8'hbb) ? reg110 : wire99))}),
              wire101[(1'h0):(1'h0)]})
            begin
              reg113 <= (&reg110);
              reg114 <= $signed(reg106[(2'h3):(2'h3)]);
              reg115 = reg104[(3'h6):(1'h1)];
            end
          else
            begin
              reg113 <= ((^~wire99) ~^ reg110[(1'h1):(1'h1)]);
              reg114 = wire101;
              reg115 = (reg107[(3'h4):(1'h1)] == (wire101[(1'h0):(1'h0)] ?
                  ($signed($signed(reg106)) && $signed($unsigned(reg104))) : (forvar103 > ((reg114 ?
                          wire99 : reg107) ?
                      (8'hb4) : (^reg107)))));
            end
          if ($unsigned(($unsigned(((reg106 ?
                  reg113 : reg105) | (reg113 >= reg110))) ?
              $unsigned(wire99[(3'h6):(2'h3)]) : (8'ha3))))
            begin
              reg116 = reg115[(1'h0):(1'h0)];
              reg117 <= reg116[(2'h2):(1'h0)];
              reg118 = {{$unsigned(((reg106 ? forvar103 : wire101) <= reg110))},
                  (&((-$unsigned(reg106)) ? wire99 : {(^reg109), (8'haa)}))};
            end
          else
            begin
              reg116 <= (reg103[(2'h2):(1'h0)] > ($signed(({reg117,
                      reg113} << ((8'hbe) ? reg116 : wire99))) ?
                  (8'h9c) : reg108));
              reg117 <= reg105[(4'hb):(1'h1)];
              reg118 <= $unsigned(wire100);
            end
          reg119 <= (reg115 ^~ (reg117[(4'ha):(4'h8)] ?
              reg115[(1'h1):(1'h1)] : reg109));
        end
      for (forvar120 = (1'h0); (forvar120 < (1'h0)); forvar120 = (forvar120 + (1'h1)))
        begin
          for (forvar121 = (1'h0); (forvar121 < (1'h0)); forvar121 = (forvar121 + (1'h1)))
            begin
              reg122 = reg106;
              reg123 <= {((~reg122) ?
                      $unsigned((wire100[(1'h0):(1'h0)] - $unsigned(reg105))) : forvar120)};
            end
        end
      reg124 = $signed((~$unsigned($unsigned(reg103))));
    end
  always
    @(posedge clk) begin
      reg125 = $signed((8'hb4));
      if ($signed(wire99[(2'h3):(1'h0)]))
        begin
          for (forvar126 = (1'h0); (forvar126 < (1'h1)); forvar126 = (forvar126 + (1'h1)))
            begin
              reg127 = $signed(reg108[(3'h4):(2'h3)]);
              reg128 = $unsigned($unsigned(reg107[(1'h1):(1'h1)]));
              reg129 = (&(wire99[(1'h0):(1'h0)] ^ $signed((8'hb2))));
              reg130 <= (&(forvar120[(1'h1):(1'h0)] ~^ $unsigned($signed(reg127[(2'h2):(1'h1)]))));
            end
          reg131 <= reg124[(3'h6):(3'h5)];
          for (forvar132 = (1'h0); (forvar132 < (3'h4)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 <= ((+($signed((|reg104)) && (8'hb2))) && (((&(reg106 ?
                      reg118 : reg130)) ?
                  ((+forvar112) == $unsigned((8'hbd))) : ($unsigned(forvar112) > (reg106 ?
                      reg110 : reg130))) || (((reg123 ? reg117 : reg113) ?
                  wire98 : $unsigned(reg110)) ^~ forvar126[(3'h4):(1'h1)])));
              reg134 = (+reg129);
              reg135 = reg111;
              reg136 = reg123[(1'h0):(1'h0)];
              reg137 = $unsigned($unsigned($unsigned(($signed(reg110) | (~reg105)))));
            end
          for (forvar138 = (1'h0); (forvar138 < (2'h3)); forvar138 = (forvar138 + (1'h1)))
            begin
              reg139 <= ((~$unsigned((~&{reg127,
                  reg103}))) < ($signed((&reg127[(2'h3):(2'h3)])) ?
                  forvar112 : (&wire101[(1'h1):(1'h1)])));
            end
          if (({(reg116 && (!reg119))} ?
              $signed(((&(8'ha6)) <<< (^~$signed(wire101)))) : wire98))
            begin
              reg140 <= reg102[(1'h0):(1'h0)];
              reg141 = reg130;
              reg142 <= reg116;
              reg143 = {(|(8'haa)), reg114[(3'h6):(3'h6)]};
            end
          else
            begin
              reg140 <= $unsigned({reg115,
                  (reg113 ?
                      (~$signed((8'ha8))) : $unsigned(reg129[(1'h1):(1'h1)]))});
              reg141 = $signed((^~wire98));
              reg142 <= {($signed(wire100) | reg107[(4'h9):(4'h8)]), reg110};
            end
        end
      else
        begin
          if (reg134[(3'h7):(1'h1)])
            begin
              reg126 <= $unsigned(((+$unsigned(reg128)) ?
                  $signed($signed(reg118[(1'h1):(1'h1)])) : reg123[(4'hf):(4'hc)]));
            end
          else
            begin
              reg126 <= $unsigned(($signed(forvar112[(1'h0):(1'h0)]) ?
                  ((^~$signed(reg126)) ?
                      (reg130 << $signed(reg142)) : forvar126[(3'h7):(3'h7)]) : {reg109[(4'h9):(2'h3)],
                      reg110[(4'h9):(3'h6)]}));
              reg127 = (($signed($unsigned($unsigned(reg141))) >>> (8'hac)) + ((({reg125,
                  reg119} != reg127) ^ reg133[(1'h1):(1'h1)]) & $signed(($signed(reg119) <= $unsigned(reg115)))));
              reg128 = $signed(($signed(($signed(reg123) == {reg134,
                  (8'hbf)})) ^~ reg131));
              reg129 = $signed(wire99);
              reg130 <= reg117;
            end
          reg131 <= {(^$unsigned($signed((~^reg124)))),
              ($signed(($signed(reg130) ~^ (~|reg139))) * (^((reg130 < reg115) >= (|reg108))))};
          if ($signed($unsigned((reg123 ?
              (~&(reg129 <<< forvar121)) : $unsigned((-(8'ha6)))))))
            begin
              reg132 = (+reg137[(3'h4):(3'h4)]);
              reg133 <= $unsigned($signed((!$signed((-reg141)))));
            end
          else
            begin
              reg132 <= (8'hb9);
              reg133 = (+(~&(!{$signed(forvar126)})));
              reg134 = reg116[(2'h2):(2'h2)];
            end
          for (forvar135 = (1'h0); (forvar135 < (3'h4)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= ((reg122[(1'h1):(1'h1)] ^~ (reg128 && (~{reg124}))) > ((8'ha8) * $signed($unsigned(reg118))));
              reg137 <= $signed((+{(~&(^~forvar112))}));
              reg138 <= $unsigned(reg140[(2'h3):(2'h3)]);
              reg139 = ($signed($signed($signed({reg119,
                  reg107}))) | reg131[(3'h6):(3'h4)]);
            end
        end
    end
  assign wire144 = (((((~reg118) ?
                           $signed(reg113) : $signed(reg126)) ^ $unsigned(reg111)) ^~ $signed(reg117)) ?
                       $signed($unsigned((|(+(8'hb5))))) : (~&$unsigned($unsigned((~wire98)))));
  assign wire145 = $signed($signed({$unsigned($unsigned(reg113))}));
  always
    @(posedge clk) begin
      for (forvar146 = (1'h0); (forvar146 < (2'h3)); forvar146 = (forvar146 + (1'h1)))
        begin
          for (forvar147 = (1'h0); (forvar147 < (1'h0)); forvar147 = (forvar147 + (1'h1)))
            begin
              reg148 = (^(reg113 ?
                  (!((reg113 & reg127) ?
                      $unsigned(wire145) : {forvar126,
                          wire145})) : reg129[(2'h2):(1'h0)]));
            end
          if ((~&forvar147[(1'h0):(1'h0)]))
            begin
              reg149 = $unsigned((^~(reg104[(3'h6):(2'h3)] && (reg138 ?
                  ((8'hac) ? forvar132 : forvar146) : (~&reg128)))));
              reg150 <= (wire101 ?
                  $signed(reg111) : ({{reg118[(2'h2):(2'h2)]}} ?
                      $unsigned($unsigned(reg118[(1'h1):(1'h0)])) : $unsigned(({reg124,
                          reg141} * (reg118 ? wire99 : (8'hae))))));
              reg151 = (~&$signed(reg134[(1'h1):(1'h1)]));
              reg152 <= $signed({$unsigned((8'hb5))});
              reg153 <= (&reg108);
            end
          else
            begin
              reg149 = (((-$unsigned(wire100[(2'h3):(2'h3)])) ?
                  reg117[(4'hc):(4'h9)] : reg143) || reg143[(3'h5):(3'h5)]);
              reg150 = $signed(((({reg153} ?
                  (+reg136) : $unsigned((7'h45))) <= ((reg153 >> wire101) == {forvar112})) << $signed(((~|reg118) ?
                  $signed(reg133) : (|reg152)))));
              reg151 = $unsigned(reg102);
            end
          for (forvar154 = (1'h0); (forvar154 < (1'h0)); forvar154 = (forvar154 + (1'h1)))
            begin
              reg155 <= (+reg139[(4'h8):(2'h3)]);
              reg156 <= ((+({{wire99}, (reg135 ? reg136 : reg128)} ?
                  (~|(reg113 ?
                      (8'hb1) : reg117)) : $signed($signed(reg118)))) & reg116);
              reg157 <= (((8'hb9) + ((wire145[(1'h1):(1'h0)] ?
                          reg103 : (reg138 ? reg110 : (8'ha1))) ?
                      ({reg105, reg103} ^ (&reg113)) : ((reg127 ?
                              wire145 : reg141) ?
                          (reg105 >> reg143) : (reg140 >= reg124)))) ?
                  $unsigned(({{forvar126}, {(8'ha2)}} * reg140)) : (8'hb1));
            end
        end
      for (forvar158 = (1'h0); (forvar158 < (3'h4)); forvar158 = (forvar158 + (1'h1)))
        begin
          for (forvar159 = (1'h0); (forvar159 < (1'h0)); forvar159 = (forvar159 + (1'h1)))
            begin
              reg160 <= (wire101[(1'h1):(1'h0)] ?
                  reg133[(3'h4):(2'h3)] : ($signed(wire145) ~^ ((8'hb4) ?
                      reg132[(1'h1):(1'h1)] : reg123[(3'h7):(3'h5)])));
              reg161 <= ($signed((forvar146[(3'h7):(2'h2)] ?
                      $signed((!reg134)) : (reg133 ?
                          reg114 : reg125[(3'h4):(1'h1)]))) ?
                  wire145 : ($signed($unsigned($signed(forvar138))) ?
                      ($signed(reg123[(4'hb):(4'h8)]) ?
                          reg107[(4'hb):(3'h6)] : ((reg115 ^~ (8'ha1)) ~^ (reg157 ?
                              wire101 : reg137))) : (reg155 * {(^(8'hb3)),
                          (~reg105)})));
              reg162 <= {reg157[(1'h1):(1'h1)], reg157[(4'h8):(4'h8)]};
              reg163 = reg107[(2'h2):(2'h2)];
            end
          reg164 = $signed((reg127[(2'h3):(2'h3)] < ((~^((7'h40) ~^ (7'h46))) >> $unsigned(reg130[(3'h5):(3'h5)]))));
          for (forvar165 = (1'h0); (forvar165 < (1'h0)); forvar165 = (forvar165 + (1'h1)))
            begin
              reg166 <= ($unsigned({((^reg115) != {(7'h40), reg119}),
                      {(&reg108)}}) ?
                  $unsigned({reg128}) : $unsigned((($signed(wire144) ?
                          $signed(reg110) : forvar154[(4'hb):(2'h3)]) ?
                      ((!reg108) >= $signed(reg130)) : (~^{reg125}))));
              reg167 = $signed((~^($signed(reg105[(3'h6):(3'h4)]) ?
                  ((forvar138 ? reg129 : reg111) ?
                      $unsigned(reg116) : $unsigned(reg108)) : $signed((forvar159 != reg105)))));
              reg168 = (!reg155[(4'hc):(4'h9)]);
            end
          reg169 = (reg133[(3'h7):(3'h4)] ?
              $signed(reg148[(4'h9):(3'h7)]) : ({($unsigned(forvar103) ?
                      ((7'h41) ~^ reg135) : $unsigned((8'had)))} && reg143[(1'h0):(1'h0)]));
        end
      if (((($unsigned((forvar132 ? wire99 : reg132)) ?
          (-(reg141 ?
              reg117 : wire145)) : $signed((reg138 >> forvar158))) != reg140) <<< ((!reg169) || (((reg139 ?
          reg114 : reg148) | forvar103[(4'he):(4'hc)]) - forvar103))))
        begin
          if (forvar126)
            begin
              reg170 <= $signed($unsigned($unsigned($unsigned(forvar154))));
            end
          else
            begin
              reg170 <= reg142[(1'h0):(1'h0)];
              reg171 <= (8'hb0);
              reg172 = $unsigned($signed(($signed((+wire98)) ?
                  (reg116[(1'h0):(1'h0)] - $unsigned(reg167)) : reg148[(4'he):(1'h1)])));
              reg173 <= $unsigned($signed($signed(reg169[(3'h6):(3'h6)])));
              reg174 = $unsigned((wire101[(1'h0):(1'h0)] ^ $unsigned((8'ha8))));
            end
          reg175 <= reg114;
          reg176 <= $unsigned($signed($unsigned((reg140 ?
              (reg143 ? reg174 : reg119) : forvar132[(4'h9):(4'h9)]))));
          for (forvar177 = (1'h0); (forvar177 < (1'h0)); forvar177 = (forvar177 + (1'h1)))
            begin
              reg178 = ($signed(reg135[(2'h3):(1'h0)]) ?
                  ($unsigned((-(&reg170))) ~^ {reg156[(1'h1):(1'h1)]}) : reg128[(1'h0):(1'h0)]);
              reg179 = (reg164 >>> $signed(((8'h9f) == ($signed(forvar154) ?
                  $signed(reg164) : (+reg123)))));
              reg180 <= reg125;
            end
        end
      else
        begin
          reg170 <= reg141;
          for (forvar171 = (1'h0); (forvar171 < (2'h2)); forvar171 = (forvar171 + (1'h1)))
            begin
              reg172 <= wire144;
              reg173 = ($unsigned((^$signed({reg172,
                  forvar165}))) >= {$signed((((8'hba) ?
                      reg152 : reg160) ^ (wire145 ? reg170 : forvar103))),
                  ($unsigned(reg137) ?
                      ((forvar126 | reg161) ~^ $signed(wire100)) : $signed((reg110 - reg174)))});
              reg174 <= (|(&(~&reg173)));
            end
          if (wire100[(5'h15):(4'h8)])
            begin
              reg175 = reg135;
              reg176 = reg179;
              reg177 <= reg131;
              reg178 = ((~^$signed((|reg155))) ?
                  reg172[(3'h7):(1'h0)] : $signed(($unsigned(((8'hbc) & reg175)) ?
                      (reg125[(3'h5):(2'h3)] >>> $unsigned(reg111)) : ((~&reg124) ?
                          (-reg152) : $unsigned(reg117)))));
            end
          else
            begin
              reg175 <= forvar121;
              reg176 <= reg140[(3'h6):(1'h0)];
              reg177 <= reg151;
              reg178 <= (~&(8'hbe));
              reg179 = {wire145[(2'h2):(2'h2)]};
            end
        end
      for (forvar181 = (1'h0); (forvar181 < (2'h3)); forvar181 = (forvar181 + (1'h1)))
        begin
          for (forvar182 = (1'h0); (forvar182 < (1'h1)); forvar182 = (forvar182 + (1'h1)))
            begin
              reg183 = ({(^reg162[(4'hb):(4'h8)]),
                  reg119[(3'h7):(1'h0)]} == reg155[(4'hc):(4'h8)]);
              reg184 <= (reg166[(1'h0):(1'h0)] ?
                  reg180 : (^reg168[(3'h4):(1'h1)]));
              reg185 = ($signed($unsigned(reg179)) ?
                  {$unsigned(((wire99 == reg153) ?
                          reg162[(4'he):(4'hd)] : forvar146[(3'h5):(2'h2)]))} : (8'hbf));
            end
        end
      for (forvar186 = (1'h0); (forvar186 < (2'h3)); forvar186 = (forvar186 + (1'h1)))
        begin
          if ({reg140[(3'h6):(2'h3)], forvar146})
            begin
              reg187 <= forvar147[(3'h5):(3'h4)];
              reg188 <= ((reg132 ?
                      (&(+$signed(forvar181))) : (~(-$signed(reg123)))) ?
                  ($unsigned($unsigned((reg185 - forvar154))) ?
                      reg117[(1'h1):(1'h0)] : ($unsigned($unsigned(reg172)) >>> (reg103[(1'h0):(1'h0)] ?
                          $signed(reg129) : (reg125 >>> (8'hb1))))) : ($unsigned((^~$signed(reg148))) != (!(reg174 < ((8'h9c) < reg149)))));
              reg189 = reg122;
            end
          else
            begin
              reg187 = (8'hab);
              reg188 = reg141[(4'he):(3'h6)];
            end
          for (forvar190 = (1'h0); (forvar190 < (1'h1)); forvar190 = (forvar190 + (1'h1)))
            begin
              reg191 = (($unsigned((~reg134[(4'hd):(4'h9)])) >= (reg115[(4'hb):(4'h8)] << ((~forvar190) != reg160))) * (8'hb6));
              reg192 = $unsigned({$signed($signed($unsigned((7'h40))))});
              reg193 = $unsigned($signed(reg179[(2'h3):(2'h2)]));
            end
        end
    end
  assign wire194 = reg129;
  assign wire195 = $signed($unsigned(reg134[(2'h3):(2'h3)]));
  assign wire196 = (^reg117[(4'h9):(3'h4)]);
  assign wire197 = (reg189 ? reg127 : $unsigned((~^(&$unsigned(reg185)))));
endmodule

module module278
#( parameter param442 = ((^({(~|(8'hb6)), ((7'h45) - (8'h9f))} ? (~|(^~(8'haa))) : ({(8'hac), (8'ha2)} << ((8'hb9) ? (8'ha0) : (8'hb1))))) ? (~|(!(+(!(7'h40))))) : ((+(^{(8'ha7)})) ? ((((7'h46) ? (8'ha3) : (7'h46)) - ((8'haa) ? (8'hb5) : (8'hb1))) ? {((8'hb6) + (8'hb6)), (~&(7'h42))} : (((8'hab) ? (7'h43) : (8'hb1)) >> (^(8'h9e)))) : ((((8'hbf) > (8'hb8)) ? {(7'h41)} : {(7'h44), (8'hae)}) - (((8'ha2) ? (8'ha8) : (8'ha2)) << ((8'h9c) & (8'ha0)))))) )
(y, clk, wire282, wire281, wire280, wire279);
  output wire [(32'h7d7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire282;
  input wire signed [(2'h2):(1'h0)] wire281;
  input wire signed [(5'h12):(1'h0)] wire280;
  input wire [(3'h6):(1'h0)] wire279;
  wire [(4'hb):(1'h0)] wire441;
  wire [(4'h8):(1'h0)] wire440;
  wire [(4'hb):(1'h0)] wire439;
  wire [(3'h4):(1'h0)] wire438;
  reg signed [(2'h3):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg432 = (1'h0);
  reg [(4'hf):(1'h0)] forvar427 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg436 = (1'h0);
  reg [(2'h2):(1'h0)] reg435 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg434 = (1'h0);
  reg [(3'h7):(1'h0)] reg433 = (1'h0);
  reg [(5'h13):(1'h0)] forvar432 = (1'h0);
  reg [(3'h6):(1'h0)] reg431 = (1'h0);
  reg [(4'hf):(1'h0)] reg430 = (1'h0);
  reg [(2'h2):(1'h0)] reg429 = (1'h0);
  reg [(5'h12):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg427 = (1'h0);
  reg [(5'h12):(1'h0)] reg426 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg425 = (1'h0);
  reg [(2'h2):(1'h0)] reg424 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg423 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg422 = (1'h0);
  reg [(3'h5):(1'h0)] reg421 = (1'h0);
  reg [(5'h15):(1'h0)] reg420 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg419 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg418 = (1'h0);
  reg [(2'h3):(1'h0)] forvar417 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg415 = (1'h0);
  reg [(4'hb):(1'h0)] reg414 = (1'h0);
  reg [(5'h10):(1'h0)] reg413 = (1'h0);
  reg [(4'hb):(1'h0)] reg412 = (1'h0);
  reg [(4'h9):(1'h0)] reg411 = (1'h0);
  reg [(3'h6):(1'h0)] reg410 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg409 = (1'h0);
  reg signed [(4'he):(1'h0)] reg408 = (1'h0);
  reg [(3'h4):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg404 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg403 = (1'h0);
  reg signed [(4'he):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg400 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar399 = (1'h0);
  reg signed [(4'he):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg398 = (1'h0);
  reg [(3'h4):(1'h0)] reg397 = (1'h0);
  reg [(5'h10):(1'h0)] reg396 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg395 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg394 = (1'h0);
  reg [(3'h7):(1'h0)] forvar393 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg392 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg391 = (1'h0);
  reg [(4'hd):(1'h0)] reg390 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar389 = (1'h0);
  reg [(5'h11):(1'h0)] forvar388 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg387 = (1'h0);
  reg [(4'ha):(1'h0)] reg386 = (1'h0);
  reg signed [(4'he):(1'h0)] reg385 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar384 = (1'h0);
  reg [(4'hd):(1'h0)] reg383 = (1'h0);
  reg [(4'h9):(1'h0)] reg382 = (1'h0);
  reg [(4'hc):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg380 = (1'h0);
  reg [(3'h6):(1'h0)] forvar379 = (1'h0);
  reg [(3'h4):(1'h0)] reg378 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg377 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg376 = (1'h0);
  reg [(5'h13):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg373 = (1'h0);
  reg signed [(4'he):(1'h0)] reg372 = (1'h0);
  reg [(4'he):(1'h0)] forvar371 = (1'h0);
  reg [(5'h10):(1'h0)] reg370 = (1'h0);
  reg signed [(4'he):(1'h0)] reg369 = (1'h0);
  reg [(4'h8):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg367 = (1'h0);
  reg [(4'ha):(1'h0)] reg366 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg365 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg363 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg359 = (1'h0);
  reg [(4'ha):(1'h0)] forvar358 = (1'h0);
  reg signed [(4'he):(1'h0)] reg362 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg361 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg360 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar359 = (1'h0);
  reg [(2'h3):(1'h0)] reg358 = (1'h0);
  reg [(4'hd):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg356 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg355 = (1'h0);
  reg [(2'h3):(1'h0)] reg354 = (1'h0);
  reg [(3'h7):(1'h0)] forvar353 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg352 = (1'h0);
  reg [(3'h5):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg350 = (1'h0);
  reg [(4'h9):(1'h0)] reg349 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg348 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg347 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar346 = (1'h0);
  reg [(4'he):(1'h0)] forvar340 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg344 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg343 = (1'h0);
  reg [(3'h5):(1'h0)] reg342 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg340 = (1'h0);
  reg signed [(4'he):(1'h0)] reg339 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg338 = (1'h0);
  reg [(4'ha):(1'h0)] reg337 = (1'h0);
  wire [(4'he):(1'h0)] wire336;
  wire signed [(5'h11):(1'h0)] wire335;
  wire signed [(4'h8):(1'h0)] wire334;
  reg [(3'h7):(1'h0)] reg333 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg332 = (1'h0);
  reg [(3'h4):(1'h0)] reg331 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg330 = (1'h0);
  reg [(5'h14):(1'h0)] reg329 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg327 = (1'h0);
  reg [(4'hc):(1'h0)] reg326 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg325 = (1'h0);
  reg [(4'hc):(1'h0)] reg324 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg323 = (1'h0);
  reg [(5'h14):(1'h0)] reg322 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg321 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg320 = (1'h0);
  reg [(4'hd):(1'h0)] reg319 = (1'h0);
  reg [(5'h15):(1'h0)] forvar318 = (1'h0);
  reg [(5'h13):(1'h0)] reg317 = (1'h0);
  reg [(3'h6):(1'h0)] reg316 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg315 = (1'h0);
  reg [(2'h3):(1'h0)] forvar314 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar304 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg313 = (1'h0);
  reg [(4'hb):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg310 = (1'h0);
  reg [(4'ha):(1'h0)] forvar309 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg308 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg307 = (1'h0);
  reg [(4'ha):(1'h0)] reg306 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg305 = (1'h0);
  reg [(4'hf):(1'h0)] reg304 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire303;
  wire [(3'h7):(1'h0)] wire302;
  reg signed [(4'h9):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg299 = (1'h0);
  reg [(4'ha):(1'h0)] reg298 = (1'h0);
  reg [(5'h14):(1'h0)] reg297 = (1'h0);
  reg [(4'ha):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg295 = (1'h0);
  reg [(4'he):(1'h0)] reg294 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg293 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg292 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg291 = (1'h0);
  reg [(5'h12):(1'h0)] reg290 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg289 = (1'h0);
  reg [(2'h3):(1'h0)] reg288 = (1'h0);
  reg [(3'h6):(1'h0)] reg287 = (1'h0);
  reg [(4'hb):(1'h0)] reg286 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg285 = (1'h0);
  reg [(5'h14):(1'h0)] reg284 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire283;
  assign y = {wire441,
                 wire440,
                 wire439,
                 wire438,
                 reg437,
                 reg432,
                 forvar427,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 forvar432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 forvar417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 forvar399,
                 reg393,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 forvar393,
                 reg392,
                 reg391,
                 reg390,
                 forvar389,
                 forvar388,
                 reg387,
                 reg386,
                 reg385,
                 forvar384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 forvar379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 forvar371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 reg359,
                 forvar358,
                 reg362,
                 reg361,
                 reg360,
                 forvar359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 forvar353,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 forvar346,
                 forvar340,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 wire336,
                 wire335,
                 wire334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 forvar318,
                 reg317,
                 reg316,
                 reg315,
                 forvar314,
                 forvar304,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 forvar309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 wire303,
                 wire302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 wire283,
                 (1'h0)};
  assign wire283 = ($unsigned({$signed((~^wire279)),
                       (wire279 ?
                           (wire282 ^ wire280) : (8'hb7))}) >>> wire280[(4'h8):(2'h3)]);
  always
    @(posedge clk) begin
      reg284 = wire281;
      reg285 <= (~|wire280[(4'ha):(1'h0)]);
      if ((+wire282))
        begin
          if ($unsigned(reg284))
            begin
              reg286 <= $signed($unsigned($signed(reg285[(4'hd):(1'h0)])));
              reg287 <= reg286[(3'h5):(1'h0)];
              reg288 = ({(((wire282 ? reg286 : (8'h9f)) ?
                          (^(8'ha8)) : reg284[(5'h13):(2'h3)]) ?
                      ({wire279,
                          reg287} - wire283) : $unsigned(wire281[(2'h2):(1'h1)])),
                  wire281} == $signed((reg287[(3'h4):(1'h0)] - $signed($signed(reg286)))));
            end
          else
            begin
              reg286 <= reg285[(2'h3):(1'h0)];
            end
          reg289 = (reg285 + (!($unsigned({(7'h45),
              reg285}) ~^ (((8'hb7) > wire279) + $unsigned(reg284)))));
          reg290 <= $unsigned($unsigned({reg288[(2'h3):(2'h2)]}));
        end
      else
        begin
          reg286 <= $unsigned(((($signed(wire279) ?
                  (!wire279) : wire279[(2'h3):(1'h0)]) ?
              (wire279[(2'h3):(1'h0)] ?
                  {reg290} : (wire283 << reg286)) : wire280) ^ (wire283[(2'h3):(2'h3)] & ($signed(reg284) ?
              (wire280 << reg290) : (reg287 | (7'h43))))));
          if (reg286[(3'h5):(3'h4)])
            begin
              reg287 <= $signed(reg285);
              reg288 = ($signed((~|$unsigned($signed(reg286)))) & ((8'hb4) && (~&((reg289 + reg289) << reg287))));
              reg289 = $signed((($unsigned(reg284) ?
                      {(reg285 || reg284)} : reg284[(3'h5):(3'h5)]) ?
                  (({(8'hb2),
                      wire282} > (reg285 * wire283)) & $unsigned(((8'hbe) ?
                      (8'hbd) : wire282))) : $unsigned((8'ha7))));
              reg290 <= reg285[(4'hb):(3'h7)];
              reg291 <= reg289;
            end
          else
            begin
              reg287 = {($signed($signed((wire280 <<< (8'hb9)))) & $unsigned((^~(8'hab)))),
                  (reg287[(3'h6):(3'h6)] >>> reg287)};
            end
          if ((wire282[(3'h4):(2'h2)] ?
              $unsigned((((|reg286) ? {wire279} : (8'had)) || {(|reg284),
                  wire282})) : ($signed(reg288[(1'h1):(1'h1)]) + (^~(reg285 || reg286[(3'h6):(2'h2)])))))
            begin
              reg292 = $unsigned((wire283 ?
                  (~$unsigned((reg291 >> wire280))) : reg290[(3'h5):(2'h2)]));
              reg293 = $unsigned(wire281[(1'h1):(1'h0)]);
              reg294 <= wire280[(3'h4):(3'h4)];
              reg295 = reg291[(4'h8):(3'h6)];
              reg296 = $unsigned((~($unsigned(reg292[(2'h3):(1'h0)]) > {(reg294 ~^ reg286)})));
            end
          else
            begin
              reg292 = (&reg293);
              reg293 = reg293[(1'h1):(1'h1)];
              reg294 <= reg288[(2'h2):(1'h0)];
              reg295 <= $signed($signed({wire281}));
              reg296 <= wire281[(2'h2):(1'h0)];
            end
          if (((&$unsigned($signed((8'ha1)))) ?
              $signed((+{$signed(reg295), $unsigned(reg294)})) : reg296))
            begin
              reg297 = $signed((~^(reg289 ?
                  (7'h41) : $signed($signed((8'hae))))));
              reg298 <= reg296[(4'h9):(1'h0)];
              reg299 <= $unsigned(($unsigned(reg286[(2'h3):(2'h2)]) >= (8'hbf)));
              reg300 = $unsigned(reg297);
            end
          else
            begin
              reg297 <= wire281;
              reg298 = reg287;
            end
        end
      reg301 = $unsigned((-{($signed(reg296) && {reg291})}));
    end
  assign wire302 = {$unsigned(reg285[(4'hb):(4'h8)])};
  assign wire303 = {$signed($signed(((~|wire280) ?
                           (reg284 - reg285) : wire302[(3'h7):(3'h6)])))};
  always
    @(posedge clk) begin
      if ((((&(reg284 & ((8'haa) << reg287))) ?
              (reg285 ~^ $unsigned(reg298[(4'h9):(3'h4)])) : (^reg288[(1'h0):(1'h0)])) ?
          $signed($unsigned((reg287[(1'h0):(1'h0)] ?
              (reg300 != reg298) : (wire302 ?
                  wire283 : reg293)))) : ($unsigned($signed(((8'hab) ~^ reg285))) ?
              (reg296 ?
                  wire279 : ($signed(reg294) ^~ (|wire302))) : reg289[(3'h6):(1'h1)])))
        begin
          if ($unsigned($signed($unsigned($unsigned($signed(wire303))))))
            begin
              reg304 <= (reg287[(3'h4):(3'h4)] ?
                  $signed(($unsigned($unsigned((8'hb9))) ^~ $signed((-(8'ha7))))) : $unsigned(reg299));
              reg305 <= (8'haa);
              reg306 = (($signed(reg292) ^~ $signed(reg290[(5'h12):(2'h2)])) ?
                  $signed($unsigned((reg286 <<< $unsigned(reg287)))) : ((8'hb1) ?
                      wire302 : (!($signed((8'hbf)) ?
                          $signed((8'hb5)) : {reg284, reg298}))));
              reg307 <= $signed($signed((reg284 & (^~reg301))));
              reg308 <= $unsigned($unsigned($signed($unsigned($signed((7'h40))))));
            end
          else
            begin
              reg304 = $unsigned((^reg291));
              reg305 = $unsigned((&{(reg294 ?
                      reg286 : (reg298 ? reg284 : reg304)),
                  $signed(((8'ha8) ^~ reg297))}));
              reg306 <= (^reg299);
            end
          for (forvar309 = (1'h0); (forvar309 < (3'h4)); forvar309 = (forvar309 + (1'h1)))
            begin
              reg310 = ((!(+reg288[(1'h1):(1'h1)])) ?
                  (-reg284[(4'hd):(3'h7)]) : ((((reg286 ?
                          wire303 : reg292) <<< (reg304 ? reg299 : reg306)) ?
                      reg287 : $signed(((8'hbc) ?
                          reg298 : wire283))) != (($signed(reg284) & $signed(reg290)) <<< $signed($signed(reg307)))));
              reg311 <= ($signed((~|reg297)) ?
                  ((~^{(~&reg285), (&reg298)}) ?
                      ($unsigned((+forvar309)) ?
                          $signed($unsigned(wire281)) : $unsigned(reg306)) : ((~^$signed(reg304)) & $signed((&(8'ha2))))) : (+reg287));
              reg312 <= $signed(reg296[(2'h3):(2'h2)]);
              reg313 <= $unsigned((($signed((|wire281)) << $signed(reg295)) >= {(reg295 ?
                      $signed(reg295) : $signed(reg305)),
                  reg307[(4'hc):(2'h3)]}));
            end
        end
      else
        begin
          for (forvar304 = (1'h0); (forvar304 < (2'h3)); forvar304 = (forvar304 + (1'h1)))
            begin
              reg305 <= reg306[(1'h0):(1'h0)];
            end
        end
      for (forvar314 = (1'h0); (forvar314 < (2'h3)); forvar314 = (forvar314 + (1'h1)))
        begin
          if ($unsigned((wire303[(3'h7):(3'h6)] == ((&{(8'h9d)}) | $signed((+forvar314))))))
            begin
              reg315 = ((reg300[(1'h0):(1'h0)] ?
                      $unsigned((reg308 == forvar314)) : (8'hb9)) ?
                  $signed((forvar309 - ($signed(reg284) ?
                      wire280 : {reg307}))) : (((^(reg284 ? wire283 : reg313)) ?
                      ($signed(reg287) ?
                          reg305 : (^~reg296)) : $unsigned($unsigned(wire281))) - reg310[(4'hd):(1'h0)]));
            end
          else
            begin
              reg315 <= (reg305[(1'h0):(1'h0)] ?
                  {(~&$unsigned((reg297 == (8'hb0))))} : (&((8'hae) ?
                      reg305 : $signed(reg307[(3'h5):(3'h4)]))));
            end
          reg316 = reg293[(2'h2):(1'h0)];
          reg317 = (!(reg288[(1'h1):(1'h1)] >= $unsigned(reg313[(1'h1):(1'h0)])));
          for (forvar318 = (1'h0); (forvar318 < (3'h4)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg319 <= reg289[(3'h5):(2'h3)];
              reg320 = $signed((^~{$unsigned((wire302 || wire280))}));
              reg321 = $signed((!$signed($signed(reg293))));
              reg322 = reg308;
            end
          reg323 = $signed({(8'hbb)});
        end
      if (reg288[(2'h2):(2'h2)])
        begin
          if ($unsigned($signed(reg295[(4'hd):(4'h9)])))
            begin
              reg324 <= reg321;
              reg325 = $signed(((~&((reg292 && reg323) >>> (reg317 | reg301))) * $unsigned(($signed(reg284) >> {(8'hbc),
                  reg285}))));
              reg326 = reg296[(2'h3):(1'h1)];
              reg327 = {{(!reg297[(4'he):(4'hc)])}};
              reg328 = (~^$unsigned($signed($unsigned($unsigned((8'hb0))))));
            end
          else
            begin
              reg324 <= ((~^{$signed($signed(reg306))}) & ($unsigned(reg321) - ($unsigned(reg327) ?
                  reg316[(3'h6):(1'h1)] : {(forvar314 ? (8'had) : reg315)})));
              reg325 = (~{(reg285 ? $signed(reg326) : reg313[(3'h6):(2'h3)])});
              reg326 <= $unsigned(($unsigned((-reg310[(1'h1):(1'h1)])) ?
                  $unsigned($unsigned((reg301 && reg294))) : reg325));
            end
          reg329 = (+$unsigned(({(8'ha4)} ^~ reg296)));
          reg330 <= $signed((reg322 ?
              {$signed((reg310 << reg326))} : $signed(reg325)));
          reg331 = $signed(reg324);
        end
      else
        begin
          if (reg321)
            begin
              reg324 <= $signed({reg319});
              reg325 <= reg330[(4'h9):(3'h5)];
              reg326 <= reg319;
            end
          else
            begin
              reg324 = (reg290[(4'h9):(3'h7)] + (reg312[(3'h5):(3'h5)] ?
                  (((reg292 ~^ reg329) >> reg323[(2'h3):(1'h1)]) || (^(reg293 ?
                      wire281 : forvar314))) : ((~|reg306[(2'h3):(1'h1)]) && (~^$signed((8'hb2))))));
              reg325 <= (&wire283);
              reg326 <= reg308[(4'hb):(4'hb)];
              reg327 = $signed(reg329[(4'ha):(2'h3)]);
            end
          reg328 <= reg316;
          if (reg289[(3'h4):(3'h4)])
            begin
              reg329 <= wire283;
              reg330 = (($signed({{(8'ha0)}}) ?
                      $signed(reg324[(4'h8):(3'h5)]) : $unsigned((~|(wire282 << reg315)))) ?
                  {{((!(8'ha1)) * {reg298, forvar304}),
                          (-$signed(wire302))}} : wire283);
              reg331 <= (~&reg327[(4'hb):(2'h2)]);
              reg332 <= $signed($unsigned(((reg293 ?
                      reg284[(2'h2):(2'h2)] : $unsigned(wire279)) ?
                  $signed($signed(reg285)) : $signed((~|reg288)))));
            end
          else
            begin
              reg329 <= $signed(((((reg305 ? reg316 : reg317) ?
                  (+reg306) : reg328[(4'hc):(1'h0)]) && $signed($unsigned(reg307))) <<< $signed(($signed((7'h44)) | reg294[(3'h5):(1'h0)]))));
            end
        end
      reg333 <= reg320;
    end
  assign wire334 = reg292;
  assign wire335 = (wire280[(4'hb):(4'h8)] ?
                       $unsigned(reg317) : $unsigned((wire281[(1'h0):(1'h0)] ?
                           $signed($signed((8'hb3))) : $unsigned($signed(reg316)))));
  assign wire336 = (reg325[(4'h9):(4'h9)] ?
                       reg321[(2'h2):(2'h2)] : $unsigned(reg324));
  always
    @(posedge clk) begin
      reg337 = reg313;
    end
  always
    @(posedge clk) begin
      reg338 <= ({(~^$unsigned({reg328})), (7'h42)} ^ (wire281[(2'h2):(1'h1)] ?
          reg288 : {(+$unsigned(wire282)), reg324}));
      reg339 = (~|$signed($unsigned($signed({reg330}))));
      if (wire280[(1'h0):(1'h0)])
        begin
          if (reg286)
            begin
              reg340 <= $unsigned(({$signed(reg333)} <= reg311));
              reg341 <= ($signed($unsigned(wire335[(5'h11):(3'h5)])) && reg315);
              reg342 = $unsigned($signed($signed($unsigned(((8'hb8) ?
                  (8'haa) : (8'hb4))))));
              reg343 = ((~reg325) >>> (wire334[(2'h3):(2'h3)] < ((wire302[(1'h1):(1'h1)] ?
                      reg310 : (reg341 ? reg312 : (7'h46))) ?
                  reg341 : reg296)));
            end
          else
            begin
              reg340 = ({$unsigned((8'hb9))} ?
                  $unsigned(wire279[(2'h3):(1'h0)]) : reg340[(4'hd):(4'h9)]);
              reg341 <= ($unsigned((wire336 ?
                  reg285[(3'h5):(2'h3)] : ($signed(reg330) + reg319))) ~^ (&wire335));
              reg342 <= reg289;
              reg343 = reg330;
              reg344 = reg300[(5'h11):(3'h5)];
            end
          reg345 <= reg338[(4'ha):(4'h9)];
        end
      else
        begin
          for (forvar340 = (1'h0); (forvar340 < (1'h1)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 = (&reg338);
              reg342 = $unsigned($signed($signed(forvar340[(1'h1):(1'h1)])));
              reg343 <= (|reg299);
              reg344 = (^$signed(($unsigned((~|reg344)) ?
                  $signed($unsigned(wire280)) : reg329)));
              reg345 = reg298;
            end
          for (forvar346 = (1'h0); (forvar346 < (2'h2)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 = reg292;
              reg348 <= (^~{((((7'h42) ? (8'ha2) : reg310) ?
                          (wire334 >>> reg321) : $unsigned(reg319)) ?
                      ($unsigned((8'ha5)) >>> (reg293 == reg311)) : {$signed(wire302),
                          $unsigned((7'h45))}),
                  (!reg288)});
              reg349 = ($unsigned((reg284 ?
                  ((reg300 ?
                      (8'hb6) : (8'h9d)) <<< reg325[(2'h2):(2'h2)]) : $signed(((8'hae) <<< reg328)))) ~^ reg307[(4'hb):(4'h8)]);
              reg350 = reg297[(1'h0):(1'h0)];
              reg351 = reg288;
            end
          reg352 <= reg286;
          for (forvar353 = (1'h0); (forvar353 < (1'h1)); forvar353 = (forvar353 + (1'h1)))
            begin
              reg354 <= $signed(($signed(((~|reg327) || $signed(reg299))) ?
                  wire334[(2'h2):(1'h1)] : reg307));
              reg355 = (reg350[(4'hf):(1'h1)] ^ {(($signed(forvar314) ?
                      (&reg341) : reg341) ~^ wire279),
                  $unsigned(((^~(8'hb7)) < $signed(reg298)))});
              reg356 = ((8'hbd) ?
                  $signed({reg341[(2'h3):(1'h0)]}) : (~|$signed(reg343)));
            end
          reg357 = reg339[(4'he):(4'hd)];
        end
      if ({reg328[(4'hc):(2'h3)]})
        begin
          reg358 = $unsigned(reg344[(3'h5):(1'h0)]);
          for (forvar359 = (1'h0); (forvar359 < (3'h4)); forvar359 = (forvar359 + (1'h1)))
            begin
              reg360 <= ((8'hbb) ^ $signed((~^forvar340[(3'h5):(3'h4)])));
              reg361 <= reg320[(1'h1):(1'h1)];
              reg362 = ($unsigned(reg355[(2'h2):(1'h0)]) ?
                  reg329 : {$unsigned($signed(reg320))});
            end
        end
      else
        begin
          for (forvar358 = (1'h0); (forvar358 < (2'h2)); forvar358 = (forvar358 + (1'h1)))
            begin
              reg359 <= forvar304[(3'h6):(2'h2)];
              reg360 = (8'hb8);
              reg361 = (7'h40);
            end
          reg362 = reg341[(4'hb):(2'h3)];
          if (reg343)
            begin
              reg363 = (&{reg349[(1'h1):(1'h1)]});
              reg364 <= ((+$unsigned(reg284)) <= reg313[(3'h7):(3'h4)]);
              reg365 = (reg344 ? wire302 : {$unsigned(wire280)});
            end
          else
            begin
              reg363 <= (forvar314[(1'h0):(1'h0)] - $unsigned($unsigned({((8'hac) == reg360)})));
              reg364 <= ($unsigned(reg312[(4'h8):(3'h7)]) ?
                  {(~^{reg323})} : $unsigned((&$signed((reg300 < reg311)))));
              reg365 <= (reg329[(4'h8):(2'h3)] << {$signed((|(~^reg329))),
                  $unsigned(wire279)});
              reg366 = reg296;
            end
          if ($signed(reg293))
            begin
              reg367 = (8'hb7);
              reg368 <= $signed((7'h40));
              reg369 <= $signed(reg347);
            end
          else
            begin
              reg367 = reg341;
              reg368 <= wire335[(1'h1):(1'h0)];
              reg369 = $signed(({reg338, ((~(8'ha3)) * (+reg367))} ?
                  reg289 : (&(|(+reg317)))));
              reg370 = $unsigned(((8'hb6) ? (!forvar318) : $signed({reg342})));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar371 = (1'h0); (forvar371 < (1'h0)); forvar371 = (forvar371 + (1'h1)))
        begin
          if (reg313)
            begin
              reg372 = $unsigned($unsigned((((reg357 <= reg327) ?
                  (reg348 <= (7'h45)) : {reg319}) != (^$signed(reg288)))));
              reg373 <= ($unsigned($signed($signed($unsigned(reg326)))) ?
                  reg348 : ((($unsigned(reg357) ?
                              $unsigned(reg298) : (~|(8'ha0))) ?
                          {(reg300 ? reg340 : reg322),
                              reg363[(5'h11):(4'ha)]} : ((!reg357) ?
                              (~|reg351) : (~&reg354))) ?
                      (($unsigned((8'hb1)) - forvar346) ?
                          ((~|reg297) || $unsigned(wire303)) : {(reg306 << reg301)}) : $unsigned(((reg319 ?
                          reg329 : (8'hb1)) * forvar318))));
              reg374 <= $unsigned((reg307 ?
                  $signed($signed((|reg354))) : reg338[(1'h1):(1'h0)]));
              reg375 <= wire280[(3'h6):(1'h0)];
              reg376 <= forvar318[(3'h5):(2'h3)];
            end
          else
            begin
              reg372 <= reg324;
            end
          reg377 <= {({reg365[(2'h2):(1'h0)], $signed(reg315[(2'h2):(1'h1)])} ?
                  (-(|reg316[(3'h5):(3'h4)])) : forvar318[(5'h12):(4'h9)])};
          reg378 = forvar314[(1'h1):(1'h0)];
          for (forvar379 = (1'h0); (forvar379 < (1'h1)); forvar379 = (forvar379 + (1'h1)))
            begin
              reg380 = reg357[(4'ha):(4'h8)];
              reg381 <= reg294;
              reg382 = ((((reg301 || (~reg315)) ?
                          ({reg323} ^ reg326) : reg338) ?
                      reg374 : $unsigned(reg359)) ?
                  reg351[(2'h3):(2'h3)] : $unsigned((reg319 >= forvar359)));
              reg383 <= forvar358[(1'h0):(1'h0)];
            end
          for (forvar384 = (1'h0); (forvar384 < (1'h1)); forvar384 = (forvar384 + (1'h1)))
            begin
              reg385 <= reg358[(2'h2):(2'h2)];
              reg386 <= reg348[(3'h6):(1'h0)];
              reg387 = (reg312 ?
                  $signed((reg337[(1'h0):(1'h0)] - $unsigned(reg297))) : $unsigned((+(8'hb3))));
            end
        end
      for (forvar388 = (1'h0); (forvar388 < (1'h0)); forvar388 = (forvar388 + (1'h1)))
        begin
          for (forvar389 = (1'h0); (forvar389 < (2'h2)); forvar389 = (forvar389 + (1'h1)))
            begin
              reg390 = $unsigned(reg308[(4'hf):(3'h5)]);
              reg391 = reg328;
              reg392 = wire280[(4'ha):(4'h9)];
            end
        end
    end
  always
    @(posedge clk) begin
      if ((reg326 || (-{reg391[(4'h9):(3'h6)]})))
        begin
          for (forvar393 = (1'h0); (forvar393 < (3'h4)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 <= ($signed($signed(((reg387 - reg378) == $signed(reg361)))) ?
                  ({reg381[(4'ha):(3'h6)]} <<< reg294) : reg286[(1'h0):(1'h0)]);
              reg395 = {(8'hbf),
                  (reg298 ?
                      (($signed(reg394) ?
                              $signed(forvar318) : $signed(reg344)) ?
                          $signed((reg368 ?
                              reg324 : reg310)) : $unsigned((reg288 ?
                              reg284 : reg341))) : ({(reg342 ?
                              (7'h45) : (8'ha7)),
                          $unsigned(forvar304)} | (reg339[(3'h6):(1'h0)] ?
                          (reg299 ?
                              (8'hb8) : reg373) : reg385[(4'hb):(4'ha)])))};
              reg396 = $signed((^~(reg340 ?
                  (!((8'haf) ?
                      forvar358 : (8'haf))) : ((~reg315) + $unsigned(reg394)))));
              reg397 = (&(&(((reg289 << forvar318) || $unsigned(reg358)) >= (reg361 ?
                  (reg305 == reg304) : (forvar393 - reg349)))));
            end
          reg398 <= reg291[(3'h4):(1'h1)];
        end
      else
        begin
          reg393 <= {((&$unsigned($signed(reg317))) && ((reg331[(1'h1):(1'h0)] ?
                  reg362 : (^~(8'hb9))) < ((^reg372) != $signed(reg370)))),
              reg380};
          if ($signed(($unsigned($unsigned((^~(7'h46)))) ?
              (!(^~{reg339, wire283})) : (!reg311[(4'hc):(4'hc)]))))
            begin
              reg394 <= $unsigned((+$signed(reg316[(3'h6):(2'h3)])));
              reg395 <= (~^(reg372[(4'h8):(2'h2)] ^ $signed($unsigned(reg345))));
              reg396 <= reg390[(4'ha):(3'h5)];
              reg397 = (~reg326);
              reg398 = (8'hb5);
            end
          else
            begin
              reg394 <= reg378[(3'h4):(2'h2)];
            end
          for (forvar399 = (1'h0); (forvar399 < (2'h2)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg400 = ({$signed($signed({reg365})),
                  $signed((reg339 ?
                      $unsigned(reg345) : $signed(reg310)))} < (~|$unsigned(reg300)));
              reg401 = reg332[(3'h4):(2'h3)];
              reg402 = ($unsigned(reg385[(3'h7):(3'h4)]) | reg377);
              reg403 <= wire283;
              reg404 <= ($unsigned((((^~reg327) * {reg292, reg374}) ?
                      reg316 : (reg343 ? reg366[(4'h8):(3'h7)] : (|reg378)))) ?
                  (|forvar304) : (~^(~&(~(forvar359 ? reg305 : forvar371)))));
            end
          reg405 <= (~^(~{$signed($unsigned((8'h9c)))}));
          if ({$unsigned($signed($unsigned((reg376 ^~ reg352)))),
              ((reg310[(3'h5):(1'h1)] ^~ reg338) < forvar384)})
            begin
              reg406 = $unsigned(reg340[(5'h10):(1'h1)]);
              reg407 = (|(7'h44));
              reg408 <= {$unsigned(reg325),
                  (-($signed($unsigned(reg284)) <= $signed(reg400)))};
              reg409 = ((+$signed(reg397[(1'h0):(1'h0)])) ~^ $signed((($unsigned((8'h9d)) * reg338) > $unsigned($unsigned(reg337)))));
              reg410 = reg320[(3'h4):(2'h2)];
            end
          else
            begin
              reg406 <= $signed($signed((+$unsigned({forvar353}))));
              reg407 <= reg362;
            end
        end
      if (({reg312[(4'h9):(3'h4)],
              (((~|forvar399) ?
                  reg364 : (wire335 ?
                      (8'h9c) : reg310)) >>> ((reg299 << wire281) ?
                  reg360 : $unsigned((8'ha2))))} ?
          reg351[(3'h4):(1'h0)] : {(~&reg410), (!reg364[(3'h4):(1'h1)])}))
        begin
          if ((($unsigned((((8'ha5) ? (8'hab) : reg355) ?
                      $unsigned(reg408) : reg323)) ?
                  $unsigned((-reg345)) : $signed($signed((!reg286)))) ?
              reg299 : ($signed($unsigned(reg351)) ^~ reg373)))
            begin
              reg411 <= {{(reg321[(2'h2):(1'h1)] ~^ ({reg329, reg343} ?
                          reg368 : $unsigned(reg343)))}};
              reg412 = reg381[(4'h9):(4'h8)];
              reg413 <= $signed(reg376);
              reg414 <= $unsigned($signed($signed(reg354[(1'h1):(1'h0)])));
              reg415 = reg294;
            end
          else
            begin
              reg411 <= (((((reg392 ? reg375 : forvar340) && (reg348 ?
                      reg356 : reg317)) << ($unsigned(reg397) ?
                      forvar304[(1'h1):(1'h1)] : $signed(reg347))) <<< $unsigned($unsigned((&reg330)))) ?
                  $signed($signed($signed({reg402}))) : $unsigned($unsigned(reg299)));
              reg412 <= $unsigned(($unsigned(reg342[(1'h1):(1'h1)]) >= ($signed((~&forvar353)) ?
                  ((~|reg295) ?
                      reg364 : (wire279 | reg381)) : $unsigned(forvar318))));
            end
        end
      else
        begin
          reg411 = ((reg396 ?
              ($unsigned((reg329 ^~ reg325)) ?
                  $signed((reg323 ?
                      reg320 : reg372)) : $unsigned(reg369)) : (($unsigned((7'h40)) << {forvar388,
                      reg362}) ?
                  reg364 : (8'ha1))) ^~ $unsigned((^($unsigned(reg400) ?
              (reg402 ~^ reg413) : ((7'h41) ? (8'ha6) : reg363)))));
          if (reg327)
            begin
              reg412 <= (|(~&forvar393));
              reg413 = $unsigned($signed((($signed(reg349) << reg304) ?
                  reg290[(4'h8):(1'h0)] : (8'ha0))));
              reg414 <= ((($unsigned((reg315 ^~ reg354)) ?
                  (reg332[(3'h5):(3'h4)] ?
                      reg325 : ((8'h9c) ?
                          forvar318 : reg316)) : ($signed(forvar379) - reg395[(1'h1):(1'h1)])) == $signed(reg410[(3'h4):(2'h3)])) && reg375[(4'h9):(3'h4)]);
              reg415 <= forvar346[(2'h3):(1'h1)];
            end
          else
            begin
              reg412 <= reg370[(4'hb):(3'h6)];
            end
          reg416 <= reg311;
          for (forvar417 = (1'h0); (forvar417 < (1'h1)); forvar417 = (forvar417 + (1'h1)))
            begin
              reg418 = (((reg287 ?
                      wire283[(3'h4):(1'h0)] : $signed($unsigned(reg316))) ?
                  $signed((reg323 & (|reg347))) : reg369[(4'h8):(3'h7)]) >>> forvar309);
              reg419 = (~^reg328[(4'he):(3'h6)]);
              reg420 = ((({forvar340} << {$unsigned(reg337)}) >>> ($unsigned(reg385[(2'h2):(1'h1)]) ?
                      (8'ha7) : $signed((reg354 > reg342)))) ?
                  reg308[(5'h13):(4'h8)] : $signed(((~^forvar340[(4'h9):(2'h3)]) & {reg321})));
              reg421 = $signed({((|$unsigned(reg349)) || wire280[(3'h7):(2'h2)]),
                  $signed(reg288)});
              reg422 = wire279;
            end
          if ((((((reg301 ? wire279 : wire303) <<< (reg285 ?
                  forvar304 : (8'hb6))) >> $unsigned((^~reg364))) <<< {{(reg402 ?
                          reg304 : reg387),
                      reg377},
                  ({reg286} ? $signed(reg398) : ((8'ha5) == reg383))}) ?
              $unsigned((forvar346 ?
                  reg372[(1'h0):(1'h0)] : ($unsigned(reg313) ?
                      reg331[(2'h3):(2'h3)] : (reg342 >> reg313)))) : reg401[(2'h3):(2'h2)]))
            begin
              reg423 = $unsigned($unsigned(reg324));
              reg424 <= reg385;
              reg425 = $unsigned($signed($unsigned((wire303 ^ wire282[(3'h6):(1'h1)]))));
              reg426 = forvar358[(3'h4):(1'h0)];
            end
          else
            begin
              reg423 = reg392[(4'hc):(4'h8)];
              reg424 = (^~{reg406,
                  ($signed((~reg347)) ?
                      reg420 : ((reg420 <= wire281) ?
                          $unsigned(reg320) : (reg395 & (8'hb6))))});
              reg425 = reg287[(2'h3):(2'h2)];
              reg426 = wire334;
            end
        end
      if ($unsigned($signed($unsigned(reg387[(1'h1):(1'h0)]))))
        begin
          if (reg330)
            begin
              reg427 <= $signed((reg404 ?
                  (!(^$signed(reg368))) : (($unsigned(reg307) ?
                          wire303 : (reg374 >> (7'h42))) ?
                      $unsigned((reg312 ?
                          reg299 : wire282)) : ($signed(reg409) >>> (reg349 <= reg351)))));
              reg428 <= ({((|reg308) ?
                      $signed((~reg408)) : ((forvar314 || reg390) ?
                          $signed(forvar359) : (reg289 ? forvar353 : reg293))),
                  reg310} < reg326[(3'h4):(2'h2)]);
              reg429 = ({reg359} ?
                  ($signed(reg321) || $unsigned($unsigned(reg350))) : $unsigned((^reg323)));
            end
          else
            begin
              reg427 = {(7'h45), (+{{$unsigned((8'h9d))}, (~(7'h46))})};
            end
          reg430 <= $signed((forvar358 ? $unsigned(reg316) : reg356));
          reg431 = {reg373};
          for (forvar432 = (1'h0); (forvar432 < (2'h3)); forvar432 = (forvar432 + (1'h1)))
            begin
              reg433 = reg368;
              reg434 = (reg307 <= reg429[(2'h2):(2'h2)]);
              reg435 = forvar379[(1'h1):(1'h1)];
              reg436 <= ($signed($signed({$signed(reg351)})) ?
                  ($signed($signed(reg428)) ?
                      (($unsigned(reg340) ? (~&reg386) : $signed((8'haf))) ?
                          reg397[(3'h4):(1'h0)] : $signed(reg339[(4'he):(2'h3)])) : reg338) : (7'h44));
            end
        end
      else
        begin
          for (forvar427 = (1'h0); (forvar427 < (2'h2)); forvar427 = (forvar427 + (1'h1)))
            begin
              reg428 <= (((($signed(reg422) ?
                          reg284[(4'h9):(1'h1)] : $signed(reg404)) ?
                      reg403[(1'h1):(1'h1)] : ((forvar388 ?
                          reg365 : reg311) + ((8'hbf) || (8'hb6)))) ?
                  (|(reg284 <<< reg345[(1'h0):(1'h0)])) : wire279[(1'h1):(1'h0)]) + $signed($signed((8'hbd))));
              reg429 <= reg329[(3'h4):(2'h2)];
              reg430 <= $unsigned((-$signed($signed($signed(reg289)))));
              reg431 = $unsigned($signed(forvar432));
            end
          reg432 = (~$unsigned((!$signed((reg420 < reg386)))));
        end
      reg437 = reg429[(1'h0):(1'h0)];
    end
  assign wire438 = $signed((&{$unsigned((reg394 > reg305)),
                       {$signed(reg426), reg320}}));
  assign wire439 = (((|(8'hb5)) ?
                           reg310 : $signed(($unsigned(reg437) & reg398[(1'h1):(1'h1)]))) ?
                       (~&reg355[(4'hb):(3'h7)]) : {$unsigned(reg311),
                           ((~^{reg405, reg431}) ?
                               ({reg329,
                                   reg411} * $unsigned(wire302)) : ($signed(reg351) ?
                                   $unsigned(reg396) : {reg393, (8'hae)}))});
  assign wire440 = $signed((reg393 - ((8'hbc) ? reg315 : (!(^reg312)))));
  assign wire441 = (reg427 | $unsigned(($signed(((8'hbe) ? (8'ha3) : reg337)) ?
                       $unsigned(reg327[(4'he):(3'h4)]) : (((7'h44) >>> reg380) < {reg368,
                           reg297}))));
endmodule