(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param2701 = (7'h4d), 
parameter param2702 = (param2701 ? (({((8'hae) != param2701), (7'h44)} + ((&param2701) ? {param2701} : (param2701 ? param2701 : param2701))) ? (((param2701 * param2701) - (+(8'hb7))) < (!(^param2701))) : (param2701 >>> {(param2701 ? param2701 : param2701), (~param2701)})) : (param2701 ? (~&(param2701 ? (param2701 ? param2701 : param2701) : (param2701 ? param2701 : param2701))) : ((~&{param2701}) ? (((8'ha2) ? param2701 : param2701) ^ param2701) : param2701))))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h144b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire0;
  input wire [(5'h1c):(1'h0)] wire1;
  input wire [(4'h8):(1'h0)] wire2;
  input wire [(5'h1a):(1'h0)] wire3;
  input wire [(5'h1d):(1'h0)] wire4;
  wire [(4'he):(1'h0)] wire2654;
  wire signed [(4'h9):(1'h0)] wire2653;
  wire signed [(4'h9):(1'h0)] wire2651;
  wire [(4'ha):(1'h0)] wire2508;
  wire signed [(4'he):(1'h0)] wire42;
  wire signed [(3'h5):(1'h0)] wire2453;
  reg [(5'h13):(1'h0)] reg2700 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2697 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2696 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2695 = (1'h0);
  reg [(5'h19):(1'h0)] reg2680 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2678 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2691 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2689 = (1'h0);
  reg [(4'hb):(1'h0)] reg2688 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2687 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2683 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2682 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2677 = (1'h0);
  reg [(5'h18):(1'h0)] reg2676 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2674 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2669 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2665 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2664 = (1'h0);
  reg [(4'he):(1'h0)] reg2661 = (1'h0);
  reg [(5'h12):(1'h0)] reg2660 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2659 = (1'h0);
  reg [(5'h1a):(1'h0)] reg5 = (1'h0);
  reg [(5'h1c):(1'h0)] reg6 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg8 = (1'h0);
  reg [(4'he):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg18 = (1'h0);
  reg [(5'h11):(1'h0)] reg22 = (1'h0);
  reg [(5'h1f):(1'h0)] reg25 = (1'h0);
  reg [(5'h13):(1'h0)] reg27 = (1'h0);
  reg [(5'h1c):(1'h0)] reg29 = (1'h0);
  reg [(5'h10):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg33 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg34 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg36 = (1'h0);
  reg [(5'h16):(1'h0)] reg2456 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2458 = (1'h0);
  reg [(4'hb):(1'h0)] reg2459 = (1'h0);
  reg [(4'hc):(1'h0)] reg2461 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2463 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2466 = (1'h0);
  reg [(5'h14):(1'h0)] reg2468 = (1'h0);
  reg [(5'h18):(1'h0)] reg2472 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2474 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2475 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2478 = (1'h0);
  reg [(4'hf):(1'h0)] reg2480 = (1'h0);
  reg [(4'h8):(1'h0)] reg2486 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2487 = (1'h0);
  reg [(4'hc):(1'h0)] reg2489 = (1'h0);
  reg [(4'hf):(1'h0)] reg2491 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2492 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2496 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2497 = (1'h0);
  reg [(4'hc):(1'h0)] reg2498 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2499 = (1'h0);
  reg [(5'h19):(1'h0)] reg2503 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2504 = (1'h0);
  reg [(5'h19):(1'h0)] reg2510 = (1'h0);
  reg [(5'h15):(1'h0)] reg2513 = (1'h0);
  reg [(2'h3):(1'h0)] reg2512 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2515 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2517 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2521 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2524 = (1'h0);
  reg [(3'h4):(1'h0)] reg2525 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2526 = (1'h0);
  reg [(4'hf):(1'h0)] reg2528 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2529 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2531 = (1'h0);
  reg [(5'h13):(1'h0)] reg2533 = (1'h0);
  reg [(4'hd):(1'h0)] reg2534 = (1'h0);
  reg [(4'h9):(1'h0)] reg2535 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2540 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2542 = (1'h0);
  reg [(5'h19):(1'h0)] reg2544 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2546 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2547 = (1'h0);
  reg [(3'h5):(1'h0)] reg2549 = (1'h0);
  reg [(4'he):(1'h0)] reg2551 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2552 = (1'h0);
  reg [(5'h19):(1'h0)] reg2553 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2555 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2556 = (1'h0);
  reg [(5'h10):(1'h0)] reg2557 = (1'h0);
  reg [(4'hd):(1'h0)] reg2559 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2560 = (1'h0);
  reg [(4'he):(1'h0)] reg2564 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2565 = (1'h0);
  reg [(4'h8):(1'h0)] reg2566 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2567 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2568 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2569 = (1'h0);
  reg [(5'h19):(1'h0)] reg2572 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2573 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2575 = (1'h0);
  reg [(4'hf):(1'h0)] reg2576 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2578 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2582 = (1'h0);
  reg [(3'h6):(1'h0)] reg2584 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2586 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2588 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2593 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2595 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2600 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2601 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2602 = (1'h0);
  reg [(4'ha):(1'h0)] reg2604 = (1'h0);
  reg [(5'h17):(1'h0)] reg2605 = (1'h0);
  reg [(4'hf):(1'h0)] reg2606 = (1'h0);
  reg [(4'hf):(1'h0)] reg2608 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2610 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2612 = (1'h0);
  reg [(5'h14):(1'h0)] reg2613 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2614 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2617 = (1'h0);
  reg [(5'h16):(1'h0)] reg2622 = (1'h0);
  reg [(3'h6):(1'h0)] reg2624 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2626 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2628 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2632 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2633 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2636 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2639 = (1'h0);
  reg [(4'ha):(1'h0)] reg2643 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2648 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2650 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2699 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2698 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2689 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2694 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2693 = (1'h0);
  reg [(2'h2):(1'h0)] reg2692 = (1'h0);
  reg [(5'h14):(1'h0)] reg2690 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2686 = (1'h0);
  reg [(4'hf):(1'h0)] reg2685 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2684 = (1'h0);
  reg [(4'hb):(1'h0)] reg2681 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2680 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2679 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2678 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2675 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2673 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2672 = (1'h0);
  reg [(5'h17):(1'h0)] reg2671 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2670 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2668 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2667 = (1'h0);
  reg [(4'ha):(1'h0)] reg2666 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2658 = (1'h0);
  reg [(5'h11):(1'h0)] reg2657 = (1'h0);
  reg [(4'hf):(1'h0)] reg2663 = (1'h0);
  reg [(5'h19):(1'h0)] reg2662 = (1'h0);
  reg [(4'ha):(1'h0)] reg2658 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2657 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2656 = (1'h0);
  reg [(4'h8):(1'h0)] reg2649 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2647 = (1'h0);
  reg [(5'h15):(1'h0)] reg2646 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2645 = (1'h0);
  reg [(5'h16):(1'h0)] reg2644 = (1'h0);
  reg [(2'h3):(1'h0)] reg2642 = (1'h0);
  reg [(5'h18):(1'h0)] reg2641 = (1'h0);
  reg [(4'hc):(1'h0)] reg2640 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2638 = (1'h0);
  reg [(5'h16):(1'h0)] reg2637 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar2635 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2634 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2631 = (1'h0);
  reg [(4'ha):(1'h0)] reg2630 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2629 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2627 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2625 = (1'h0);
  reg [(5'h10):(1'h0)] reg2623 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2621 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2620 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2619 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2618 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2616 = (1'h0);
  reg [(3'h6):(1'h0)] reg2615 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2606 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2611 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2609 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2607 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2603 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2599 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2598 = (1'h0);
  reg [(5'h16):(1'h0)] reg2597 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2596 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2594 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2592 = (1'h0);
  reg [(5'h16):(1'h0)] reg2591 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2590 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2589 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2587 = (1'h0);
  reg [(5'h15):(1'h0)] reg2585 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar2583 = (1'h0);
  reg [(3'h5):(1'h0)] reg2581 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2580 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2570 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2566 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2579 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2577 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2574 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2571 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2570 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2563 = (1'h0);
  reg [(5'h15):(1'h0)] reg2562 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2561 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2558 = (1'h0);
  reg [(5'h16):(1'h0)] forvar2554 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2550 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2545 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2548 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2545 = (1'h0);
  reg [(3'h6):(1'h0)] reg2543 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2541 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2539 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2538 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2537 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2536 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2532 = (1'h0);
  reg [(2'h2):(1'h0)] reg2530 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2527 = (1'h0);
  reg [(4'hb):(1'h0)] reg2523 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2522 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2520 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2519 = (1'h0);
  reg [(5'h10):(1'h0)] reg2518 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2516 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2514 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar2512 = (1'h0);
  reg [(3'h7):(1'h0)] reg2511 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2509 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2507 = (1'h0);
  reg [(3'h5):(1'h0)] reg2500 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2506 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2505 = (1'h0);
  reg [(5'h10):(1'h0)] reg2502 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2501 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2500 = (1'h0);
  reg [(4'ha):(1'h0)] reg2495 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2494 = (1'h0);
  reg [(2'h2):(1'h0)] reg2493 = (1'h0);
  reg [(3'h7):(1'h0)] reg2490 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2488 = (1'h0);
  reg [(5'h10):(1'h0)] reg2485 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2484 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2483 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2482 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2481 = (1'h0);
  reg [(3'h5):(1'h0)] reg2479 = (1'h0);
  reg [(4'hd):(1'h0)] reg2477 = (1'h0);
  reg [(4'ha):(1'h0)] reg2476 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2473 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2471 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar2470 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2469 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2467 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2465 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2464 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2462 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2457 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2456 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2460 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2457 = (1'h0);
  reg [(4'ha):(1'h0)] reg2455 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg41 = (1'h0);
  reg [(5'h1c):(1'h0)] reg40 = (1'h0);
  reg [(4'hf):(1'h0)] reg39 = (1'h0);
  reg [(5'h1e):(1'h0)] reg38 = (1'h0);
  reg [(4'hd):(1'h0)] reg37 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar35 = (1'h0);
  reg [(3'h6):(1'h0)] forvar32 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg21 = (1'h0);
  reg [(4'ha):(1'h0)] forvar20 = (1'h0);
  reg [(2'h2):(1'h0)] reg19 = (1'h0);
  reg [(5'h19):(1'h0)] forvar16 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg15 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg13 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg11 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg9 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg7 = (1'h0);
  assign y = {wire2654,
                 wire2653,
                 wire2651,
                 wire2508,
                 wire42,
                 wire2453,
                 reg2700,
                 reg2697,
                 reg2696,
                 reg2695,
                 reg2680,
                 reg2678,
                 reg2691,
                 reg2689,
                 reg2688,
                 reg2687,
                 reg2683,
                 reg2682,
                 reg2677,
                 reg2676,
                 reg2674,
                 reg2669,
                 reg2665,
                 reg2664,
                 reg2661,
                 reg2660,
                 reg2659,
                 reg5,
                 reg6,
                 reg8,
                 reg12,
                 reg17,
                 reg18,
                 reg22,
                 reg25,
                 reg27,
                 reg29,
                 reg30,
                 reg31,
                 reg33,
                 reg34,
                 reg36,
                 reg2456,
                 reg2458,
                 reg2459,
                 reg2461,
                 reg2463,
                 reg2466,
                 reg2468,
                 reg2472,
                 reg2474,
                 reg2475,
                 reg2478,
                 reg2480,
                 reg2486,
                 reg2487,
                 reg2489,
                 reg2491,
                 reg2492,
                 reg2496,
                 reg2497,
                 reg2498,
                 reg2499,
                 reg2503,
                 reg2504,
                 reg2510,
                 reg2513,
                 reg2512,
                 reg2515,
                 reg2517,
                 reg2521,
                 reg2524,
                 reg2525,
                 reg2526,
                 reg2528,
                 reg2529,
                 reg2531,
                 reg2533,
                 reg2534,
                 reg2535,
                 reg2540,
                 reg2542,
                 reg2544,
                 reg2546,
                 reg2547,
                 reg2549,
                 reg2551,
                 reg2552,
                 reg2553,
                 reg2555,
                 reg2556,
                 reg2557,
                 reg2559,
                 reg2560,
                 reg2564,
                 reg2565,
                 reg2566,
                 reg2567,
                 reg2568,
                 reg2569,
                 reg2572,
                 reg2573,
                 reg2575,
                 reg2576,
                 reg2578,
                 reg2582,
                 reg2584,
                 reg2586,
                 reg2588,
                 reg2593,
                 reg2595,
                 reg2600,
                 reg2601,
                 reg2602,
                 reg2604,
                 reg2605,
                 reg2606,
                 reg2608,
                 reg2610,
                 reg2612,
                 reg2613,
                 reg2614,
                 reg2617,
                 reg2622,
                 reg2624,
                 reg2626,
                 reg2628,
                 reg2632,
                 reg2633,
                 reg2636,
                 reg2639,
                 reg2643,
                 reg2648,
                 reg2650,
                 reg2699,
                 reg2698,
                 forvar2689,
                 reg2694,
                 reg2693,
                 reg2692,
                 reg2690,
                 reg2686,
                 reg2685,
                 reg2684,
                 reg2681,
                 forvar2680,
                 reg2679,
                 forvar2678,
                 reg2675,
                 reg2673,
                 reg2672,
                 reg2671,
                 reg2670,
                 reg2668,
                 forvar2667,
                 reg2666,
                 forvar2658,
                 reg2657,
                 reg2663,
                 reg2662,
                 reg2658,
                 forvar2657,
                 reg2656,
                 reg2649,
                 reg2647,
                 reg2646,
                 reg2645,
                 reg2644,
                 reg2642,
                 reg2641,
                 reg2640,
                 reg2638,
                 reg2637,
                 forvar2635,
                 reg2634,
                 reg2631,
                 reg2630,
                 forvar2629,
                 reg2627,
                 reg2625,
                 reg2623,
                 reg2621,
                 reg2620,
                 forvar2619,
                 reg2618,
                 forvar2616,
                 reg2615,
                 forvar2606,
                 reg2611,
                 reg2609,
                 reg2607,
                 reg2603,
                 reg2599,
                 forvar2598,
                 reg2597,
                 forvar2596,
                 reg2594,
                 reg2592,
                 reg2591,
                 reg2590,
                 reg2589,
                 reg2587,
                 reg2585,
                 forvar2583,
                 reg2581,
                 forvar2580,
                 reg2570,
                 forvar2566,
                 reg2579,
                 reg2577,
                 reg2574,
                 reg2571,
                 forvar2570,
                 reg2563,
                 reg2562,
                 reg2561,
                 reg2558,
                 forvar2554,
                 forvar2550,
                 forvar2545,
                 reg2548,
                 reg2545,
                 reg2543,
                 reg2541,
                 reg2539,
                 reg2538,
                 reg2537,
                 reg2536,
                 reg2532,
                 reg2530,
                 reg2527,
                 reg2523,
                 reg2522,
                 reg2520,
                 reg2519,
                 reg2518,
                 reg2516,
                 reg2514,
                 forvar2512,
                 reg2511,
                 reg2509,
                 reg2507,
                 reg2500,
                 reg2506,
                 reg2505,
                 reg2502,
                 reg2501,
                 forvar2500,
                 reg2495,
                 reg2494,
                 reg2493,
                 reg2490,
                 reg2488,
                 reg2485,
                 reg2484,
                 forvar2483,
                 reg2482,
                 forvar2481,
                 reg2479,
                 reg2477,
                 reg2476,
                 reg2473,
                 reg2471,
                 forvar2470,
                 reg2469,
                 forvar2467,
                 reg2465,
                 reg2464,
                 reg2462,
                 reg2457,
                 forvar2456,
                 reg2460,
                 forvar2457,
                 reg2455,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 forvar35,
                 forvar32,
                 reg28,
                 reg26,
                 reg24,
                 reg23,
                 reg21,
                 forvar20,
                 reg19,
                 forvar16,
                 reg15,
                 reg14,
                 reg13,
                 reg11,
                 reg10,
                 reg9,
                 reg7,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire3)
        begin
          if ((7'h4e))
            begin
              reg5 <= (wire1[(4'h9):(3'h4)] ~^ wire3);
              reg6 <= wire4[(4'ha):(4'h8)];
              reg7 = wire4[(1'h0):(1'h0)];
              reg8 <= (~($signed(((wire4 ? reg6 : wire0) ?
                  (wire1 == reg5) : {reg7,
                      wire0})) == $signed((reg6[(4'hd):(1'h1)] > (8'hbd)))));
              reg9 = (-$unsigned((&((~^wire4) ?
                  (-reg7) : wire3[(5'h14):(4'ha)]))));
              reg10 = reg6[(1'h1):(1'h1)];
              reg11 = $unsigned($unsigned((~^$unsigned(reg5[(3'h6):(2'h2)]))));
            end
          else
            begin
              reg7 = $signed({{reg5[(4'hc):(3'h4)],
                      (wire4 + (reg10 ? (8'hab) : (8'hbf)))},
                  wire1});
              reg8 <= ((wire2 * wire2[(3'h5):(2'h2)]) ^~ $unsigned({($unsigned(reg9) ^ {(8'hb8),
                      wire0}),
                  reg6[(5'h15):(4'h8)]}));
              reg9 = reg8[(3'h6):(2'h3)];
              reg12 <= (((^~$signed(((7'h40) & reg9))) ?
                      ($signed((reg10 <<< reg7)) * $unsigned((wire3 ?
                          wire4 : reg11))) : reg6[(5'h18):(2'h2)]) ?
                  reg11[(3'h5):(2'h2)] : ($signed({(reg8 << reg6),
                          $signed(wire4)}) ?
                      wire1[(5'h19):(4'he)] : ({(reg5 ^~ wire4)} ?
                          (~|(8'h9f)) : reg7[(4'hd):(1'h0)])));
              reg13 = reg9[(4'ha):(3'h4)];
              reg14 = (&$signed(reg10[(3'h6):(1'h0)]));
            end
          reg15 = $signed(((reg8[(5'h17):(1'h0)] ?
              (wire1 ? (|(8'hbb)) : reg9[(1'h1):(1'h0)]) : ($unsigned(wire3) ?
                  (reg9 ? wire3 : (7'h49)) : (reg9 != reg10))) <<< (wire2 ?
              $unsigned(reg11[(1'h0):(1'h0)]) : (8'ha9))));
          for (forvar16 = (1'h0); (forvar16 < (2'h2)); forvar16 = (forvar16 + (1'h1)))
            begin
              reg17 <= ($signed($signed(($unsigned(reg12) <<< {reg11,
                  reg14,
                  reg5}))) <<< reg7);
              reg18 <= {{$signed((reg13 ?
                          reg6[(4'hf):(2'h2)] : $unsigned((8'hb7))))},
                  wire1};
              reg19 = (reg7[(5'h17):(3'h6)] ?
                  $unsigned({$unsigned($signed(reg12))}) : reg6);
            end
        end
      else
        begin
          reg5 <= $unsigned($signed($signed($signed($unsigned(reg18)))));
        end
      for (forvar20 = (1'h0); (forvar20 < (3'h6)); forvar20 = (forvar20 + (1'h1)))
        begin
          reg21 = ((7'h55) || ($signed({((7'h58) ?
                  reg10 : reg9)}) && (&{reg17[(2'h3):(2'h2)]})));
        end
      reg22 <= $unsigned(((&(reg10 ?
          (reg14 ? reg19 : wire2) : $signed(reg11))) && ({{reg7}} ?
          $unsigned((reg19 - wire3)) : $unsigned((reg5 ? reg14 : reg14)))));
      reg23 = reg7[(5'h19):(4'hd)];
      if ((reg9 ?
          ($signed($signed((wire0 != wire3))) ?
              $signed(reg5) : $unsigned((7'h52))) : reg17[(5'h18):(5'h11)]))
        begin
          if ((({reg21[(3'h6):(1'h0)], $signed(reg17), reg9} ?
              $unsigned(reg8[(5'h10):(4'hb)]) : (~&(+$signed(reg21)))) < ((reg13 ?
                  $unsigned($unsigned(wire0)) : $unsigned(reg23[(4'h9):(3'h6)])) ?
              $unsigned(((~^wire3) ?
                  reg13 : $unsigned((8'ha5)))) : ($signed(wire0[(3'h4):(3'h4)]) ?
                  $unsigned(reg13[(3'h5):(1'h0)]) : $unsigned({reg15,
                      reg6,
                      reg9})))))
            begin
              reg24 = (reg23 >= reg19);
              reg25 <= ($signed(reg12[(4'h9):(3'h6)]) + $unsigned((8'h9d)));
              reg26 = reg8[(2'h3):(2'h3)];
            end
          else
            begin
              reg25 <= reg13[(1'h1):(1'h0)];
              reg26 = ($signed($unsigned(reg14[(3'h4):(1'h0)])) ?
                  $signed(reg25[(4'h8):(3'h4)]) : (forvar20 ?
                      (reg9[(3'h7):(3'h5)] ?
                          ($signed(reg12) >= $signed(reg6)) : reg24[(4'hb):(1'h1)]) : reg24));
            end
        end
      else
        begin
          reg24 = reg18;
          if (reg17[(1'h1):(1'h0)])
            begin
              reg26 = $unsigned($signed(forvar20));
            end
          else
            begin
              reg25 <= reg21[(3'h5):(1'h0)];
              reg27 <= (8'haa);
              reg28 = ((-$signed(((wire0 ? wire4 : reg18) ?
                  $unsigned(wire0) : (reg14 ? reg24 : reg24)))) || reg26);
              reg29 <= $signed((~&(($signed(reg22) + (~reg17)) ?
                  $unsigned(wire3) : reg11[(4'ha):(2'h3)])));
              reg30 <= $signed($unsigned(wire2));
            end
          reg31 <= (~^reg23);
        end
      for (forvar32 = (1'h0); (forvar32 < (3'h4)); forvar32 = (forvar32 + (1'h1)))
        begin
          reg33 <= (($signed($unsigned((|reg15))) ^~ (((-reg8) >= (reg5 >> reg25)) || $signed(((7'h4d) ?
                  reg23 : reg19)))) ?
              $unsigned(($signed((reg8 & forvar32)) >> $unsigned(reg15))) : $unsigned((-($unsigned(forvar16) ?
                  $unsigned(wire3) : (7'h42)))));
          reg34 <= $unsigned((forvar20 ?
              ((reg18 ? reg26 : reg14[(2'h3):(1'h1)]) <<< ({reg5,
                      reg18,
                      forvar20} ?
                  reg31[(2'h3):(1'h1)] : (reg23 ?
                      (8'h9e) : (7'h55)))) : $signed({(reg26 <= (7'h55))})));
        end
      for (forvar35 = (1'h0); (forvar35 < (3'h4)); forvar35 = (forvar35 + (1'h1)))
        begin
          reg36 <= ($unsigned(reg31[(3'h7):(1'h0)]) ~^ reg27[(3'h6):(2'h2)]);
          if ((reg19 ? $unsigned(reg24[(4'h9):(2'h3)]) : reg30[(4'hd):(4'h9)]))
            begin
              reg37 = reg22;
              reg38 = ((&(7'h4b)) >= ((+$signed((reg27 ?
                  (7'h49) : forvar16))) << (reg18 ?
                  reg19 : $signed({reg28, reg14}))));
              reg39 = $signed($signed(reg27));
              reg40 = {$unsigned(((+$signed((8'hb9))) ?
                      (reg11 ? (wire3 ? reg37 : wire3) : reg19) : ((~&(8'hbd)) ?
                          reg31[(3'h7):(3'h7)] : {forvar32}))),
                  reg34};
            end
          else
            begin
              reg37 = (reg17[(5'h12):(3'h4)] ?
                  $unsigned(reg24[(4'h8):(3'h7)]) : $unsigned($unsigned(reg14)));
            end
        end
    end
  always
    @(posedge clk) begin
      reg41 = {reg25[(5'h18):(4'hc)],
          (((-(reg34 && wire3)) << ($unsigned(reg31) - $unsigned(wire2))) ?
              (^~((reg25 << reg12) < (^reg17))) : (~^$signed((reg33 | reg25)))),
          ((!(reg17 ?
              (wire3 - reg29) : (wire3 ?
                  reg30 : reg12))) >>> ($unsigned((reg34 ? (7'h58) : reg30)) ?
              (+(^reg29)) : ({reg12, (8'had), reg22} >= $signed(reg8))))};
    end
  assign wire42 = ((&((!$unsigned(reg31)) > (((7'h50) ~^ reg33) | ((7'h4e) >> reg34)))) ^~ ($signed((~^(reg17 ?
                          reg31 : reg33))) ?
                      reg34[(1'h1):(1'h0)] : reg22));
  module43 #() modinst2454 (wire2453, clk, reg36, reg27, reg31, reg5, wire3);
  always
    @(posedge clk) begin
      reg2455 = {{(^~wire2[(3'h4):(3'h4)]),
              $unsigned((|(reg5 ? (7'h49) : wire0)))},
          (~&(({reg22, reg17} >>> ((8'ha5) ? (7'h4c) : (7'h51))) ?
              $unsigned(reg17[(4'hb):(4'h8)]) : (8'hbd))),
          (reg33[(1'h0):(1'h0)] ^ (~&$signed(reg8[(5'h11):(4'ha)])))};
      if (($unsigned((!($unsigned((7'h53)) ?
          {reg34} : $signed((8'hbf))))) + (!reg2455)))
        begin
          reg2456 <= ($unsigned($unsigned((|reg18[(4'h9):(4'h8)]))) >>> ((~^($unsigned((8'ha1)) ~^ $signed(reg30))) ?
              ((wire2453[(3'h5):(1'h0)] ? $unsigned(wire2453) : (-reg31)) ?
                  reg36[(4'hf):(4'h9)] : ($unsigned(wire1) ?
                      (wire3 & wire2) : $signed((7'h49)))) : $unsigned($signed($unsigned((8'ha2))))));
          for (forvar2457 = (1'h0); (forvar2457 < (1'h0)); forvar2457 = (forvar2457 + (1'h1)))
            begin
              reg2458 <= reg33[(3'h6):(3'h4)];
              reg2459 <= $signed($unsigned((&wire2[(3'h6):(1'h0)])));
              reg2460 = {{((~|(wire0 ?
                          reg8 : reg33)) << (((7'h43) >>> wire3) || $signed(reg5))),
                      (wire3[(3'h6):(1'h1)] << ($signed(wire2) < (wire0 ?
                          reg36 : reg33))),
                      (((8'hb1) ?
                          $unsigned(reg5) : (reg36 < reg30)) > $signed($signed(reg22)))}};
            end
        end
      else
        begin
          for (forvar2456 = (1'h0); (forvar2456 < (1'h1)); forvar2456 = (forvar2456 + (1'h1)))
            begin
              reg2457 = (8'hba);
              reg2460 = reg31[(2'h3):(1'h0)];
              reg2461 <= (reg29 + $signed({(reg2458[(2'h2):(2'h2)] >> $unsigned((8'hb9))),
                  (wire42 >>> {reg12}),
                  reg5[(3'h4):(1'h0)]}));
            end
          if ((($signed(wire4) ?
                  $signed(reg34[(2'h3):(1'h1)]) : ($unsigned((wire3 ^ reg22)) ?
                      $signed((^reg2456)) : ($unsigned((8'hba)) ?
                          reg33 : {forvar2456, reg25, forvar2456}))) ?
              $signed($unsigned((reg2458 & $unsigned(reg6)))) : $unsigned((^(!$signed(reg27))))))
            begin
              reg2462 = ((8'ha7) ?
                  ((~{{reg5, reg25, wire1},
                      reg30[(4'ha):(3'h4)]}) || wire2) : $signed($unsigned($signed(((7'h4d) ?
                      reg2456 : (8'h9e))))));
              reg2463 <= (reg29 ?
                  ($unsigned($signed($unsigned(reg34))) >>> reg5[(2'h3):(2'h3)]) : $signed($unsigned($signed($unsigned(reg2461)))));
              reg2464 = (reg2456 ?
                  reg34[(1'h0):(1'h0)] : (($signed($signed(wire4)) != {(~(8'ha9)),
                      (reg18 == reg29),
                      (reg29 + reg31)}) > wire4));
              reg2465 = (+($signed(($unsigned(reg33) != reg36)) >> $signed($signed((wire2453 == reg31)))));
            end
          else
            begin
              reg2462 = (|reg2460[(3'h7):(3'h6)]);
            end
          reg2466 <= (~((+(!reg34)) || reg5[(3'h5):(1'h0)]));
          for (forvar2467 = (1'h0); (forvar2467 < (2'h3)); forvar2467 = (forvar2467 + (1'h1)))
            begin
              reg2468 <= (~|reg29);
              reg2469 = reg8;
            end
        end
      for (forvar2470 = (1'h0); (forvar2470 < (2'h2)); forvar2470 = (forvar2470 + (1'h1)))
        begin
          reg2471 = wire1;
          reg2472 <= $signed((forvar2457[(5'h10):(4'hc)] >> (reg2465[(3'h6):(1'h0)] > reg2468)));
          reg2473 = reg2465[(4'ha):(4'h8)];
          if (reg2463[(5'h1a):(5'h19)])
            begin
              reg2474 <= reg18;
              reg2475 <= {(forvar2456 ?
                      forvar2456 : $signed({(^~reg18), {reg36}, wire2453}))};
              reg2476 = (($signed(({wire4} >>> $signed(reg5))) ^~ $unsigned({reg29[(4'hf):(2'h2)]})) || $signed($signed(reg8)));
              reg2477 = reg2469[(5'h1b):(5'h16)];
              reg2478 <= ((((((8'hbf) ? reg12 : (7'h54)) ?
                          $unsigned(reg29) : $unsigned(wire4)) <= reg2475) ?
                      (wire2[(3'h4):(1'h1)] ?
                          (~&(reg34 ?
                              reg2477 : forvar2467)) : ($unsigned(reg33) ^~ reg2457[(1'h0):(1'h0)])) : (^($unsigned(forvar2470) ?
                          (~|forvar2456) : {reg2458, reg2463, reg2469}))) ?
                  (reg2466[(5'h15):(3'h6)] != ($unsigned(wire1) ?
                      ($unsigned((8'h9e)) <<< reg2473) : (~reg29))) : ((|$signed((reg2466 ^ reg2463))) << ($signed($signed((8'hb7))) ?
                      (^(wire42 ?
                          reg36 : reg27)) : ((wire42 < wire0) >> (reg25 >= (8'h9c))))));
              reg2479 = reg2464;
            end
          else
            begin
              reg2474 <= {((~^(forvar2470[(4'hc):(3'h7)] > $unsigned(reg29))) ?
                      $signed(($signed(wire4) != (~^wire2453))) : (-reg2462))};
              reg2476 = $signed((($unsigned((reg2458 <<< (7'h4b))) ?
                      ((^~reg17) & {reg34}) : (~|(reg2478 ?
                          (8'haf) : (8'hb8)))) ?
                  (reg31 + ($unsigned(reg5) && $unsigned(wire3))) : reg2457[(2'h2):(1'h1)]));
              reg2478 <= reg2462[(4'hf):(3'h5)];
              reg2480 <= $signed($unsigned($signed(wire3)));
            end
          for (forvar2481 = (1'h0); (forvar2481 < (1'h1)); forvar2481 = (forvar2481 + (1'h1)))
            begin
              reg2482 = $signed(reg2469[(4'hc):(1'h1)]);
            end
          for (forvar2483 = (1'h0); (forvar2483 < (3'h4)); forvar2483 = (forvar2483 + (1'h1)))
            begin
              reg2484 = $unsigned(((({forvar2456,
                      reg2455} >>> reg2477[(1'h1):(1'h0)]) ?
                  reg18 : $unsigned({reg2468,
                      reg31,
                      forvar2456})) & ((7'h51) || reg2466[(5'h15):(4'h9)])));
              reg2485 = (8'ha1);
              reg2486 <= $unsigned(($unsigned(((~^reg2474) << (8'hb3))) == ({$unsigned((7'h56)),
                  reg2485,
                  $signed((7'h48))} | ($signed(reg27) ?
                  $signed(reg2478) : {reg2482}))));
              reg2487 <= (((^~reg2479) ?
                  reg2461 : reg27[(4'hc):(4'h8)]) ^~ $signed((reg2456 - ((wire42 >> wire4) ?
                  (reg6 && (7'h46)) : {reg8}))));
            end
        end
      if (($unsigned((~&$signed({(8'hb6),
          reg2466}))) << ((~^$signed(((7'h49) ^ reg2462))) != (^~forvar2483[(3'h7):(2'h3)]))))
        begin
          reg2488 = wire0[(2'h2):(2'h2)];
          if (reg25[(5'h1e):(5'h1c)])
            begin
              reg2489 <= (($signed((|(^(8'ha2)))) ?
                      $signed({(8'hb2),
                          {reg2473}}) : {(-(forvar2457 * (8'hba))),
                          (reg31[(3'h4):(2'h2)] ?
                              (^reg2477) : (reg2471 - reg2485)),
                          wire2453}) ?
                  (~(reg2487 ~^ ($signed(reg2468) ?
                      $signed((8'hab)) : reg2461[(1'h0):(1'h0)]))) : $signed(((!(~reg2456)) ?
                      ((reg2486 ^ reg30) << {(8'ha8),
                          reg2458,
                          reg22}) : ((reg2459 ? forvar2470 : reg2463) ?
                          (&(8'hbe)) : reg2463))));
              reg2490 = forvar2483;
              reg2491 <= reg2488[(4'h8):(1'h0)];
              reg2492 <= reg18;
            end
          else
            begin
              reg2490 = reg2482;
              reg2493 = (^(-((~&(~&reg2468)) ?
                  ((+reg2456) <<< $signed(wire2453)) : $unsigned($signed(reg29)))));
              reg2494 = (!reg12);
              reg2495 = ((forvar2481[(1'h1):(1'h1)] ?
                      (-(wire3[(4'he):(3'h5)] ?
                          {reg6,
                              (8'ha5),
                              reg2462} : (^forvar2481))) : (reg17[(3'h7):(3'h5)] ~^ forvar2467[(3'h7):(3'h5)])) ?
                  ($signed(reg2485[(3'h4):(1'h0)]) ?
                      {$signed($signed(reg2475))} : (~&reg2476)) : ((~&$unsigned($signed((8'hbb)))) ^~ ($signed(((8'h9f) <<< (7'h52))) >= (((7'h4b) ?
                      reg2482 : reg2472) | ((8'hac) << reg2476)))));
              reg2496 <= ($signed((^~($unsigned(reg2491) ?
                  (~|reg2479) : (~|reg25)))) <= ($signed($unsigned($signed(reg2460))) ?
                  $signed(((|reg34) ?
                      $signed(reg2494) : (!wire42))) : $signed((~|(reg2461 ?
                      reg2474 : reg8)))));
              reg2497 <= (|$unsigned(reg2484));
              reg2498 <= $unsigned((reg2486 ?
                  ((^~reg2495) ?
                      (reg2462 >= {wire0,
                          reg2466,
                          reg2493}) : $unsigned((~reg6))) : (7'h50)));
            end
          reg2499 <= (^~$signed(reg2488[(2'h2):(1'h1)]));
          for (forvar2500 = (1'h0); (forvar2500 < (2'h3)); forvar2500 = (forvar2500 + (1'h1)))
            begin
              reg2501 = $signed($unsigned((+(~^(-reg2479)))));
              reg2502 = $signed((reg2494[(4'ha):(2'h3)] ?
                  forvar2456 : (reg2501 ? reg2460 : $signed((8'hb6)))));
              reg2503 <= wire3;
              reg2504 <= ({{($signed(reg18) ? (!forvar2470) : reg22),
                          reg2493,
                          $signed(((8'h9e) ? wire3 : reg29))}} ?
                  reg2490[(3'h4):(1'h0)] : reg2495[(1'h1):(1'h0)]);
              reg2505 = wire2[(3'h7):(3'h4)];
              reg2506 = $unsigned(wire2);
            end
        end
      else
        begin
          if ((~^$signed((|{(+reg18), reg2499}))))
            begin
              reg2488 = ($unsigned(($signed((reg2492 ? reg2479 : reg2480)) ?
                      $signed((reg2487 ^ reg2466)) : $unsigned((~|reg2496)))) ?
                  (~|$signed($signed((reg2466 >= wire2453)))) : (!(|wire42[(3'h6):(1'h0)])));
              reg2490 = reg2498;
              reg2491 <= {((-$unsigned((reg2473 <= reg2464))) ?
                      (+reg12[(3'h7):(3'h5)]) : ((7'h43) <= {reg2505})),
                  ($signed((^$signed(wire2453))) ^~ ($unsigned({(8'hb5),
                          forvar2500}) ?
                      $unsigned(reg2464) : ({reg2457} ?
                          $unsigned(reg2463) : $unsigned((8'ha5)))))};
              reg2492 <= (|($unsigned($signed((reg2487 ?
                  reg2499 : reg2477))) ^~ $unsigned($unsigned((reg2473 ~^ wire2453)))));
            end
          else
            begin
              reg2488 = $signed($signed((8'hb1)));
              reg2489 <= $signed(($unsigned($unsigned((reg34 >>> (7'h41)))) && (-$unsigned($signed(reg2473)))));
              reg2491 <= ($signed({((reg2501 << wire0) && reg12),
                      (~&(~&(8'had)))}) ?
                  $signed(((reg2491[(4'he):(4'h8)] || ((8'hbd) || wire0)) ?
                      reg2476 : ((reg2496 ? (8'hbf) : reg2457) ?
                          (reg2496 ?
                              reg2505 : reg2480) : (&reg2455)))) : {(^{(8'ha8),
                          $unsigned(reg2462)}),
                      (reg2477[(3'h6):(3'h5)] << {wire2453,
                          (~^reg2497),
                          (reg2502 ? (7'h51) : wire3)}),
                      wire1[(5'h18):(1'h1)]});
              reg2493 = (-(^~$signed(forvar2456)));
              reg2494 = {(reg31[(5'h15):(4'h8)] ?
                      (!$signed({forvar2481,
                          (7'h4c),
                          reg2486})) : reg18[(4'he):(3'h4)]),
                  $unsigned($signed($signed(reg2496[(3'h5):(1'h1)])))};
              reg2495 = $unsigned((^(+({reg2477, reg22, forvar2483} ?
                  $signed(reg2456) : (reg2503 ? (7'h58) : reg2475)))));
            end
          reg2496 <= reg2458[(5'h12):(4'he)];
          if ((reg2497 <<< reg2477))
            begin
              reg2497 <= (((-reg2476[(4'h9):(3'h5)]) ?
                      reg36 : reg2487[(5'h1a):(5'h1a)]) ?
                  $unsigned($unsigned($unsigned((|reg2503)))) : (reg2486 ?
                      forvar2500[(4'h9):(1'h0)] : forvar2467));
              reg2500 = reg27[(1'h1):(1'h0)];
            end
          else
            begin
              reg2500 = reg2492;
              reg2501 = {(^(^$signed((wire0 == reg2497)))),
                  (({$unsigned(reg2498)} ?
                          ((reg2491 - wire0) < reg18[(4'hf):(2'h3)]) : ((~|reg2484) >> reg31)) ?
                      ((reg2473 ? reg34 : reg25) ?
                          $signed((reg2469 > reg2502)) : {(~^reg17),
                              (wire1 ? reg2463 : reg6)}) : (^((reg2499 ?
                          reg2466 : reg2474) << (+wire2)))),
                  reg2472};
              reg2502 = ($unsigned({(reg30 ?
                          $unsigned(reg5) : {(8'ha8), reg2487, reg2466}),
                      $signed(reg2475),
                      $unsigned(wire2)}) ?
                  reg2498 : ({reg2499,
                      (!(reg33 ? reg2488 : reg2465))} > reg2497));
            end
          reg2505 = (reg2474 ?
              ((reg33[(4'he):(4'hb)] >> $unsigned($unsigned(reg2461))) << wire0) : (&$signed((~^forvar2470))));
          reg2506 = $signed($unsigned($unsigned((^~forvar2467[(3'h5):(1'h1)]))));
        end
      reg2507 = $signed($unsigned(reg2464[(1'h1):(1'h1)]));
    end
  assign wire2508 = $signed(((reg2486[(1'h0):(1'h0)] ?
                        ((8'ha4) * (|reg5)) : (wire2 + (8'h9d))) <= reg2472[(3'h4):(2'h2)]));
  always
    @(posedge clk) begin
      reg2509 = (|reg2456);
      if ((^~(~^{$signed(reg22[(4'hc):(4'h8)]), $signed((^~reg2504))})))
        begin
          reg2510 <= (((-(-{reg2498, reg2496, (8'ha1)})) ?
              $signed(reg2474) : $unsigned((+reg2496))) >= $unsigned(reg2496));
          reg2511 = $signed(reg2463[(2'h3):(2'h2)]);
          for (forvar2512 = (1'h0); (forvar2512 < (3'h4)); forvar2512 = (forvar2512 + (1'h1)))
            begin
              reg2513 <= reg2511;
              reg2514 = reg2478;
            end
        end
      else
        begin
          reg2511 = (($signed($unsigned($signed(reg17))) ?
              ((((8'h9f) ?
                  (8'hbb) : reg2486) << $unsigned((7'h4f))) >> reg30[(4'h9):(3'h6)]) : ($signed((reg2456 ?
                      reg2463 : reg2474)) ?
                  ((wire3 ?
                      (8'hb8) : reg2514) <<< $signed(reg2461)) : ((~&(8'hbb)) | (~^wire1)))) ~^ (reg25[(5'h1f):(4'h8)] ?
              $unsigned($unsigned((reg2497 ~^ reg8))) : reg2503));
          if ($signed(($unsigned(((|(8'hb1)) ?
                  $unsigned((8'hba)) : reg5[(5'h15):(5'h14)])) ?
              {reg2504,
                  $signed((reg2510 || reg2503))} : (((reg2468 == reg31) && reg22[(1'h0):(1'h0)]) ?
                  reg2478[(5'h14):(5'h13)] : (&$signed(reg29))))))
            begin
              reg2512 <= reg2504[(4'h9):(3'h4)];
              reg2513 <= reg2466[(5'h11):(2'h2)];
              reg2514 = (^~$unsigned(reg2474[(2'h2):(1'h1)]));
              reg2515 <= $signed((wire42[(4'h8):(4'h8)] * $signed(reg2503[(4'hc):(2'h3)])));
              reg2516 = $signed(((reg2474[(3'h4):(2'h2)] | reg31) | (($unsigned(reg2466) > wire1[(5'h18):(5'h13)]) > (~$unsigned(reg2486)))));
              reg2517 <= (-(7'h46));
            end
          else
            begin
              reg2514 = (7'h48);
              reg2515 <= $unsigned(reg12);
              reg2516 = ($unsigned($unsigned(reg2458)) ?
                  ($signed((~^$unsigned(reg5))) <<< $unsigned($unsigned({reg2456,
                      reg6,
                      reg29}))) : wire2453);
              reg2517 <= (((reg2458 ?
                  $signed(reg29[(4'hd):(3'h6)]) : ((reg2461 ?
                          reg2486 : reg2475) ?
                      (reg2492 ?
                          reg2456 : reg2511) : $signed(reg17))) - reg5) <<< $unsigned((reg2458[(4'h8):(1'h0)] & $unsigned((reg2487 ?
                  reg2517 : reg5)))));
            end
        end
      if ($unsigned(((~&(|reg2461)) ?
          reg2486 : {$signed((-wire2)),
              ({reg2459, forvar2512} ?
                  $signed(reg2463) : (wire1 ? reg2499 : wire0))})))
        begin
          reg2518 = $signed(reg2468[(4'hc):(2'h2)]);
        end
      else
        begin
          if (reg2498)
            begin
              reg2518 = {reg2463};
            end
          else
            begin
              reg2518 = $signed((8'hb0));
              reg2519 = reg2515[(2'h2):(1'h1)];
              reg2520 = reg2509[(3'h6):(3'h6)];
              reg2521 <= wire42[(3'h5):(3'h4)];
              reg2522 = ((reg2504[(3'h4):(3'h4)] ?
                  wire4 : (&$unsigned(reg2459))) + {$unsigned((^~reg2513[(4'hb):(4'h8)]))});
              reg2523 = $signed($unsigned($unsigned(({(8'h9d),
                  reg2478} >= reg31))));
            end
          if (($signed({(8'ha6)}) | $unsigned($signed($signed({reg2486,
              reg6,
              reg2523})))))
            begin
              reg2524 <= (reg33 <= $unsigned(reg34[(1'h1):(1'h0)]));
              reg2525 <= $signed(($unsigned(wire3[(2'h2):(2'h2)]) ?
                  reg2513[(3'h6):(3'h4)] : (7'h57)));
              reg2526 <= (&(({{reg31}, reg2524, (reg33 ? (8'h9d) : reg2521)} ?
                      (~&reg25[(2'h3):(1'h0)]) : reg2503[(5'h10):(4'ha)]) ?
                  ($unsigned(reg2461[(3'h4):(2'h3)]) ?
                      ({(8'ha0)} ?
                          reg2497[(2'h2):(1'h1)] : (~wire2453)) : ($signed(reg18) != $signed(reg2504))) : $signed(((7'h46) | (+reg2510)))));
            end
          else
            begin
              reg2527 = reg2524;
              reg2528 <= reg25[(1'h1):(1'h1)];
              reg2529 <= reg2518[(4'he):(4'hb)];
              reg2530 = (^$signed({(reg2518[(3'h7):(1'h0)] + (^reg2529))}));
              reg2531 <= $unsigned(reg2510);
              reg2532 = {$unsigned(reg27[(2'h3):(2'h2)])};
            end
          if ($unsigned({(8'hbc)}))
            begin
              reg2533 <= ($signed((^~($unsigned(reg2510) ?
                  (reg27 < reg2491) : (reg2513 * reg36)))) + wire2508);
              reg2534 <= (~|($unsigned($signed({reg2531, (8'ha0), reg2530})) ?
                  reg2531[(3'h4):(3'h4)] : $unsigned((reg17[(3'h7):(1'h1)] ?
                      $signed(reg2478) : reg2512))));
              reg2535 <= $signed((reg17[(5'h17):(5'h14)] ?
                  $unsigned((^~(^~reg2503))) : reg2525));
            end
          else
            begin
              reg2533 <= ((((|{reg2459,
                      reg2513,
                      reg18}) ^~ $signed($unsigned(reg2529))) ^ (-$unsigned((reg2528 ?
                      reg2532 : reg2529)))) ?
                  (-((reg2531 ^~ $signed(reg2480)) ?
                      $signed((reg2514 ?
                          wire2508 : (7'h51))) : reg2535)) : $signed({$unsigned((reg2474 >> reg2456))}));
              reg2534 <= reg2475[(3'h4):(3'h4)];
              reg2535 <= ((&reg2522) ~^ reg22);
              reg2536 = wire1[(4'hf):(3'h4)];
              reg2537 = {reg2474};
              reg2538 = {reg12[(4'he):(4'hd)],
                  $unsigned($signed((~reg2474[(3'h4):(2'h2)]))),
                  ({{reg2511}} ?
                      (+(^{reg31, reg2497, wire42})) : (reg2496[(4'h9):(2'h3)] ?
                          $unsigned(reg2478) : reg2520))};
              reg2539 = ($unsigned($unsigned($unsigned((reg2509 ?
                      (7'h4a) : reg2530)))) ?
                  ((~|wire1[(5'h1c):(3'h5)]) ?
                      $unsigned((7'h4e)) : reg2525) : $signed($signed(($unsigned(reg2504) ?
                      (!reg2513) : {wire2508}))));
            end
        end
      reg2540 <= (reg25 ?
          {(((reg2497 != wire2) == $signed(reg2492)) >>> (~(reg2512 >= reg2528)))} : (+(+(~$unsigned(reg2530)))));
      reg2541 = (reg2498 + (wire2453[(3'h5):(2'h3)] ?
          ($unsigned((reg34 ?
              reg2478 : reg2458)) && (+$signed((8'ha7)))) : reg2504));
    end
  always
    @(posedge clk) begin
      if ($unsigned((reg2510 << (reg2496[(3'h7):(3'h4)] >= {(reg2499 ?
              reg2466 : reg2503),
          (&reg2512),
          $unsigned(reg2517)}))))
        begin
          if (((^(&$signed({reg2517}))) ^ reg17[(4'hd):(1'h1)]))
            begin
              reg2542 <= (+$unsigned((~((~|reg22) + (~(8'hbb))))));
            end
          else
            begin
              reg2543 = $signed((reg2456 ?
                  ($unsigned(reg2489) ?
                      {$unsigned(wire2453),
                          $unsigned(reg33)} : (reg34 > (8'h9d))) : (~&reg2491[(3'h7):(2'h3)])));
              reg2544 <= ({{(~(reg2504 ? reg27 : reg2459)),
                          $unsigned((reg2497 >>> (8'hab)))},
                      ({reg2504} ?
                          ((reg25 ? reg2498 : reg5) ?
                              reg31 : ((8'ha9) ^ wire2)) : (((8'ha4) ?
                              reg17 : reg8) * $signed(reg22))),
                      wire0[(1'h0):(1'h0)]} ?
                  reg34 : (!reg2504));
              reg2545 = $unsigned({$unsigned((~$signed(reg2474)))});
              reg2546 <= (reg2543[(3'h6):(3'h5)] ?
                  ((reg2461 ?
                      (^reg2491[(3'h5):(3'h5)]) : (~|(reg2468 ?
                          reg2544 : reg2491))) * reg2524[(3'h7):(3'h7)]) : reg2512[(1'h0):(1'h0)]);
              reg2547 <= $unsigned($signed((~&((~&(7'h55)) ?
                  $signed((8'hb3)) : $signed((7'h58))))));
              reg2548 = $signed((|($unsigned(reg2480[(4'hd):(4'hd)]) ?
                  {(reg8 || (7'h4f))} : reg2496[(3'h7):(1'h0)])));
              reg2549 <= reg2533[(3'h5):(1'h0)];
            end
        end
      else
        begin
          if ($unsigned((~|reg2499[(1'h0):(1'h0)])))
            begin
              reg2543 = (~|($unsigned(((~&reg27) ^ $signed(reg5))) | $signed($unsigned($unsigned(reg34)))));
            end
          else
            begin
              reg2543 = ($signed(reg2486) ? $signed(wire3) : (7'h4e));
              reg2544 <= reg2512;
            end
          for (forvar2545 = (1'h0); (forvar2545 < (3'h5)); forvar2545 = (forvar2545 + (1'h1)))
            begin
              reg2546 <= $unsigned($unsigned({($unsigned(reg2468) != (~^reg2524)),
                  (reg2533 ? $signed(reg5) : reg2478[(4'hc):(2'h2)]),
                  reg2531[(4'hd):(4'hb)]}));
            end
          reg2547 <= ($unsigned((reg33 + $unsigned($unsigned((8'hb0))))) << {{(reg2496[(4'h8):(4'h8)] + (reg29 ?
                      reg29 : reg2461))},
              reg27,
              ((~$signed(reg2529)) ?
                  reg2486[(3'h7):(3'h4)] : ((reg22 ~^ reg2512) ?
                      (reg2489 & reg2525) : $signed(wire2)))});
          reg2548 = $signed(reg2472[(4'h9):(2'h3)]);
          reg2549 <= wire2;
          for (forvar2550 = (1'h0); (forvar2550 < (2'h3)); forvar2550 = (forvar2550 + (1'h1)))
            begin
              reg2551 <= $unsigned(($signed((|(~reg2548))) >= ((~|((7'h4d) ?
                  reg2492 : (8'hbe))) - reg18)));
              reg2552 <= wire2508;
            end
        end
      reg2553 <= (~|($signed((+(reg2463 ^~ reg2466))) ^ (+(8'ha5))));
      if (wire3[(4'he):(4'ha)])
        begin
          for (forvar2554 = (1'h0); (forvar2554 < (1'h1)); forvar2554 = (forvar2554 + (1'h1)))
            begin
              reg2555 <= reg27;
              reg2556 <= $unsigned(((~^($unsigned(reg33) >= (reg2478 ^~ reg2504))) != $signed($unsigned((&reg2472)))));
              reg2557 <= ({{reg2528[(3'h5):(1'h0)],
                      wire0[(2'h2):(1'h0)],
                      reg2546[(4'hd):(1'h1)]}} >= ($unsigned(reg2526) | $signed(reg12[(4'hd):(4'hb)])));
              reg2558 = (reg2456 ?
                  $unsigned($signed($signed((reg2533 && (7'h44))))) : $signed(((reg2543 ^~ reg2499) ?
                      (8'hae) : $signed((reg2544 == (7'h51))))));
              reg2559 <= (-{$unsigned($unsigned(reg2480)),
                  $signed((|(forvar2550 ? wire0 : reg2486)))});
              reg2560 <= $unsigned(reg2510);
              reg2561 = (reg2474[(1'h0):(1'h0)] ?
                  {(((reg18 ?
                          reg2498 : reg2474) ^~ (reg2475 + reg6)) != reg2474)} : (~{((reg2543 == wire0) >> reg2510[(2'h3):(1'h1)])}));
            end
          if ({$signed((^(((8'hb5) == reg5) - {wire2453, reg6, reg2491})))})
            begin
              reg2562 = (&$signed($unsigned($unsigned({reg2525}))));
              reg2563 = $unsigned((reg2456[(5'h16):(4'h9)] ?
                  $signed(($signed(reg2480) == $signed(reg2487))) : ($signed(reg2533[(5'h10):(4'h8)]) ?
                      $unsigned((reg25 ?
                          reg31 : reg8)) : {reg2544[(5'h17):(1'h0)],
                          ((8'hbf) ? reg2486 : reg6)})));
              reg2564 <= $signed(reg2547);
            end
          else
            begin
              reg2564 <= $unsigned((({reg34[(1'h1):(1'h1)],
                  reg2563[(5'h13):(4'h8)],
                  {reg2512}} == $signed(reg2564[(4'hd):(4'ha)])) - $unsigned(((!(8'hb1)) ?
                  (reg2526 ? wire42 : reg2542) : $signed(reg2474)))));
              reg2565 <= $unsigned((+reg2472[(2'h2):(1'h1)]));
              reg2566 <= (reg2496[(2'h3):(2'h3)] ?
                  ({(^~(&reg29))} ?
                      ((7'h52) ?
                          {$signed((8'hb4)),
                              $unsigned(reg2512),
                              $signed((7'h55))} : $unsigned({reg2526,
                              reg2486})) : (reg2564 - reg2533[(2'h2):(2'h2)])) : reg8[(4'hc):(1'h0)]);
              reg2567 <= $unsigned(($unsigned(reg2487) ?
                  (reg2486 ^ ({reg2551,
                      wire1,
                      reg2498} + $signed(wire3))) : reg29[(4'hd):(4'hb)]));
              reg2568 <= $unsigned((forvar2550 < reg2503[(5'h10):(4'hd)]));
              reg2569 <= $unsigned(reg2556[(3'h5):(3'h5)]);
            end
          for (forvar2570 = (1'h0); (forvar2570 < (2'h2)); forvar2570 = (forvar2570 + (1'h1)))
            begin
              reg2571 = (|{(^$unsigned((reg2486 ? reg2561 : reg2564)))});
              reg2572 <= $signed($signed(($signed((reg2559 + reg2543)) ?
                  $unsigned($unsigned(reg2491)) : $signed((reg2566 ?
                      reg2503 : (7'h56))))));
              reg2573 <= $signed((((((8'ha8) ? (8'hb6) : reg2555) <<< reg31) ?
                  {((7'h4a) || wire2),
                      reg2526,
                      reg2521[(5'h11):(3'h5)]} : $unsigned(reg2528[(4'h9):(3'h5)])) == $unsigned($unsigned((reg2472 == reg2492)))));
              reg2574 = $signed((~|$signed(wire4[(4'he):(4'he)])));
              reg2575 <= (reg2468 && reg2548);
              reg2576 <= $unsigned((7'h44));
            end
          reg2577 = reg2540;
          reg2578 <= reg2547[(3'h7):(3'h6)];
          reg2579 = reg2552[(3'h4):(1'h1)];
        end
      else
        begin
          for (forvar2554 = (1'h0); (forvar2554 < (3'h6)); forvar2554 = (forvar2554 + (1'h1)))
            begin
              reg2555 <= reg2571[(2'h3):(2'h3)];
              reg2558 = ({(&forvar2554),
                      (reg2577 || {wire2508}),
                      $signed((7'h49))} ?
                  $signed($unsigned((reg2548 ?
                      reg2504[(1'h0):(1'h0)] : reg2578[(1'h1):(1'h0)]))) : ($signed((reg2491[(4'hf):(4'ha)] ?
                      reg2512 : reg2503[(4'h8):(1'h0)])) > (!($unsigned(reg2489) <<< $signed(reg2459)))));
              reg2559 <= {$unsigned($unsigned(forvar2545[(4'hc):(4'ha)])),
                  (^~reg17),
                  $unsigned($unsigned($unsigned(reg2574)))};
              reg2560 <= $unsigned((~|$signed({$unsigned(reg2535), (|reg5)})));
              reg2564 <= $unsigned(reg2560[(3'h6):(3'h6)]);
              reg2565 <= reg2556[(2'h3):(1'h1)];
            end
          for (forvar2566 = (1'h0); (forvar2566 < (1'h0)); forvar2566 = (forvar2566 + (1'h1)))
            begin
              reg2570 = reg2531;
              reg2572 <= reg22[(1'h1):(1'h0)];
              reg2573 <= $signed(reg2499[(5'h13):(3'h6)]);
              reg2574 = (reg2496[(1'h0):(1'h0)] - (^~$unsigned((reg25 ?
                  (reg5 != reg2472) : $signed(reg2543)))));
              reg2575 <= (-{(reg2577[(1'h1):(1'h0)] == $unsigned($signed(reg2547)))});
              reg2577 = $unsigned((^((^~reg25) ^ reg2557)));
              reg2579 = reg18;
            end
          for (forvar2580 = (1'h0); (forvar2580 < (3'h6)); forvar2580 = (forvar2580 + (1'h1)))
            begin
              reg2581 = (reg2461[(4'h8):(4'h8)] ? wire2 : reg2563);
              reg2582 <= (((^~(&(~(8'hb4)))) << reg2525[(1'h0):(1'h0)]) ?
                  ((reg2559 > (reg5[(5'h13):(4'h8)] << (reg6 && reg2496))) ?
                      $unsigned($unsigned($signed((8'ha8)))) : (reg2567[(3'h5):(3'h5)] ?
                          reg36 : $signed((reg2560 ?
                              reg25 : (7'h4f))))) : (({(reg2531 <= reg2531)} ?
                      $signed((reg2472 | reg2544)) : ({reg2487} - $signed(reg2568))) * wire2508));
            end
          for (forvar2583 = (1'h0); (forvar2583 < (2'h2)); forvar2583 = (forvar2583 + (1'h1)))
            begin
              reg2584 <= wire3[(5'h19):(4'h8)];
              reg2585 = $signed(reg2475[(2'h3):(1'h1)]);
              reg2586 <= ((^~wire2508) ?
                  {$unsigned(reg2556[(1'h0):(1'h0)]),
                      (^(reg2555 < (reg2552 ? reg2472 : (7'h54)))),
                      $unsigned(($signed(reg2568) * (~&wire4)))} : $signed((^~({reg2560,
                      reg2468,
                      reg2577} ^ $unsigned(reg2458)))));
              reg2587 = reg2569[(4'hd):(1'h0)];
              reg2588 <= reg2555[(3'h4):(1'h1)];
              reg2589 = $unsigned($signed($unsigned(reg30)));
            end
          if (({($signed((reg27 ?
                  reg2525 : wire3)) >> $signed((^~reg2547)))} <= reg2459))
            begin
              reg2590 = reg2531[(4'hd):(2'h3)];
            end
          else
            begin
              reg2590 = $unsigned($unsigned(reg31[(4'hf):(4'h9)]));
              reg2591 = $unsigned((^((reg2510 ?
                  $unsigned(reg2558) : $signed(reg2531)) >> (~reg2565[(3'h4):(1'h1)]))));
              reg2592 = reg2555[(2'h2):(1'h0)];
              reg2593 <= ($signed((wire1 ? {(~reg2513)} : (8'haa))) ?
                  $signed($signed(reg2468[(5'h11):(1'h0)])) : reg2574);
              reg2594 = {($unsigned(((reg31 > reg2588) ?
                      {reg2567} : (-reg2573))) <<< (~&(((8'hb6) ?
                      reg2565 : (8'hbd)) && (reg2497 ? (8'hbb) : reg2524)))),
                  (!(reg2466 ?
                      reg2586[(3'h4):(3'h4)] : {wire42[(2'h3):(2'h2)]}))};
              reg2595 <= (^{$unsigned(reg2588[(4'he):(3'h5)]),
                  ((wire1 ?
                      reg2589 : (reg2480 ?
                          (8'had) : reg2504)) <<< $unsigned({reg2529})),
                  (($unsigned(reg2584) << $unsigned((7'h4f))) ?
                      ((reg2524 || reg2548) != (reg34 > reg2591)) : reg2496)});
            end
        end
      for (forvar2596 = (1'h0); (forvar2596 < (3'h6)); forvar2596 = (forvar2596 + (1'h1)))
        begin
          reg2597 = {$signed(reg2524),
              {(((7'h4a) >= (+reg2468)) >> $signed((forvar2583 ?
                      wire3 : reg2528)))}};
          for (forvar2598 = (1'h0); (forvar2598 < (1'h1)); forvar2598 = (forvar2598 + (1'h1)))
            begin
              reg2599 = (8'ha6);
            end
          if ($unsigned($signed($unsigned(reg2570[(4'hb):(3'h5)]))))
            begin
              reg2600 <= ((($signed(reg2513[(5'h10):(3'h4)]) > ((reg2582 ?
                  reg2552 : reg2581) + ((7'h46) ~^ reg2572))) & wire42) * {$signed((7'h55)),
                  (reg2542 ^ reg2591)});
              reg2601 <= ($unsigned((8'hbf)) ?
                  $signed((($unsigned(reg2549) ? $unsigned(reg2461) : reg2498) ?
                      $unsigned($unsigned(reg2459)) : (|$signed(wire3)))) : {(|{reg2524}),
                      reg2581[(2'h2):(2'h2)],
                      ($signed(reg2574) < wire1[(2'h2):(1'h1)])});
              reg2602 <= (~|(forvar2554[(5'h15):(3'h6)] ?
                  reg29[(5'h14):(5'h13)] : ((reg2458[(5'h16):(3'h5)] ?
                      reg2560 : reg2601) + ($unsigned(forvar2583) <<< wire4))));
            end
          else
            begin
              reg2603 = (~&({((reg2542 & reg17) >= forvar2570[(3'h5):(3'h4)])} ?
                  $signed((^~(reg2573 & (8'ha6)))) : (+$signed({reg2573}))));
            end
          reg2604 <= reg18[(4'ha):(4'ha)];
        end
      reg2605 <= (|($signed((+$signed((7'h50)))) ~^ reg25[(5'h19):(4'he)]));
      if ((!$unsigned(reg2566)))
        begin
          if ((~reg2584[(1'h1):(1'h1)]))
            begin
              reg2606 <= ({$signed(forvar2566[(4'ha):(4'h9)])} << reg2498[(2'h3):(2'h3)]);
              reg2607 = ($unsigned($signed(reg2461[(2'h2):(1'h0)])) ?
                  reg2531[(3'h7):(3'h5)] : reg2576[(3'h5):(2'h2)]);
              reg2608 <= reg2599[(4'hd):(2'h3)];
            end
          else
            begin
              reg2607 = $unsigned(reg2557[(2'h3):(1'h1)]);
              reg2609 = reg2607[(1'h0):(1'h0)];
              reg2610 <= (((($signed(reg29) ? (^~reg2568) : reg2587) ?
                          {reg2587[(3'h5):(1'h0)],
                              (reg2472 >> (7'h47))} : $signed($signed(reg2600))) ?
                      (reg2521 >> $unsigned(forvar2570[(2'h2):(1'h1)])) : $unsigned($unsigned({forvar2554,
                          reg2491}))) ?
                  ((7'h51) ?
                      ($unsigned((~reg31)) + (!$unsigned(reg2551))) : reg2568[(2'h3):(2'h3)]) : $signed({((forvar2570 ?
                              (7'h44) : reg2570) ?
                          reg2496[(4'h8):(1'h0)] : (reg2568 ?
                              reg2474 : reg2585)),
                      reg34[(2'h3):(1'h1)],
                      (8'ha3)}));
              reg2611 = reg2512;
            end
        end
      else
        begin
          for (forvar2606 = (1'h0); (forvar2606 < (3'h6)); forvar2606 = (forvar2606 + (1'h1)))
            begin
              reg2607 = (|reg2552[(4'h8):(3'h4)]);
              reg2608 <= (reg2499 != (^reg30[(4'hd):(4'hd)]));
              reg2609 = {reg2570};
              reg2610 <= ($signed((reg2582 > $signed((^reg2573)))) ?
                  ($signed(((-reg2468) ~^ reg2498)) ?
                      $unsigned(($signed(reg2461) ?
                          $unsigned(reg2480) : reg2566)) : reg2478) : reg2575);
              reg2612 <= $unsigned({$signed({(+reg2588), (^reg2510)}),
                  (~|((wire3 >= reg2609) ?
                      reg2475[(1'h1):(1'h0)] : $unsigned(reg2504))),
                  reg31[(5'h13):(3'h7)]});
              reg2613 <= $unsigned((($signed($signed(reg2528)) ?
                      reg2472[(2'h3):(1'h1)] : reg2525) ?
                  $unsigned($signed(wire2453[(2'h3):(2'h3)])) : (~^((!wire2) & $signed(reg2604)))));
            end
          if ($unsigned($unsigned($unsigned({$unsigned((8'h9d)),
              reg2594[(2'h3):(1'h0)],
              reg2578[(1'h1):(1'h0)]}))))
            begin
              reg2614 <= ((|reg34) * ($signed((~(forvar2566 ?
                  reg2575 : forvar2606))) ^ (((reg2526 ?
                  reg2587 : wire1) + reg2515) >= {$signed((7'h58)),
                  forvar2583[(4'hf):(3'h5)]})));
            end
          else
            begin
              reg2615 = $unsigned(($signed(reg29[(4'hc):(4'hb)]) >> $signed(reg2546)));
            end
          for (forvar2616 = (1'h0); (forvar2616 < (3'h6)); forvar2616 = (forvar2616 + (1'h1)))
            begin
              reg2617 <= wire42;
              reg2618 = (!(^~$unsigned(reg2472)));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2619 = (1'h0); (forvar2619 < (3'h6)); forvar2619 = (forvar2619 + (1'h1)))
        begin
          if ((((8'ha5) > $unsigned(((reg2613 + reg2535) ?
              (reg2531 ?
                  (7'h56) : wire1) : reg2533[(1'h1):(1'h1)]))) ^ reg2588[(5'h1c):(5'h19)]))
            begin
              reg2620 = $unsigned(reg2463[(5'h18):(4'hb)]);
              reg2621 = (|((((|reg2576) * $unsigned(reg2612)) ?
                  reg2512[(1'h1):(1'h0)] : reg17) >> $unsigned((~^reg2569[(2'h2):(1'h1)]))));
            end
          else
            begin
              reg2622 <= $unsigned(reg2513[(2'h3):(2'h2)]);
              reg2623 = $unsigned(({(-$unsigned(reg34))} ?
                  {{(reg2496 ?
                              reg2582 : reg2551)}} : $signed(wire3[(3'h5):(2'h2)])));
            end
          if (reg2600[(4'h8):(4'h8)])
            begin
              reg2624 <= $signed($unsigned($unsigned($unsigned({reg2521,
                  reg2582,
                  reg2542}))));
              reg2625 = (($signed((7'h41)) ?
                      (~|((reg2472 << reg2608) >>> (~|reg2489))) : (7'h53)) ?
                  $unsigned(($signed((reg2549 * reg33)) & ((^(8'hb2)) ?
                      (~^reg30) : $unsigned(wire2453)))) : (^reg29));
              reg2626 <= $unsigned($signed(((reg2458 == reg2492[(3'h5):(3'h5)]) > reg2492[(1'h1):(1'h1)])));
            end
          else
            begin
              reg2625 = ((~|reg36[(3'h6):(1'h0)]) <= ({(|(7'h4f)),
                      (!(7'h49)),
                      {(!reg2525), reg2623, (~|reg2623)}} ?
                  reg2466[(5'h1a):(2'h3)] : (reg30[(1'h1):(1'h1)] > $signed($signed(reg2600)))));
              reg2627 = $unsigned(((^~$unsigned({(7'h47),
                  reg2605})) ^~ (((reg2572 <<< reg2525) ?
                      reg2510 : (reg2588 < reg2612)) ?
                  ({wire42, (7'h57), (8'h9f)} ?
                      $unsigned(reg2614) : (reg6 ?
                          reg2542 : reg2515)) : (~|(reg2567 > reg2524)))));
            end
        end
      reg2628 <= (reg2588 ?
          ({reg2613,
                  $unsigned((reg2491 ? reg2475 : reg2456)),
                  reg2564[(3'h7):(3'h6)]} ?
              reg2475[(1'h0):(1'h0)] : (((reg6 & reg2529) ^ reg2575) ?
                  (|(reg2515 ?
                      reg2458 : reg2606)) : reg2531)) : $signed(reg2513));
      for (forvar2629 = (1'h0); (forvar2629 < (1'h1)); forvar2629 = (forvar2629 + (1'h1)))
        begin
          reg2630 = $unsigned((-({(reg31 ? reg2542 : reg2613),
                  {reg2478, reg2628},
                  (reg2557 | (7'h4c))} ?
              (^$unsigned((8'ha6))) : (&$signed(reg2567)))));
          if ((^($unsigned($unsigned(reg2602)) <= (8'hbf))))
            begin
              reg2631 = reg33;
              reg2632 <= $signed(reg2486[(2'h2):(2'h2)]);
              reg2633 <= {reg2517};
            end
          else
            begin
              reg2632 <= ($unsigned(reg2631[(4'hf):(1'h1)]) ?
                  (~(~&$signed($signed(reg2544)))) : (($unsigned(((8'hb0) + reg2631)) ?
                      ((reg2588 >>> reg36) ?
                          (reg31 <= reg2632) : reg2568[(2'h3):(2'h2)]) : $signed($signed(reg2564))) == {reg2553[(3'h4):(3'h4)],
                      $unsigned($unsigned((8'ha5))),
                      $unsigned((reg2569 ? reg8 : (8'hab)))}));
            end
          reg2634 = (^~$signed($unsigned((|reg2632))));
        end
      for (forvar2635 = (1'h0); (forvar2635 < (2'h2)); forvar2635 = (forvar2635 + (1'h1)))
        begin
          if ({$signed((8'hb1)), $unsigned($unsigned({$unsigned(reg2604)}))})
            begin
              reg2636 <= ($unsigned($signed($unsigned(reg2524[(1'h0):(1'h0)]))) ?
                  ($unsigned(($unsigned(wire42) ?
                      reg2573[(5'h14):(5'h11)] : $signed(reg2593))) * $unsigned(($signed(wire2508) > {reg8}))) : reg2627);
              reg2637 = forvar2619[(4'hd):(2'h2)];
              reg2638 = $unsigned($unsigned(reg2533[(5'h10):(4'hb)]));
              reg2639 <= (~&((|$unsigned($signed(reg2610))) ?
                  reg2564 : reg2621));
              reg2640 = (~|reg2478[(4'h9):(4'h8)]);
            end
          else
            begin
              reg2636 <= reg2526[(4'hd):(3'h5)];
              reg2637 = reg2547[(4'h9):(1'h1)];
              reg2639 <= $signed(((reg2556 ^ reg22) ?
                  $signed(reg2612[(5'h16):(3'h7)]) : $unsigned($signed((~^reg34)))));
            end
          reg2641 = reg2582[(2'h2):(1'h1)];
          if (reg34)
            begin
              reg2642 = reg2555;
              reg2643 <= ($signed(((^reg2478) || (reg2578[(1'h1):(1'h0)] ?
                  (reg5 != reg2546) : (8'hbf)))) * (8'hb3));
              reg2644 = $signed((-wire0[(3'h5):(2'h2)]));
              reg2645 = reg2468[(3'h5):(3'h5)];
              reg2646 = forvar2629[(3'h5):(3'h4)];
              reg2647 = (~^$signed(reg2612));
            end
          else
            begin
              reg2643 <= wire2[(2'h3):(2'h2)];
              reg2648 <= $signed((({(reg2463 ? reg2492 : reg2627)} ?
                  {$unsigned(reg2646),
                      $unsigned(reg2566),
                      forvar2629} : $signed($unsigned(reg2515))) ^ {$signed($signed(reg2461)),
                  (~^((7'h47) ? (8'ha7) : reg36))}));
              reg2649 = reg2531;
              reg2650 <= $signed((reg2578 ?
                  reg2498[(4'h8):(2'h2)] : (~^$unsigned($signed(reg2645)))));
            end
        end
    end
  module179 #() modinst2652 (wire2651, clk, reg2632, reg30, reg2499, reg2557, reg2503, reg25);
  assign wire2653 = $unsigned(reg2624[(1'h1):(1'h0)]);
  module1961 #() modinst2655 (.wire1962(reg2487), .wire1964(reg6), .wire1965(reg2586), .y(wire2654), .wire1963(reg17), .clk(clk), .wire1966(reg2555));
  always
    @(posedge clk) begin
      if ($unsigned(reg2533))
        begin
          reg2656 = $unsigned(reg2534[(2'h2):(1'h1)]);
          for (forvar2657 = (1'h0); (forvar2657 < (2'h2)); forvar2657 = (forvar2657 + (1'h1)))
            begin
              reg2658 = (~|$signed((|($signed(reg2588) ?
                  reg2535 : reg2604[(2'h2):(1'h0)]))));
              reg2659 <= ((~&$unsigned($unsigned({reg2586,
                      reg2472,
                      reg2650}))) ?
                  (!$signed(($signed(reg2614) ?
                      (wire42 ?
                          (8'hb6) : reg2503) : reg2528[(4'ha):(1'h0)]))) : wire2654);
              reg2660 <= wire0[(3'h5):(1'h0)];
            end
          if ($unsigned($signed(reg2643)))
            begin
              reg2661 <= {(+$signed(reg2633[(4'hd):(4'ha)])), reg2588};
              reg2662 = $signed($signed(($unsigned(reg2529) ?
                  (+$signed(reg25)) : reg2512[(2'h3):(2'h3)])));
            end
          else
            begin
              reg2662 = {($signed($unsigned($signed(reg30))) ?
                      reg2643[(4'h8):(1'h1)] : $signed(reg2515[(4'hf):(4'hd)])),
                  $signed($signed({(reg27 <= reg2499)})),
                  $signed(wire2653)};
              reg2663 = (~&(+reg2499));
              reg2664 <= (7'h41);
            end
        end
      else
        begin
          reg2656 = (8'hb1);
          reg2657 = reg2608;
          for (forvar2658 = (1'h0); (forvar2658 < (2'h2)); forvar2658 = (forvar2658 + (1'h1)))
            begin
              reg2662 = (({$unsigned(reg2605[(5'h11):(4'ha)])} ?
                      reg2568 : {reg2491}) ?
                  reg2614 : (forvar2657 * {reg17[(5'h17):(5'h10)],
                      ($signed((7'h58)) ? reg2582 : (^~reg2517))}));
              reg2664 <= ($unsigned($signed($unsigned(reg2510))) & (+($signed($unsigned(reg2567)) ?
                  ((~^reg2466) == (wire1 <<< wire2453)) : {$unsigned(reg2468),
                      {(8'ha4)},
                      wire3[(3'h4):(2'h2)]})));
              reg2665 <= (reg2478 > reg2517);
            end
          reg2666 = $unsigned(reg2573);
          for (forvar2667 = (1'h0); (forvar2667 < (3'h4)); forvar2667 = (forvar2667 + (1'h1)))
            begin
              reg2668 = ({(~|(~^$signed(reg8))),
                      $unsigned($unsigned(reg2588)),
                      (reg18[(4'h9):(1'h1)] + (~$unsigned(reg2622)))} ?
                  $signed((reg2458[(4'hb):(4'ha)] ?
                      $signed((^(7'h4c))) : ($unsigned(reg2573) ~^ (reg2480 * reg2461)))) : (-reg2533));
              reg2669 <= ($signed((((reg2466 != wire3) || wire3[(4'h9):(3'h6)]) ?
                  (8'h9f) : (-(~|reg2564)))) && (reg2606[(2'h3):(2'h2)] >> $signed({(~^(7'h41)),
                  {reg2547}})));
              reg2670 = reg2573;
              reg2671 = reg2613[(4'he):(2'h2)];
              reg2672 = {(~$signed((-reg2492))),
                  $signed({$signed(reg2504), wire2653[(1'h0):(1'h0)]}),
                  {reg2503[(2'h2):(2'h2)],
                      ($signed($unsigned(reg2559)) * reg2656[(1'h0):(1'h0)]),
                      wire3[(5'h12):(4'hd)]}};
              reg2673 = reg2582;
              reg2674 <= reg2524;
            end
          reg2675 = (|((&reg31[(4'hd):(1'h1)]) - (~&reg2515[(5'h1c):(4'h9)])));
        end
      reg2676 <= ($signed((~&($unsigned(wire2653) == reg2675))) ^~ $signed(reg2458[(5'h1a):(4'hb)]));
      reg2677 <= ($signed(wire2651[(3'h5):(1'h0)]) ?
          ($signed((reg2582 <<< (+reg2639))) ?
              reg2595 : ((reg25 ?
                  reg2521 : (~^reg6)) ^ $signed(wire2651[(1'h1):(1'h0)]))) : (reg2503[(4'hf):(2'h2)] ?
              $unsigned($signed((reg2675 ? reg30 : reg2586))) : (~|reg2487)));
      if (({$unsigned({(!reg2564)})} ?
          ((!$unsigned($signed(reg2557))) == (~(reg2665[(3'h6):(1'h1)] ^~ (8'ha2)))) : (reg2600 ~^ (reg2458 ^ (~((8'ha0) >= reg2578))))))
        begin
          for (forvar2678 = (1'h0); (forvar2678 < (3'h6)); forvar2678 = (forvar2678 + (1'h1)))
            begin
              reg2679 = (8'hb1);
            end
          for (forvar2680 = (1'h0); (forvar2680 < (3'h4)); forvar2680 = (forvar2680 + (1'h1)))
            begin
              reg2681 = ($signed(((wire2653[(4'h8):(1'h1)] * (~^wire3)) + $signed((reg2547 + reg2529)))) ?
                  $signed(($signed(reg2535[(1'h1):(1'h0)]) ?
                      $unsigned(reg2496) : (&$unsigned(reg2549)))) : reg2456);
              reg2682 <= reg2660[(4'h8):(2'h2)];
              reg2683 <= ({reg2474, $signed({reg2593, $unsigned(reg2466)})} ?
                  reg2459 : ((reg2682 ?
                          {reg2675,
                              reg2551,
                              (-wire3)} : (reg2487[(1'h0):(1'h0)] & $unsigned(reg2472))) ?
                      wire0 : ((~&(-wire2653)) ?
                          (reg2517[(2'h3):(1'h0)] | wire2651) : ((7'h57) < (~reg2593)))));
              reg2684 = $unsigned($unsigned((^reg2503[(1'h1):(1'h1)])));
              reg2685 = reg2549;
            end
          reg2686 = reg2557;
          reg2687 <= $unsigned($unsigned($unsigned(((reg2661 >>> wire2651) ^~ {wire0,
              reg2524}))));
          reg2688 <= $unsigned(reg2552[(2'h2):(1'h0)]);
          if (({reg2497,
              $unsigned($unsigned(reg2648)),
              reg2604[(2'h3):(1'h1)]} != reg2602[(1'h1):(1'h1)]))
            begin
              reg2689 <= ((&reg2660[(3'h4):(1'h0)]) - ($signed($signed((reg2658 && (8'hab)))) ?
                  (-((reg2569 ?
                      (8'haa) : (7'h52)) > reg18[(5'h10):(4'ha)])) : (((reg2633 >= wire2453) <<< {reg2675,
                          (8'ha2),
                          reg2675}) ?
                      reg18[(5'h14):(4'hc)] : ((reg2564 ?
                          reg2491 : reg2662) <<< (forvar2680 >> reg2576)))));
            end
          else
            begin
              reg2690 = $signed($unsigned({((7'h56) ^~ (8'hba)),
                  $unsigned($unsigned(reg2593))}));
              reg2691 <= ($unsigned(reg2472) ?
                  $unsigned((reg2531[(5'h1a):(5'h19)] ?
                      reg2489[(3'h5):(2'h3)] : $unsigned((~&(7'h56))))) : (((|reg2478) ?
                      $signed(reg2535[(4'h9):(2'h3)]) : ({reg2628} ?
                          (reg2663 < reg2557) : reg2573[(4'he):(4'h9)])) && (reg2492 ?
                      (^~(reg2610 ? reg2546 : reg2544)) : (|$unsigned(reg8)))));
              reg2692 = {((reg2668 ?
                      reg2491 : reg2557[(3'h7):(3'h7)]) + (|reg2478))};
              reg2693 = $unsigned((~|(+(-((7'h4c) - wire2453)))));
            end
          reg2694 = (~^reg2498);
        end
      else
        begin
          reg2678 <= ((8'hbb) + (&reg2525));
          if ((reg2498 & reg2670))
            begin
              reg2679 = (({(7'h55),
                      ((8'hb6) << reg2566)} ^~ reg2540[(1'h0):(1'h0)]) ?
                  (7'h54) : wire3);
              reg2680 <= ((|(|(+$signed(reg2524)))) ?
                  ($signed(reg2475) <<< $signed(reg2692)) : {(($unsigned((8'hb0)) * $signed(reg2546)) + (reg2588 <= {reg2612,
                          reg17})),
                      (+{wire0[(2'h3):(1'h0)]})});
              reg2682 <= reg2546[(4'hc):(3'h7)];
              reg2684 = (~reg2458);
              reg2685 = $unsigned($unsigned($signed($unsigned((reg2679 ?
                  reg2458 : (7'h4b))))));
              reg2687 <= reg2672;
            end
          else
            begin
              reg2680 <= (8'ha0);
              reg2682 <= $unsigned($unsigned((reg2692 >= (~&$unsigned(reg2578)))));
            end
          reg2688 <= wire4[(5'h16):(5'h11)];
          for (forvar2689 = (1'h0); (forvar2689 < (2'h3)); forvar2689 = (forvar2689 + (1'h1)))
            begin
              reg2691 <= ((reg2694[(4'hb):(4'h9)] ?
                      wire0[(3'h4):(3'h4)] : reg6[(4'he):(2'h3)]) ?
                  $signed((reg2661 ?
                      reg2694[(4'hf):(3'h5)] : $signed((~^reg2686)))) : $signed($signed($unsigned(reg2549))));
              reg2695 <= ($signed($signed(reg2528[(4'he):(4'he)])) ?
                  (7'h40) : (~&(!reg2498[(4'h8):(3'h5)])));
              reg2696 <= (((|{reg2670}) ~^ (|(+(^reg2529)))) ?
                  $signed($signed($signed({reg2639}))) : $unsigned(($unsigned((-(8'hba))) ?
                      (reg30 ?
                          $signed(wire0) : $unsigned(reg2664)) : {reg2534})));
              reg2697 <= (reg2458[(3'h7):(1'h0)] ^ reg2617[(3'h6):(2'h2)]);
              reg2698 = ((~reg2547[(4'h8):(4'h8)]) >> reg18);
              reg2699 = reg2681;
            end
        end
      reg2700 <= ((~^(^reg2687[(4'hb):(1'h0)])) ?
          (({(|reg2683)} ?
              $signed($unsigned(wire2)) : $signed(reg2463[(3'h7):(3'h7)])) < (reg2474[(2'h2):(2'h2)] == (|$unsigned(reg2542)))) : $signed(reg18[(3'h7):(2'h3)]));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module43  (y, clk, wire48, wire47, wire46, wire45, wire44);
  output wire [(32'hbb8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h16):(1'h0)] wire48;
  input wire [(5'h13):(1'h0)] wire47;
  input wire signed [(5'h15):(1'h0)] wire46;
  input wire signed [(3'h5):(1'h0)] wire45;
  input wire signed [(2'h3):(1'h0)] wire44;
  wire signed [(5'h17):(1'h0)] wire2452;
  wire [(4'h9):(1'h0)] wire2451;
  wire signed [(4'he):(1'h0)] wire2450;
  wire [(2'h3):(1'h0)] wire2449;
  wire [(5'h17):(1'h0)] wire2448;
  wire [(4'hb):(1'h0)] wire2443;
  wire [(5'h1c):(1'h0)] wire1273;
  wire [(5'h18):(1'h0)] wire51;
  wire [(5'h13):(1'h0)] wire50;
  wire [(4'he):(1'h0)] wire49;
  wire [(5'h1f):(1'h0)] wire1392;
  wire signed [(5'h10):(1'h0)] wire1393;
  wire signed [(5'h15):(1'h0)] wire1430;
  wire signed [(4'hc):(1'h0)] wire1431;
  wire [(5'h1c):(1'h0)] wire1432;
  wire [(2'h2):(1'h0)] wire2441;
  reg [(3'h4):(1'h0)] reg2447 = (1'h0);
  reg [(4'hd):(1'h0)] reg1275 = (1'h0);
  reg [(5'h17):(1'h0)] reg1280 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1281 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1286 = (1'h0);
  reg [(5'h19):(1'h0)] reg1287 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1290 = (1'h0);
  reg [(3'h4):(1'h0)] reg1291 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1292 = (1'h0);
  reg [(5'h18):(1'h0)] reg1296 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1298 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1300 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1303 = (1'h0);
  reg [(4'ha):(1'h0)] reg1304 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1310 = (1'h0);
  reg [(4'ha):(1'h0)] reg1312 = (1'h0);
  reg [(5'h16):(1'h0)] reg1313 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1314 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1315 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1317 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1319 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1320 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1321 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1322 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1325 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1332 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1336 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1337 = (1'h0);
  reg [(5'h10):(1'h0)] reg1342 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1344 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1348 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1349 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1351 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1354 = (1'h0);
  reg [(5'h14):(1'h0)] reg1355 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1356 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1357 = (1'h0);
  reg [(4'hf):(1'h0)] reg1358 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1359 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1363 = (1'h0);
  reg [(5'h12):(1'h0)] reg1365 = (1'h0);
  reg [(5'h11):(1'h0)] reg1368 = (1'h0);
  reg [(3'h7):(1'h0)] reg1369 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1371 = (1'h0);
  reg [(4'ha):(1'h0)] reg1379 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1383 = (1'h0);
  reg [(4'hf):(1'h0)] reg1386 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1387 = (1'h0);
  reg [(5'h10):(1'h0)] reg1390 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1391 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1397 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1398 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1399 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1400 = (1'h0);
  reg [(2'h3):(1'h0)] reg1401 = (1'h0);
  reg [(3'h7):(1'h0)] reg1407 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1408 = (1'h0);
  reg [(2'h3):(1'h0)] reg1409 = (1'h0);
  reg [(5'h14):(1'h0)] reg1410 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1405 = (1'h0);
  reg [(5'h13):(1'h0)] reg1413 = (1'h0);
  reg [(3'h6):(1'h0)] reg1414 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1416 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1419 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1421 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1424 = (1'h0);
  reg [(3'h7):(1'h0)] reg1427 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1428 = (1'h0);
  reg [(3'h6):(1'h0)] reg1429 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2446 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2445 = (1'h0);
  reg [(5'h14):(1'h0)] reg2444 = (1'h0);
  reg [(2'h3):(1'h0)] reg1426 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1425 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1423 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1422 = (1'h0);
  reg [(4'hb):(1'h0)] reg1420 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1418 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1417 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1415 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1412 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1411 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1402 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1400 = (1'h0);
  reg [(4'hf):(1'h0)] reg1406 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1405 = (1'h0);
  reg [(5'h11):(1'h0)] reg1404 = (1'h0);
  reg [(5'h17):(1'h0)] reg1403 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1402 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1396 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1395 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1394 = (1'h0);
  reg [(4'hc):(1'h0)] reg1372 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1367 = (1'h0);
  reg [(3'h5):(1'h0)] reg1366 = (1'h0);
  reg [(4'ha):(1'h0)] reg1389 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1388 = (1'h0);
  reg [(5'h10):(1'h0)] reg1385 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1384 = (1'h0);
  reg [(3'h6):(1'h0)] reg1382 = (1'h0);
  reg [(5'h10):(1'h0)] reg1381 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1380 = (1'h0);
  reg [(4'he):(1'h0)] reg1378 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1377 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1376 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1375 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1374 = (1'h0);
  reg [(5'h11):(1'h0)] reg1373 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1372 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1370 = (1'h0);
  reg [(5'h18):(1'h0)] reg1367 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1366 = (1'h0);
  reg [(5'h10):(1'h0)] reg1364 = (1'h0);
  reg [(4'hb):(1'h0)] reg1362 = (1'h0);
  reg [(4'hb):(1'h0)] reg1361 = (1'h0);
  reg [(3'h5):(1'h0)] reg1360 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar1353 = (1'h0);
  reg [(4'ha):(1'h0)] reg1352 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1335 = (1'h0);
  reg [(4'hf):(1'h0)] reg1350 = (1'h0);
  reg [(5'h13):(1'h0)] reg1347 = (1'h0);
  reg [(4'hb):(1'h0)] reg1346 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1345 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1343 = (1'h0);
  reg [(4'h8):(1'h0)] reg1341 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1340 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1339 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1338 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1335 = (1'h0);
  reg [(4'h8):(1'h0)] reg1334 = (1'h0);
  reg [(4'ha):(1'h0)] reg1333 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1331 = (1'h0);
  reg [(5'h12):(1'h0)] reg1330 = (1'h0);
  reg [(5'h16):(1'h0)] reg1329 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1328 = (1'h0);
  reg [(5'h11):(1'h0)] reg1327 = (1'h0);
  reg [(5'h16):(1'h0)] reg1326 = (1'h0);
  reg [(4'hb):(1'h0)] reg1324 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1323 = (1'h0);
  reg [(4'h9):(1'h0)] reg1318 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1316 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1311 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1309 = (1'h0);
  reg [(5'h13):(1'h0)] reg1308 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1307 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1306 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1305 = (1'h0);
  reg [(3'h6):(1'h0)] reg1302 = (1'h0);
  reg [(2'h3):(1'h0)] reg1301 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1299 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1297 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1295 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1294 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1293 = (1'h0);
  reg [(3'h6):(1'h0)] reg1289 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1288 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1283 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1285 = (1'h0);
  reg [(5'h14):(1'h0)] reg1284 = (1'h0);
  reg [(5'h14):(1'h0)] reg1283 = (1'h0);
  reg [(4'h9):(1'h0)] reg1282 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1279 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1278 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1277 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1276 = (1'h0);
  assign y = {wire2452,
                 wire2451,
                 wire2450,
                 wire2449,
                 wire2448,
                 wire2443,
                 wire1273,
                 wire51,
                 wire50,
                 wire49,
                 wire1392,
                 wire1393,
                 wire1430,
                 wire1431,
                 wire1432,
                 wire2441,
                 reg2447,
                 reg1275,
                 reg1280,
                 reg1281,
                 reg1286,
                 reg1287,
                 reg1290,
                 reg1291,
                 reg1292,
                 reg1296,
                 reg1298,
                 reg1300,
                 reg1303,
                 reg1304,
                 reg1310,
                 reg1312,
                 reg1313,
                 reg1314,
                 reg1315,
                 reg1317,
                 reg1319,
                 reg1320,
                 reg1321,
                 reg1322,
                 reg1325,
                 reg1332,
                 reg1336,
                 reg1337,
                 reg1342,
                 reg1344,
                 reg1348,
                 reg1349,
                 reg1351,
                 reg1354,
                 reg1355,
                 reg1356,
                 reg1357,
                 reg1358,
                 reg1359,
                 reg1363,
                 reg1365,
                 reg1368,
                 reg1369,
                 reg1371,
                 reg1379,
                 reg1383,
                 reg1386,
                 reg1387,
                 reg1390,
                 reg1391,
                 reg1397,
                 reg1398,
                 reg1399,
                 reg1400,
                 reg1401,
                 reg1407,
                 reg1408,
                 reg1409,
                 reg1410,
                 reg1405,
                 reg1413,
                 reg1414,
                 reg1416,
                 reg1419,
                 reg1421,
                 reg1424,
                 reg1427,
                 reg1428,
                 reg1429,
                 reg2446,
                 reg2445,
                 reg2444,
                 reg1426,
                 reg1425,
                 reg1423,
                 reg1422,
                 reg1420,
                 reg1418,
                 reg1417,
                 forvar1415,
                 forvar1412,
                 reg1411,
                 reg1402,
                 forvar1400,
                 reg1406,
                 forvar1405,
                 reg1404,
                 reg1403,
                 forvar1402,
                 reg1396,
                 forvar1395,
                 forvar1394,
                 reg1372,
                 forvar1367,
                 reg1366,
                 reg1389,
                 forvar1388,
                 reg1385,
                 reg1384,
                 reg1382,
                 reg1381,
                 reg1380,
                 reg1378,
                 reg1377,
                 reg1376,
                 reg1375,
                 reg1374,
                 reg1373,
                 forvar1372,
                 reg1370,
                 reg1367,
                 forvar1366,
                 reg1364,
                 reg1362,
                 reg1361,
                 reg1360,
                 forvar1353,
                 reg1352,
                 forvar1335,
                 reg1350,
                 reg1347,
                 reg1346,
                 reg1345,
                 reg1343,
                 reg1341,
                 reg1340,
                 reg1339,
                 reg1338,
                 reg1335,
                 reg1334,
                 reg1333,
                 reg1331,
                 reg1330,
                 reg1329,
                 reg1328,
                 reg1327,
                 reg1326,
                 reg1324,
                 reg1323,
                 reg1318,
                 forvar1316,
                 forvar1311,
                 reg1309,
                 reg1308,
                 reg1307,
                 forvar1306,
                 forvar1305,
                 reg1302,
                 reg1301,
                 forvar1299,
                 reg1297,
                 reg1295,
                 reg1294,
                 reg1293,
                 reg1289,
                 reg1288,
                 forvar1283,
                 reg1285,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 (1'h0)};
  assign wire49 = (^~($unsigned({{wire47}}) & ($unsigned((wire46 ?
                      wire48 : wire44)) * wire47[(4'he):(4'he)])));
  assign wire50 = {wire46[(3'h6):(1'h1)], (7'h46)};
  assign wire51 = $signed(wire50);
  module52 #() modinst1274 (wire1273, clk, wire46, wire49, wire51, wire47, wire48);
  always
    @(posedge clk) begin
      reg1275 <= (~&$unsigned((((wire47 >= wire47) > $unsigned(wire51)) ?
          (-(wire49 ? wire44 : wire51)) : $signed((wire48 ?
              wire1273 : wire44)))));
      if (($unsigned(((wire45 > wire49) + $signed((!(8'hae))))) ?
          wire46[(4'hc):(4'ha)] : wire46[(2'h3):(1'h1)]))
        begin
          reg1276 = wire44[(1'h1):(1'h0)];
          reg1277 = reg1275;
          if ((wire49 < (($unsigned(wire48[(3'h4):(3'h4)]) >>> ($unsigned(wire49) * $unsigned(wire1273))) ?
              $signed((~|(8'had))) : {wire47,
                  $signed((wire51 >= wire50)),
                  (^~wire48)})))
            begin
              reg1278 = $unsigned($unsigned({$unsigned((~reg1276))}));
              reg1279 = (wire51 ?
                  (^$signed(((reg1275 ?
                      wire48 : wire44) < reg1276[(3'h5):(3'h4)]))) : {$signed($unsigned($signed(wire50)))});
            end
          else
            begin
              reg1278 = ((+wire51) ?
                  ($signed((^~wire44[(1'h1):(1'h0)])) ?
                      wire45[(1'h1):(1'h1)] : (reg1279 != reg1275)) : $signed(reg1279[(2'h3):(1'h0)]));
              reg1280 <= wire1273[(5'h1b):(4'h9)];
              reg1281 <= $unsigned($signed($signed(({(8'ha0)} ?
                  reg1275[(4'hb):(2'h2)] : $unsigned(reg1278)))));
              reg1282 = $signed(((7'h52) || ((+wire44) << $signed($unsigned(wire1273)))));
              reg1283 = $signed($unsigned($signed((+$signed(wire48)))));
              reg1284 = (wire45[(1'h1):(1'h0)] ?
                  wire50[(2'h3):(2'h2)] : reg1280);
            end
          reg1285 = {(~^(((reg1281 ?
                  (8'hb5) : wire1273) == (wire49 < reg1275)) * {(reg1276 ^ wire50),
                  wire50,
                  $signed(reg1281)}))};
        end
      else
        begin
          reg1280 <= reg1283;
          reg1282 = $signed($unsigned(wire49[(3'h4):(2'h2)]));
          for (forvar1283 = (1'h0); (forvar1283 < (3'h6)); forvar1283 = (forvar1283 + (1'h1)))
            begin
              reg1284 = $signed(reg1276[(4'he):(4'h8)]);
              reg1286 <= forvar1283[(3'h4):(3'h4)];
              reg1287 <= wire44;
            end
          if (forvar1283[(4'hc):(2'h3)])
            begin
              reg1288 = $unsigned(($unsigned(reg1287[(5'h13):(4'h8)]) ?
                  $unsigned({(reg1282 ? reg1284 : (8'h9d)),
                      $unsigned(wire45),
                      $signed(wire51)}) : $signed(((&wire50) <= reg1275[(1'h0):(1'h0)]))));
              reg1289 = $unsigned(wire50);
              reg1290 <= (forvar1283[(4'hf):(2'h2)] ?
                  (~|($signed(forvar1283[(5'h11):(4'hd)]) ?
                      $unsigned((wire51 << reg1289)) : $signed($unsigned(wire44)))) : $unsigned((reg1277 ?
                      ($signed(reg1278) ?
                          $signed(wire44) : reg1280[(5'h10):(3'h5)]) : ($unsigned(reg1280) - reg1285))));
              reg1291 <= (^~$unsigned(reg1285));
              reg1292 <= reg1291[(1'h0):(1'h0)];
            end
          else
            begin
              reg1290 <= reg1288;
              reg1293 = $unsigned($unsigned(($signed((wire48 > wire49)) ?
                  reg1280[(5'h10):(2'h3)] : reg1290[(5'h18):(4'he)])));
              reg1294 = reg1282;
              reg1295 = (($unsigned($unsigned($signed((8'hbe)))) <<< wire50) < {$signed((reg1281[(4'hd):(1'h0)] & (~(8'ha5)))),
                  ((reg1287 ~^ (wire50 ? reg1275 : wire45)) ?
                      $unsigned(reg1280[(2'h3):(1'h1)]) : ({reg1276,
                          wire46} ^ wire48[(4'hd):(3'h4)])),
                  $signed($signed(reg1284))});
              reg1296 <= $unsigned($unsigned($signed($unsigned((|reg1284)))));
              reg1297 = ((!forvar1283[(3'h6):(2'h2)]) ?
                  forvar1283[(4'hc):(3'h7)] : (({$signed(reg1278),
                              reg1285,
                              $unsigned(reg1289)} ?
                          (reg1275 ?
                              wire49[(3'h5):(2'h3)] : (reg1279 <<< reg1282)) : {reg1284[(4'hb):(1'h0)],
                              {reg1280}}) ?
                      reg1277[(5'h13):(5'h12)] : ((reg1289 & (reg1293 ?
                              reg1285 : reg1285)) ?
                          $signed((+wire47)) : {(wire50 + forvar1283)})));
            end
          reg1298 <= $signed($signed($signed($unsigned(reg1281[(4'he):(4'hd)]))));
          for (forvar1299 = (1'h0); (forvar1299 < (3'h5)); forvar1299 = (forvar1299 + (1'h1)))
            begin
              reg1300 <= $signed($signed((-{reg1297,
                  $unsigned(reg1298),
                  (reg1291 ^ (8'h9f))})));
              reg1301 = forvar1283[(5'h11):(5'h10)];
              reg1302 = ($signed(((+{reg1295}) >>> reg1275[(2'h2):(2'h2)])) ?
                  $unsigned((((reg1301 <= wire44) ?
                          (reg1280 >>> forvar1299) : $signed(reg1301)) ?
                      $signed({forvar1283}) : $unsigned($unsigned(wire48)))) : ($signed(reg1297[(4'ha):(4'h9)]) ?
                      (~{(8'had),
                          reg1288,
                          (reg1279 ?
                              reg1285 : reg1282)}) : $unsigned((!$signed(reg1300)))));
              reg1303 <= {wire47[(4'hb):(4'h8)],
                  (~^($signed(wire50[(2'h3):(2'h2)]) >> ($unsigned(reg1289) ?
                      reg1294[(2'h3):(2'h2)] : $signed(wire46))))};
              reg1304 <= reg1295[(4'hc):(1'h0)];
            end
        end
      for (forvar1305 = (1'h0); (forvar1305 < (3'h6)); forvar1305 = (forvar1305 + (1'h1)))
        begin
          for (forvar1306 = (1'h0); (forvar1306 < (2'h2)); forvar1306 = (forvar1306 + (1'h1)))
            begin
              reg1307 = $unsigned({(8'ha9)});
            end
        end
      reg1308 = $unsigned((reg1285 ?
          $signed(($signed(reg1287) <= (reg1276 + reg1278))) : $signed((wire47 ?
              reg1302 : $unsigned(forvar1306)))));
    end
  always
    @(posedge clk) begin
      reg1309 = (~^$unsigned((~&(-(^wire1273)))));
      reg1310 <= ($unsigned(wire1273) ~^ $unsigned(wire50[(3'h6):(3'h6)]));
      for (forvar1311 = (1'h0); (forvar1311 < (2'h3)); forvar1311 = (forvar1311 + (1'h1)))
        begin
          reg1312 <= {$signed((|($unsigned(wire1273) << (wire44 ^~ reg1309))))};
          reg1313 <= reg1296[(4'hf):(4'he)];
          reg1314 <= {reg1304,
              $signed((((reg1296 ?
                  (7'h57) : reg1300) ^~ reg1300[(5'h15):(1'h0)]) > reg1313[(3'h7):(1'h1)]))};
          reg1315 <= (reg1290 & $unsigned({wire51[(3'h4):(1'h1)]}));
        end
      for (forvar1316 = (1'h0); (forvar1316 < (2'h2)); forvar1316 = (forvar1316 + (1'h1)))
        begin
          reg1317 <= (^($signed((!(^~wire47))) >>> reg1280));
          if ({$unsigned(($unsigned(reg1281) ?
                  (7'h4c) : {$signed(reg1275), (~reg1287)})),
              (&reg1303)})
            begin
              reg1318 = $signed(wire1273);
              reg1319 <= $signed({$unsigned($signed((&reg1314)))});
              reg1320 <= wire46;
              reg1321 <= $signed({(((^~reg1313) << $signed(wire45)) ?
                      wire46[(4'hb):(4'h9)] : (~|(reg1291 ?
                          reg1280 : reg1320)))});
              reg1322 <= {($unsigned(($signed(wire47) ?
                          reg1315[(2'h2):(2'h2)] : (wire1273 ?
                              reg1298 : reg1314))) ?
                      (((reg1313 - reg1310) >= reg1281[(3'h5):(2'h3)]) ?
                          (reg1319 * (7'h58)) : {$signed(wire47),
                              (wire45 || wire46)}) : $unsigned(((reg1309 ?
                          (7'h51) : wire49) + (wire1273 ? reg1321 : reg1321)))),
                  wire50[(3'h7):(3'h4)]};
              reg1323 = (!$unsigned(forvar1316[(2'h3):(2'h3)]));
            end
          else
            begin
              reg1319 <= (|$signed((reg1292 + reg1318)));
              reg1320 <= (($unsigned((~^((8'hb8) ? wire47 : reg1315))) ?
                  (reg1317[(1'h0):(1'h0)] != ((~wire47) ?
                      (reg1323 ?
                          reg1312 : reg1286) : wire46)) : (($signed(reg1281) ?
                      (|reg1292) : (reg1286 ~^ reg1291)) ^~ ({forvar1311,
                      reg1281} * (7'h43)))) | reg1318[(1'h0):(1'h0)]);
              reg1323 = {reg1319[(3'h5):(2'h3)],
                  $signed($signed($unsigned((reg1312 ? wire48 : wire1273)))),
                  wire46[(4'he):(4'h8)]};
              reg1324 = reg1318[(1'h0):(1'h0)];
              reg1325 <= (!(($signed($unsigned(reg1314)) ?
                      reg1296 : wire44[(2'h3):(1'h1)]) ?
                  $unsigned($signed({wire44})) : (8'h9c)));
              reg1326 = $unsigned($unsigned($signed(($signed(reg1314) ?
                  reg1315 : (reg1275 ~^ forvar1311)))));
            end
          if (forvar1316[(4'hf):(2'h2)])
            begin
              reg1327 = {$unsigned($unsigned((((8'hb0) >> reg1317) ?
                      reg1280 : (wire48 & reg1309)))),
                  {$unsigned(wire51[(5'h18):(4'hb)]),
                      $unsigned(($unsigned(reg1310) ?
                          (~|reg1291) : $signed(reg1315))),
                      wire49[(3'h7):(2'h2)]}};
              reg1328 = (~^($unsigned(($unsigned(reg1324) - wire47[(5'h11):(5'h10)])) ?
                  reg1281[(4'hd):(1'h1)] : reg1317[(1'h1):(1'h1)]));
              reg1329 = {$unsigned((~^forvar1311))};
              reg1330 = $unsigned(reg1290);
              reg1331 = reg1323;
              reg1332 <= (~^{reg1327, reg1323[(1'h0):(1'h0)]});
            end
          else
            begin
              reg1332 <= $signed({$unsigned($unsigned($unsigned(reg1325))),
                  reg1310});
              reg1333 = (+(($unsigned((reg1280 ^~ reg1314)) == ($unsigned(reg1300) ?
                      (reg1281 ? (8'h9c) : reg1325) : reg1313)) ?
                  (($signed(reg1314) ?
                          $signed(wire46) : reg1322[(1'h0):(1'h0)]) ?
                      ($unsigned(reg1304) ?
                          $unsigned(reg1275) : (wire45 << reg1286)) : ((reg1328 <= wire48) || $unsigned(wire50))) : (+(^~(reg1310 << reg1329)))));
              reg1334 = reg1329[(4'hc):(4'h9)];
            end
        end
      if ((reg1292 ~^ wire1273))
        begin
          if ((($signed((reg1324 ?
              ((8'ha5) ?
                  reg1328 : reg1291) : (~reg1329))) > $unsigned($signed($signed(reg1333)))) - (~&($signed({reg1334}) && $unsigned($unsigned(wire46))))))
            begin
              reg1335 = ((~(($unsigned(reg1328) ? (^~wire50) : reg1287) ?
                      $signed({reg1304,
                          reg1312,
                          (8'ha6)}) : $signed((8'haf)))) ?
                  ((&(!(forvar1316 <<< reg1300))) ?
                      (reg1300 | reg1318[(1'h1):(1'h1)]) : (~|{$unsigned(wire46)})) : (-wire45[(3'h4):(1'h1)]));
              reg1336 <= $signed(((reg1333 ^~ (7'h42)) ?
                  wire45[(1'h1):(1'h1)] : ({(reg1329 ? (8'hbd) : reg1290),
                          $unsigned(reg1317),
                          $unsigned(reg1286)} ?
                      forvar1316[(3'h7):(2'h3)] : ($unsigned(reg1298) == $signed(reg1327)))));
            end
          else
            begin
              reg1336 <= reg1329[(5'h12):(4'h8)];
              reg1337 <= $signed((!(~$signed(reg1286[(4'hc):(1'h0)]))));
              reg1338 = $unsigned(((~&($signed(reg1318) ?
                      (&reg1280) : (reg1319 << reg1310))) ?
                  $unsigned(reg1328) : {wire45[(3'h5):(2'h3)],
                      $signed($unsigned((7'h50)))}));
              reg1339 = ({(7'h47),
                  reg1333[(3'h6):(3'h4)]} <= reg1325[(5'h14):(3'h7)]);
              reg1340 = $signed(reg1310);
              reg1341 = $signed($unsigned(($signed((reg1328 ?
                      forvar1316 : (7'h49))) ?
                  (reg1325[(5'h15):(5'h11)] ?
                      wire44 : reg1333[(1'h0):(1'h0)]) : reg1312)));
              reg1342 <= (^~reg1281);
            end
          reg1343 = (^(reg1313 ?
              wire46[(1'h1):(1'h0)] : (^($signed((8'h9d)) || (reg1335 ?
                  reg1320 : forvar1316)))));
          if ((&($signed(wire49) <= reg1324)))
            begin
              reg1344 <= reg1318[(1'h0):(1'h0)];
              reg1345 = reg1312;
              reg1346 = ($signed((~&$signed(wire44[(1'h0):(1'h0)]))) ?
                  {reg1342[(3'h4):(3'h4)]} : reg1324[(2'h2):(1'h1)]);
              reg1347 = {$signed({wire44})};
            end
          else
            begin
              reg1344 <= $signed(reg1291);
              reg1348 <= ((~^(reg1337 ?
                  $unsigned($unsigned((8'ha6))) : $signed((~|reg1303)))) + $signed((8'hba)));
              reg1349 <= ((~&(~(&reg1333[(3'h6):(1'h1)]))) << {reg1347});
              reg1350 = reg1325[(3'h5):(3'h4)];
            end
        end
      else
        begin
          for (forvar1335 = (1'h0); (forvar1335 < (3'h4)); forvar1335 = (forvar1335 + (1'h1)))
            begin
              reg1338 = (($signed(wire44) ?
                  $signed((reg1345 & $signed(forvar1311))) : ((^~wire49) > reg1344[(5'h10):(4'hb)])) ^ ($signed(($signed(reg1327) ?
                  (|reg1291) : (wire50 ?
                      reg1338 : reg1348))) && ((|(^(8'hbc))) ?
                  reg1332 : {$signed(reg1329)})));
              reg1342 <= (8'hab);
              reg1343 = (+reg1312[(2'h2):(1'h0)]);
              reg1345 = reg1281[(3'h4):(1'h0)];
            end
          reg1348 <= (((+(7'h50)) ?
              (reg1339 >>> {(reg1343 | (7'h4c)),
                  (~&(8'hb2)),
                  (reg1332 ? wire46 : (8'haf))}) : $signed(reg1334)) * reg1281);
          reg1349 <= (forvar1335 ^ (~|$unsigned({(reg1334 << reg1331),
              (-reg1347),
              (wire1273 ? reg1322 : (8'haf))})));
          reg1351 <= (~&(wire49[(3'h6):(3'h4)] & reg1322[(2'h3):(2'h3)]));
          reg1352 = reg1331[(3'h7):(3'h6)];
        end
      for (forvar1353 = (1'h0); (forvar1353 < (3'h4)); forvar1353 = (forvar1353 + (1'h1)))
        begin
          if ({((((~&reg1340) ? $signed(forvar1335) : (~&reg1318)) ?
                      $signed((reg1337 <<< reg1340)) : ({(8'h9e),
                          (7'h51),
                          reg1320} != (8'hb2))) ?
                  ((~|$unsigned(reg1286)) ?
                      reg1352 : reg1324) : $signed((&(wire48 && reg1332)))),
              $signed((reg1300 && (-$unsigned((8'had)))))})
            begin
              reg1354 <= $signed(reg1331);
              reg1355 <= (reg1342[(5'h10):(4'hc)] ?
                  reg1321[(2'h2):(2'h2)] : $signed((~|reg1340[(3'h6):(1'h0)])));
              reg1356 <= (({(~|(^~reg1275))} ^~ wire45) ?
                  reg1318 : reg1342[(2'h2):(2'h2)]);
              reg1357 <= reg1329;
              reg1358 <= $unsigned(($signed(reg1319[(1'h1):(1'h1)]) ?
                  ((~^reg1325[(5'h1e):(5'h19)]) ^~ (~(reg1334 || (7'h46)))) : (reg1340[(4'hb):(1'h0)] ?
                      $signed(reg1339[(5'h10):(4'ha)]) : reg1345)));
              reg1359 <= forvar1353[(5'h17):(4'hd)];
              reg1360 = {(reg1330 ?
                      reg1275 : $signed(({(8'h9e), reg1352} <<< (reg1324 ?
                          reg1303 : reg1344))))};
            end
          else
            begin
              reg1360 = $unsigned(reg1348[(2'h3):(2'h3)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg1361 = {((reg1317 ?
              $signed(reg1357) : $unsigned(((8'ha0) || reg1275))) <= reg1303[(2'h3):(1'h0)]),
          {$unsigned(reg1280)},
          (~(~^((!reg1304) ?
              $signed(wire46) : ((7'h55) ? reg1296 : (8'h9e)))))};
      if (reg1292[(5'h10):(2'h3)])
        begin
          reg1362 = $signed(((reg1313 ?
                  ($signed(wire50) ?
                      (~^reg1344) : $signed(reg1361)) : ((reg1313 < reg1332) ?
                      reg1332[(5'h16):(2'h2)] : {reg1313, wire1273, reg1342})) ?
              $signed((8'haa)) : $signed(reg1298)));
        end
      else
        begin
          reg1363 <= (+reg1310[(3'h7):(3'h5)]);
        end
      reg1364 = $unsigned(reg1310[(3'h4):(2'h3)]);
      if (reg1313[(4'hd):(4'ha)])
        begin
          reg1365 <= $unsigned($signed(reg1320));
          for (forvar1366 = (1'h0); (forvar1366 < (3'h5)); forvar1366 = (forvar1366 + (1'h1)))
            begin
              reg1367 = reg1321;
              reg1368 <= $signed(reg1362);
              reg1369 <= reg1317;
              reg1370 = ((8'ha4) * ({((!(8'ha5)) ?
                      reg1342[(3'h5):(3'h4)] : reg1342[(4'hf):(3'h6)])} & reg1292));
              reg1371 <= $unsigned((($unsigned(reg1356) ?
                  (&$signed(wire50)) : (reg1300[(5'h19):(5'h12)] ^ reg1300)) | (8'hb1)));
            end
          for (forvar1372 = (1'h0); (forvar1372 < (3'h5)); forvar1372 = (forvar1372 + (1'h1)))
            begin
              reg1373 = reg1357[(4'hc):(1'h1)];
              reg1374 = (|(|reg1349[(5'h14):(1'h1)]));
              reg1375 = (&reg1348[(4'h8):(2'h3)]);
              reg1376 = reg1321[(3'h4):(1'h0)];
            end
          if (($unsigned($signed((~&wire51[(4'he):(4'hd)]))) ?
              ((~|{reg1363}) == {(reg1304[(3'h5):(1'h0)] ?
                      $unsigned(reg1280) : wire45[(2'h2):(2'h2)])}) : (^{(^~(reg1296 ?
                      (7'h47) : reg1348)),
                  reg1281[(5'h11):(3'h7)]})))
            begin
              reg1377 = $unsigned($unsigned((wire49[(4'h8):(3'h5)] ?
                  reg1319[(2'h3):(2'h2)] : {(wire1273 ~^ reg1317),
                      reg1290[(2'h3):(1'h1)],
                      $signed(reg1300)})));
              reg1378 = reg1342;
              reg1379 <= $signed($signed(wire44));
              reg1380 = (reg1319[(3'h6):(3'h4)] ?
                  {(reg1317[(1'h1):(1'h0)] ?
                          ((reg1304 ~^ reg1368) ?
                              reg1312[(1'h1):(1'h1)] : (reg1310 ?
                                  reg1322 : reg1362)) : {reg1367,
                              {reg1376},
                              $signed(reg1332)}),
                      reg1312[(3'h6):(1'h1)],
                      (8'hbf)} : reg1292);
              reg1381 = $signed(($unsigned(((^~reg1380) ?
                      reg1296 : reg1363[(1'h0):(1'h0)])) ?
                  $unsigned({reg1370,
                      (reg1371 ^ forvar1366),
                      (~^(7'h49))}) : $signed(((-reg1370) + $unsigned((7'h4c))))));
              reg1382 = (reg1291 ? $signed((+{$unsigned(reg1336)})) : reg1304);
            end
          else
            begin
              reg1379 <= $unsigned($unsigned((((^reg1292) ?
                      reg1379[(3'h6):(3'h6)] : (|reg1275)) ?
                  (-{reg1365, reg1344, (8'hb1)}) : (-$unsigned(forvar1372)))));
              reg1380 = (+((&(8'hb4)) ?
                  (+reg1363[(3'h7):(3'h7)]) : $signed(((reg1358 ?
                          reg1355 : reg1362) ?
                      ((8'ha0) ? reg1310 : reg1375) : (reg1314 ~^ reg1290)))));
              reg1383 <= reg1281;
              reg1384 = $unsigned($unsigned(wire50));
              reg1385 = reg1286;
              reg1386 <= $unsigned(((^$unsigned($signed(reg1280))) & ((7'h47) >= ((wire48 | reg1356) ?
                  $unsigned(reg1383) : $unsigned(reg1374)))));
              reg1387 <= (((|(|(~&(7'h46)))) ^ (reg1319 <= reg1312[(2'h2):(1'h1)])) & $signed($unsigned($unsigned((reg1356 ?
                  reg1376 : reg1380)))));
            end
          for (forvar1388 = (1'h0); (forvar1388 < (2'h3)); forvar1388 = (forvar1388 + (1'h1)))
            begin
              reg1389 = $unsigned(reg1380[(1'h0):(1'h0)]);
              reg1390 <= {$unsigned((reg1313[(5'h13):(2'h2)] * $signed(reg1368)))};
              reg1391 <= reg1344;
            end
        end
      else
        begin
          reg1366 = ($unsigned((|$signed($signed((8'hae))))) ?
              $signed($unsigned($unsigned({wire46,
                  (8'hbe),
                  reg1275}))) : {$signed($unsigned(wire48)),
                  {reg1382[(1'h0):(1'h0)]}});
          for (forvar1367 = (1'h0); (forvar1367 < (3'h6)); forvar1367 = (forvar1367 + (1'h1)))
            begin
              reg1370 = $signed($signed((reg1336[(1'h1):(1'h0)] ?
                  $unsigned(reg1336) : (reg1325[(2'h2):(1'h0)] ?
                      (forvar1367 ? reg1351 : (7'h51)) : (8'hb3)))));
              reg1372 = reg1300[(5'h13):(5'h10)];
              reg1373 = (~^$unsigned((|reg1290)));
              reg1374 = {{$unsigned($signed({reg1298, wire51, reg1391})),
                      {$unsigned(reg1370)},
                      $signed(({reg1355, (8'ha9)} << $unsigned(reg1303)))},
                  (7'h47)};
              reg1375 = reg1348;
            end
          reg1376 = $signed(reg1356[(4'h9):(2'h2)]);
          reg1377 = $signed((^~$signed(reg1381[(4'h8):(1'h0)])));
        end
    end
  assign wire1392 = reg1320;
  assign wire1393 = {(&$unsigned((~&$signed(reg1310))))};
  always
    @(posedge clk) begin
      for (forvar1394 = (1'h0); (forvar1394 < (3'h4)); forvar1394 = (forvar1394 + (1'h1)))
        begin
          for (forvar1395 = (1'h0); (forvar1395 < (3'h5)); forvar1395 = (forvar1395 + (1'h1)))
            begin
              reg1396 = (reg1369[(1'h0):(1'h0)] * $signed((~^((reg1281 ^ reg1386) || ((7'h4e) >>> reg1321)))));
              reg1397 <= {(|reg1300[(3'h5):(1'h1)]),
                  ((wire48[(4'hc):(4'ha)] >>> (+reg1312)) ?
                      $unsigned(((wire45 ? reg1358 : reg1310) ?
                          {reg1313} : $signed(reg1317))) : reg1379[(4'h9):(4'h8)]),
                  ($unsigned(($unsigned(reg1359) ? reg1310 : (+reg1280))) ?
                      reg1391 : (&(^~$signed(reg1348))))};
            end
        end
      reg1398 <= $unsigned(($unsigned($unsigned({reg1358})) != wire1273[(4'ha):(3'h4)]));
      reg1399 <= ((({{reg1280, wire45, wire47}, $signed(reg1291)} ?
          reg1396 : $unsigned(reg1351[(3'h5):(1'h1)])) >> {reg1314[(4'h8):(2'h2)]}) - reg1332);
      if (reg1344[(4'ha):(3'h5)])
        begin
          reg1400 <= reg1281;
          reg1401 <= (8'haa);
          for (forvar1402 = (1'h0); (forvar1402 < (3'h6)); forvar1402 = (forvar1402 + (1'h1)))
            begin
              reg1403 = (~(((8'hb3) ?
                      (wire46 ^~ $unsigned(reg1296)) : (+reg1349)) ?
                  {(8'hb5),
                      $signed($signed(reg1383))} : ($signed((reg1332 & wire1393)) != reg1314)));
              reg1404 = $signed(reg1387);
            end
          for (forvar1405 = (1'h0); (forvar1405 < (3'h5)); forvar1405 = (forvar1405 + (1'h1)))
            begin
              reg1406 = (reg1292[(5'h13):(4'hc)] ?
                  (($unsigned((reg1399 || wire47)) | ($signed(wire47) ?
                      {(7'h53)} : {reg1397})) | ({reg1355[(4'ha):(2'h2)]} ?
                      $signed((reg1315 >= (7'h55))) : ($signed(wire51) ?
                          (reg1296 ? reg1356 : reg1287) : (reg1321 ?
                              reg1342 : reg1371)))) : (reg1401 ?
                      (~|((^~wire46) ?
                          $signed(wire51) : (&reg1325))) : ((7'h49) ^~ $unsigned((^reg1348)))));
              reg1407 <= forvar1394;
              reg1408 <= $signed(reg1359);
            end
          reg1409 <= $signed($signed(((reg1406 ?
                  $signed(reg1325) : ((7'h53) && reg1320)) ?
              reg1396[(2'h2):(1'h0)] : (reg1275[(1'h1):(1'h0)] ?
                  reg1310 : (+wire1393)))));
          reg1410 <= ((&(reg1287[(1'h1):(1'h1)] ?
              (~^(!reg1296)) : reg1280)) < reg1280);
        end
      else
        begin
          for (forvar1400 = (1'h0); (forvar1400 < (2'h3)); forvar1400 = (forvar1400 + (1'h1)))
            begin
              reg1402 = reg1404;
              reg1405 <= wire51[(5'h12):(5'h12)];
              reg1406 = reg1371[(3'h6):(3'h5)];
            end
          reg1411 = (($signed({$unsigned(reg1320)}) ?
                  (~^reg1286) : ($unsigned((reg1342 == reg1397)) ?
                      reg1287 : forvar1405[(2'h3):(2'h2)])) ?
              (reg1409[(2'h2):(2'h2)] ?
                  (((reg1400 ?
                      reg1336 : reg1342) > ((7'h52) ~^ wire1273)) << reg1319) : reg1379) : {($signed($unsigned(reg1342)) | $signed({wire45,
                      reg1280}))});
        end
      for (forvar1412 = (1'h0); (forvar1412 < (3'h5)); forvar1412 = (forvar1412 + (1'h1)))
        begin
          reg1413 <= $unsigned({($unsigned(reg1281) ?
                  ((+wire49) <<< $signed(reg1396)) : {(reg1320 ?
                          reg1349 : reg1321)})});
          reg1414 <= reg1351;
          for (forvar1415 = (1'h0); (forvar1415 < (1'h0)); forvar1415 = (forvar1415 + (1'h1)))
            begin
              reg1416 <= $signed($unsigned((&wire46)));
            end
          reg1417 = reg1410[(4'he):(2'h3)];
          reg1418 = reg1332;
          reg1419 <= (7'h4b);
        end
      reg1420 = (~&($signed(reg1396[(1'h0):(1'h0)]) ?
          {(-(reg1387 | forvar1395)), reg1399[(4'h8):(2'h3)]} : (^reg1405)));
      if ((8'hb1))
        begin
          reg1421 <= $unsigned($signed($unsigned($unsigned($unsigned(wire48)))));
          reg1422 = (!($signed($signed((reg1402 || (8'hb6)))) ?
              {($unsigned(reg1407) ? (^~wire1393) : reg1387),
                  (+$unsigned(reg1349))} : (forvar1415[(1'h0):(1'h0)] ~^ $signed((reg1292 == reg1321)))));
          reg1423 = $signed(wire1273[(5'h1a):(4'h9)]);
        end
      else
        begin
          if ({{(($signed(reg1368) ? reg1303 : (7'h4e)) ?
                      ((reg1296 ~^ reg1404) ?
                          (~&reg1281) : (8'hb9)) : $unsigned({reg1298,
                          (8'hab)})),
                  reg1422},
              (((^~{wire51, reg1401}) ?
                  ($unsigned(reg1398) ?
                      (~&forvar1395) : wire48[(5'h14):(3'h7)]) : $unsigned($unsigned(reg1371))) << $unsigned(($signed((7'h54)) ?
                  reg1402[(3'h6):(2'h3)] : wire1393[(3'h6):(2'h3)])))})
            begin
              reg1422 = (&{((~wire46[(4'hc):(2'h2)]) >= (^~$unsigned(reg1416))),
                  (|(~^((8'hbe) >>> reg1291))),
                  $unsigned($signed($unsigned(reg1398)))});
              reg1424 <= $signed((-forvar1394));
              reg1425 = wire51[(4'hf):(2'h2)];
              reg1426 = ((8'hb1) ^ reg1314[(5'h16):(3'h4)]);
              reg1427 <= $signed($signed(reg1313));
              reg1428 <= wire44;
            end
          else
            begin
              reg1422 = {$unsigned($unsigned(reg1401[(1'h1):(1'h0)])),
                  {$unsigned(((^wire44) ?
                          (forvar1394 ? reg1406 : reg1428) : $signed(reg1402))),
                      (wire50 + (reg1348[(2'h3):(2'h3)] ?
                          (~^reg1408) : $unsigned(reg1304))),
                      (($signed(reg1419) << reg1420) ?
                          {reg1383[(2'h3):(2'h3)],
                              (reg1425 ? reg1359 : forvar1415),
                              reg1398[(1'h0):(1'h0)]} : (~{reg1397,
                              reg1425}))}};
              reg1423 = ($unsigned($signed(forvar1412[(4'h9):(3'h7)])) ?
                  reg1383[(5'h11):(2'h3)] : (reg1315[(2'h3):(1'h0)] >> (reg1386 ?
                      reg1304[(1'h0):(1'h0)] : reg1371)));
              reg1425 = reg1409[(2'h2):(1'h0)];
              reg1426 = forvar1405[(2'h3):(2'h2)];
              reg1427 <= (-(~|forvar1394[(3'h4):(3'h4)]));
              reg1428 <= reg1411[(2'h3):(2'h2)];
              reg1429 <= $signed(forvar1402);
            end
        end
    end
  assign wire1430 = reg1298[(5'h1d):(5'h1a)];
  assign wire1431 = (|$unsigned(reg1408));
  assign wire1432 = (reg1399 != reg1400[(4'h9):(2'h3)]);
  module1433 #() modinst2442 (wire2441, clk, reg1368, reg1286, wire48, reg1387, reg1319, reg1344);
  assign wire2443 = reg1363;
  always
    @(posedge clk) begin
      reg2444 = reg1351;
      reg2445 = reg1363[(3'h7):(2'h2)];
      reg2446 = {reg1408[(1'h0):(1'h0)], reg2445};
      reg2447 <= reg1424[(3'h4):(2'h2)];
    end
  assign wire2448 = (|reg1290);
  assign wire2449 = $unsigned(($signed((reg1312 ?
                        $signed(reg1355) : (~|wire2441))) >= $unsigned($signed((reg1275 + reg1399)))));
  assign wire2450 = reg1313[(5'h15):(5'h12)];
  assign wire2451 = (reg1319[(4'h9):(3'h6)] < {$signed((reg1368[(2'h2):(2'h2)] ?
                            reg1281[(4'hc):(4'hc)] : wire1431[(1'h0):(1'h0)]))});
  assign wire2452 = $unsigned((+($unsigned($unsigned(reg1401)) <= $unsigned(wire46[(3'h7):(3'h6)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1433
#(parameter param2439 = ((~|((|(~(8'hb9))) & ((+(7'h4f)) ? (!(7'h45)) : (-(8'hb5))))) >= {({((7'h57) << (8'hbc)), {(8'ha0)}} >> (8'h9f))}), 
parameter param2440 = param2439)
(y, clk, wire1439, wire1438, wire1437, wire1436, wire1435, wire1434);
  output wire [(32'h1b3d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire1439;
  input wire [(5'h1b):(1'h0)] wire1438;
  input wire signed [(4'ha):(1'h0)] wire1437;
  input wire [(5'h1d):(1'h0)] wire1436;
  input wire [(5'h1f):(1'h0)] wire1435;
  input wire signed [(5'h1c):(1'h0)] wire1434;
  wire signed [(5'h16):(1'h0)] wire2438;
  wire signed [(5'h12):(1'h0)] wire2437;
  wire [(5'h15):(1'h0)] wire2436;
  wire [(3'h5):(1'h0)] wire2326;
  wire [(5'h1f):(1'h0)] wire2324;
  wire signed [(5'h1a):(1'h0)] wire2323;
  wire signed [(4'ha):(1'h0)] wire2321;
  wire [(5'h1e):(1'h0)] wire1906;
  wire [(4'hc):(1'h0)] wire1685;
  wire signed [(5'h13):(1'h0)] wire1684;
  wire signed [(3'h5):(1'h0)] wire1566;
  wire [(5'h1f):(1'h0)] wire1565;
  reg [(5'h10):(1'h0)] reg2432 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2431 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2427 = (1'h0);
  reg [(3'h7):(1'h0)] reg2423 = (1'h0);
  reg [(5'h11):(1'h0)] reg2422 = (1'h0);
  reg [(5'h18):(1'h0)] reg2421 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2418 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2417 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2416 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2413 = (1'h0);
  reg [(5'h16):(1'h0)] reg2412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2408 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2407 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2403 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2402 = (1'h0);
  reg [(5'h16):(1'h0)] reg2399 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2397 = (1'h0);
  reg [(4'he):(1'h0)] reg2396 = (1'h0);
  reg [(3'h6):(1'h0)] reg2395 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2391 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2389 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2388 = (1'h0);
  reg [(4'hd):(1'h0)] reg2385 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2384 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2382 = (1'h0);
  reg [(5'h10):(1'h0)] reg2375 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2374 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2371 = (1'h0);
  reg [(4'he):(1'h0)] reg2365 = (1'h0);
  reg [(5'h15):(1'h0)] reg2363 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2361 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2357 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2355 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2351 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2349 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2348 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2345 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2341 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2340 = (1'h0);
  reg [(5'h11):(1'h0)] reg2337 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2330 = (1'h0);
  reg [(5'h11):(1'h0)] reg2328 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2327 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2325 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1681 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1676 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1675 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1674 = (1'h0);
  reg [(5'h14):(1'h0)] reg1673 = (1'h0);
  reg [(5'h17):(1'h0)] reg1672 = (1'h0);
  reg [(4'he):(1'h0)] reg1670 = (1'h0);
  reg [(5'h19):(1'h0)] reg1668 = (1'h0);
  reg [(4'h9):(1'h0)] reg1667 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1666 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1663 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1661 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1659 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1658 = (1'h0);
  reg [(5'h19):(1'h0)] reg1657 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1651 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1647 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1645 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1644 = (1'h0);
  reg [(5'h12):(1'h0)] reg1642 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1636 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1633 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1630 = (1'h0);
  reg [(4'h9):(1'h0)] reg1628 = (1'h0);
  reg [(4'hf):(1'h0)] reg1626 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1625 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1624 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1623 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1621 = (1'h0);
  reg [(5'h10):(1'h0)] reg1618 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1617 = (1'h0);
  reg [(3'h6):(1'h0)] reg1611 = (1'h0);
  reg [(2'h2):(1'h0)] reg1608 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1602 = (1'h0);
  reg [(2'h3):(1'h0)] reg1601 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1600 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1599 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1596 = (1'h0);
  reg [(4'ha):(1'h0)] reg1594 = (1'h0);
  reg [(3'h5):(1'h0)] reg1593 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1592 = (1'h0);
  reg [(3'h5):(1'h0)] reg1587 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1585 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1584 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1567 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1582 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1581 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1578 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1576 = (1'h0);
  reg [(5'h10):(1'h0)] reg1572 = (1'h0);
  reg [(5'h10):(1'h0)] reg1569 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1568 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1564 = (1'h0);
  reg [(5'h18):(1'h0)] reg1561 = (1'h0);
  reg [(3'h4):(1'h0)] reg1559 = (1'h0);
  reg [(4'ha):(1'h0)] reg1557 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1554 = (1'h0);
  reg [(5'h15):(1'h0)] reg1551 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1550 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1549 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1548 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1546 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1545 = (1'h0);
  reg [(5'h18):(1'h0)] reg1541 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1539 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1538 = (1'h0);
  reg [(4'ha):(1'h0)] reg1537 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1536 = (1'h0);
  reg [(4'he):(1'h0)] reg1533 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1530 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1528 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1522 = (1'h0);
  reg [(3'h4):(1'h0)] reg1521 = (1'h0);
  reg [(5'h15):(1'h0)] reg1517 = (1'h0);
  reg [(4'ha):(1'h0)] reg1512 = (1'h0);
  reg [(4'h8):(1'h0)] reg1510 = (1'h0);
  reg [(5'h10):(1'h0)] reg1508 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1505 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1503 = (1'h0);
  reg [(5'h15):(1'h0)] reg1502 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1501 = (1'h0);
  reg [(4'ha):(1'h0)] reg1499 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1498 = (1'h0);
  reg [(4'h9):(1'h0)] reg1496 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1495 = (1'h0);
  reg [(3'h4):(1'h0)] reg1494 = (1'h0);
  reg [(5'h19):(1'h0)] reg1492 = (1'h0);
  reg [(4'h9):(1'h0)] reg1491 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1489 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1486 = (1'h0);
  reg [(5'h19):(1'h0)] reg1484 = (1'h0);
  reg [(5'h13):(1'h0)] reg1477 = (1'h0);
  reg [(5'h10):(1'h0)] reg1476 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1473 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1472 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1470 = (1'h0);
  reg [(2'h3):(1'h0)] reg1469 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1464 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1463 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1460 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1459 = (1'h0);
  reg [(5'h10):(1'h0)] reg1457 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1456 = (1'h0);
  reg [(5'h15):(1'h0)] reg1455 = (1'h0);
  reg [(2'h3):(1'h0)] reg1452 = (1'h0);
  reg [(5'h12):(1'h0)] reg1450 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1449 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1447 = (1'h0);
  reg [(4'ha):(1'h0)] reg1446 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1445 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1444 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1442 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1441 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1910 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1911 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1915 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1916 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1918 = (1'h0);
  reg [(3'h6):(1'h0)] reg1919 = (1'h0);
  reg [(3'h4):(1'h0)] reg1920 = (1'h0);
  reg [(4'hd):(1'h0)] reg1925 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1927 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1928 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1930 = (1'h0);
  reg [(5'h17):(1'h0)] reg1932 = (1'h0);
  reg [(5'h11):(1'h0)] reg1935 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1936 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1938 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1940 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1942 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1948 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1949 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1951 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1952 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1953 = (1'h0);
  reg [(4'ha):(1'h0)] reg1957 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1958 = (1'h0);
  reg [(5'h12):(1'h0)] reg1959 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1960 = (1'h0);
  reg [(3'h6):(1'h0)] reg2435 = (1'h0);
  reg [(5'h16):(1'h0)] reg2434 = (1'h0);
  reg [(5'h14):(1'h0)] reg2433 = (1'h0);
  reg [(4'he):(1'h0)] reg2430 = (1'h0);
  reg [(4'hf):(1'h0)] reg2429 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2428 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2426 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2425 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2424 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2420 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2419 = (1'h0);
  reg [(3'h4):(1'h0)] reg2415 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2414 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2411 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2410 = (1'h0);
  reg [(5'h14):(1'h0)] reg2409 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2406 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2405 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2404 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2401 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2400 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2398 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2394 = (1'h0);
  reg [(4'hb):(1'h0)] reg2393 = (1'h0);
  reg [(5'h16):(1'h0)] reg2392 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2390 = (1'h0);
  reg [(4'hd):(1'h0)] reg2387 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2386 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2383 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2381 = (1'h0);
  reg [(5'h14):(1'h0)] reg2380 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2379 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2378 = (1'h0);
  reg [(4'hc):(1'h0)] reg2377 = (1'h0);
  reg [(5'h13):(1'h0)] reg2376 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2373 = (1'h0);
  reg [(3'h5):(1'h0)] reg2372 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2370 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2369 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2368 = (1'h0);
  reg [(4'hd):(1'h0)] reg2367 = (1'h0);
  reg [(5'h11):(1'h0)] reg2366 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2364 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2362 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2360 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2359 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2358 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2356 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2354 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2353 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2352 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2350 = (1'h0);
  reg [(5'h10):(1'h0)] reg2347 = (1'h0);
  reg [(5'h11):(1'h0)] reg2346 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2344 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2343 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2342 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2339 = (1'h0);
  reg [(5'h17):(1'h0)] reg2338 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2336 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2335 = (1'h0);
  reg [(4'he):(1'h0)] reg2334 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2333 = (1'h0);
  reg [(4'h9):(1'h0)] reg2332 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2327 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2331 = (1'h0);
  reg [(4'hf):(1'h0)] reg2329 = (1'h0);
  reg [(3'h6):(1'h0)] reg1956 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1955 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1954 = (1'h0);
  reg [(3'h6):(1'h0)] reg1950 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1947 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1946 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1945 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1944 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1943 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1941 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1937 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1929 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1939 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1937 = (1'h0);
  reg [(2'h2):(1'h0)] reg1934 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1933 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1931 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1929 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1926 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1924 = (1'h0);
  reg [(5'h19):(1'h0)] reg1923 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1922 = (1'h0);
  reg [(5'h11):(1'h0)] reg1921 = (1'h0);
  reg [(5'h16):(1'h0)] reg1917 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1914 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1913 = (1'h0);
  reg [(4'hb):(1'h0)] reg1912 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1909 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1908 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1683 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1682 = (1'h0);
  reg [(3'h4):(1'h0)] reg1680 = (1'h0);
  reg [(5'h19):(1'h0)] reg1679 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1678 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar1677 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1671 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1669 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1665 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1664 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1662 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1660 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1656 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1655 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1654 = (1'h0);
  reg [(4'hf):(1'h0)] reg1653 = (1'h0);
  reg [(4'ha):(1'h0)] reg1652 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1650 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1649 = (1'h0);
  reg [(5'h14):(1'h0)] reg1648 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1646 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1643 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1641 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1640 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1639 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1638 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1637 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1631 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1628 = (1'h0);
  reg [(3'h7):(1'h0)] reg1627 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1635 = (1'h0);
  reg [(5'h15):(1'h0)] reg1634 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1632 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1631 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1629 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1627 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1622 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1620 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1619 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1616 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1615 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1614 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1613 = (1'h0);
  reg [(3'h5):(1'h0)] reg1612 = (1'h0);
  reg [(5'h12):(1'h0)] reg1610 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1609 = (1'h0);
  reg [(3'h6):(1'h0)] reg1607 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1606 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1605 = (1'h0);
  reg [(4'h8):(1'h0)] reg1604 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1603 = (1'h0);
  reg [(3'h7):(1'h0)] reg1598 = (1'h0);
  reg [(3'h6):(1'h0)] reg1597 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1595 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1591 = (1'h0);
  reg [(3'h6):(1'h0)] reg1590 = (1'h0);
  reg [(4'hb):(1'h0)] reg1589 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1588 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1586 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1583 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1577 = (1'h0);
  reg [(2'h2):(1'h0)] reg1580 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1579 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1577 = (1'h0);
  reg [(5'h18):(1'h0)] reg1575 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1574 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1573 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1571 = (1'h0);
  reg [(3'h7):(1'h0)] reg1570 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1567 = (1'h0);
  reg [(3'h5):(1'h0)] reg1563 = (1'h0);
  reg [(2'h2):(1'h0)] reg1562 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1560 = (1'h0);
  reg [(5'h12):(1'h0)] reg1558 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1556 = (1'h0);
  reg [(4'ha):(1'h0)] reg1555 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1553 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1552 = (1'h0);
  reg [(3'h4):(1'h0)] reg1547 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1544 = (1'h0);
  reg [(4'hf):(1'h0)] reg1543 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1542 = (1'h0);
  reg [(4'hc):(1'h0)] reg1540 = (1'h0);
  reg [(2'h3):(1'h0)] reg1535 = (1'h0);
  reg [(4'ha):(1'h0)] reg1534 = (1'h0);
  reg [(2'h2):(1'h0)] reg1532 = (1'h0);
  reg [(4'h8):(1'h0)] reg1531 = (1'h0);
  reg [(4'ha):(1'h0)] reg1529 = (1'h0);
  reg [(4'h9):(1'h0)] reg1527 = (1'h0);
  reg [(5'h17):(1'h0)] reg1526 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1525 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1524 = (1'h0);
  reg [(4'hc):(1'h0)] reg1523 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1520 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1519 = (1'h0);
  reg [(3'h4):(1'h0)] reg1518 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1516 = (1'h0);
  reg [(4'hf):(1'h0)] reg1515 = (1'h0);
  reg [(5'h10):(1'h0)] reg1514 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1513 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1511 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1509 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1507 = (1'h0);
  reg [(4'hf):(1'h0)] reg1506 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1504 = (1'h0);
  reg [(5'h15):(1'h0)] reg1500 = (1'h0);
  reg [(5'h16):(1'h0)] reg1497 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1493 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1490 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1488 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1487 = (1'h0);
  reg [(3'h5):(1'h0)] reg1485 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1483 = (1'h0);
  reg [(5'h14):(1'h0)] reg1482 = (1'h0);
  reg [(5'h14):(1'h0)] reg1481 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1480 = (1'h0);
  reg [(4'he):(1'h0)] reg1479 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1478 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1475 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1474 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1471 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar1468 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1467 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1466 = (1'h0);
  reg [(5'h14):(1'h0)] reg1465 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1462 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1461 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1458 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1454 = (1'h0);
  reg [(4'hb):(1'h0)] reg1453 = (1'h0);
  reg [(4'hb):(1'h0)] reg1451 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1448 = (1'h0);
  reg [(4'h8):(1'h0)] reg1443 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1440 = (1'h0);
  assign y = {wire2438,
                 wire2437,
                 wire2436,
                 wire2326,
                 wire2324,
                 wire2323,
                 wire2321,
                 wire1906,
                 wire1685,
                 wire1684,
                 wire1566,
                 wire1565,
                 reg2432,
                 reg2431,
                 reg2427,
                 reg2423,
                 reg2422,
                 reg2421,
                 reg2418,
                 reg2417,
                 reg2416,
                 reg2413,
                 reg2412,
                 reg2408,
                 reg2407,
                 reg2403,
                 reg2402,
                 reg2399,
                 reg2397,
                 reg2396,
                 reg2395,
                 reg2391,
                 reg2389,
                 reg2388,
                 reg2385,
                 reg2384,
                 reg2382,
                 reg2375,
                 reg2374,
                 reg2371,
                 reg2365,
                 reg2363,
                 reg2361,
                 reg2357,
                 reg2355,
                 reg2351,
                 reg2349,
                 reg2348,
                 reg2345,
                 reg2341,
                 reg2340,
                 reg2337,
                 reg2330,
                 reg2328,
                 reg2327,
                 reg2325,
                 reg1681,
                 reg1676,
                 reg1675,
                 reg1674,
                 reg1673,
                 reg1672,
                 reg1670,
                 reg1668,
                 reg1667,
                 reg1666,
                 reg1663,
                 reg1661,
                 reg1659,
                 reg1658,
                 reg1657,
                 reg1651,
                 reg1647,
                 reg1645,
                 reg1644,
                 reg1642,
                 reg1636,
                 reg1633,
                 reg1630,
                 reg1628,
                 reg1626,
                 reg1625,
                 reg1624,
                 reg1623,
                 reg1621,
                 reg1618,
                 reg1617,
                 reg1611,
                 reg1608,
                 reg1602,
                 reg1601,
                 reg1600,
                 reg1599,
                 reg1596,
                 reg1594,
                 reg1593,
                 reg1592,
                 reg1587,
                 reg1585,
                 reg1584,
                 reg1567,
                 reg1582,
                 reg1581,
                 reg1578,
                 reg1576,
                 reg1572,
                 reg1569,
                 reg1568,
                 reg1564,
                 reg1561,
                 reg1559,
                 reg1557,
                 reg1554,
                 reg1551,
                 reg1550,
                 reg1549,
                 reg1548,
                 reg1546,
                 reg1545,
                 reg1541,
                 reg1539,
                 reg1538,
                 reg1537,
                 reg1536,
                 reg1533,
                 reg1530,
                 reg1528,
                 reg1522,
                 reg1521,
                 reg1517,
                 reg1512,
                 reg1510,
                 reg1508,
                 reg1505,
                 reg1503,
                 reg1502,
                 reg1501,
                 reg1499,
                 reg1498,
                 reg1496,
                 reg1495,
                 reg1494,
                 reg1492,
                 reg1491,
                 reg1489,
                 reg1486,
                 reg1484,
                 reg1477,
                 reg1476,
                 reg1473,
                 reg1472,
                 reg1470,
                 reg1469,
                 reg1464,
                 reg1463,
                 reg1460,
                 reg1459,
                 reg1457,
                 reg1456,
                 reg1455,
                 reg1452,
                 reg1450,
                 reg1449,
                 reg1447,
                 reg1446,
                 reg1445,
                 reg1444,
                 reg1442,
                 reg1441,
                 reg1910,
                 reg1911,
                 reg1915,
                 reg1916,
                 reg1918,
                 reg1919,
                 reg1920,
                 reg1925,
                 reg1927,
                 reg1928,
                 reg1930,
                 reg1932,
                 reg1935,
                 reg1936,
                 reg1938,
                 reg1940,
                 reg1942,
                 reg1948,
                 reg1949,
                 reg1951,
                 reg1952,
                 reg1953,
                 reg1957,
                 reg1958,
                 reg1959,
                 reg1960,
                 reg2435,
                 reg2434,
                 reg2433,
                 reg2430,
                 reg2429,
                 reg2428,
                 forvar2426,
                 reg2425,
                 forvar2424,
                 reg2420,
                 reg2419,
                 reg2415,
                 forvar2414,
                 reg2411,
                 reg2410,
                 reg2409,
                 forvar2406,
                 reg2405,
                 reg2404,
                 forvar2401,
                 reg2400,
                 reg2398,
                 reg2394,
                 reg2393,
                 reg2392,
                 reg2390,
                 reg2387,
                 reg2386,
                 reg2383,
                 reg2381,
                 reg2380,
                 reg2379,
                 forvar2378,
                 reg2377,
                 reg2376,
                 reg2373,
                 reg2372,
                 reg2370,
                 reg2369,
                 reg2368,
                 reg2367,
                 reg2366,
                 reg2364,
                 reg2362,
                 reg2360,
                 reg2359,
                 reg2358,
                 reg2356,
                 reg2354,
                 reg2353,
                 reg2352,
                 forvar2350,
                 reg2347,
                 reg2346,
                 reg2344,
                 forvar2343,
                 reg2342,
                 reg2339,
                 reg2338,
                 reg2336,
                 forvar2335,
                 reg2334,
                 reg2333,
                 reg2332,
                 forvar2327,
                 reg2331,
                 reg2329,
                 reg1956,
                 reg1955,
                 reg1954,
                 reg1950,
                 reg1947,
                 reg1946,
                 reg1945,
                 reg1944,
                 reg1943,
                 reg1941,
                 reg1937,
                 forvar1929,
                 reg1939,
                 forvar1937,
                 reg1934,
                 reg1933,
                 reg1931,
                 reg1929,
                 reg1926,
                 reg1924,
                 reg1923,
                 reg1922,
                 reg1921,
                 reg1917,
                 reg1914,
                 reg1913,
                 reg1912,
                 reg1909,
                 forvar1908,
                 reg1683,
                 reg1682,
                 reg1680,
                 reg1679,
                 reg1678,
                 forvar1677,
                 reg1671,
                 forvar1669,
                 forvar1665,
                 forvar1664,
                 reg1662,
                 reg1660,
                 reg1656,
                 reg1655,
                 forvar1654,
                 reg1653,
                 reg1652,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1646,
                 forvar1643,
                 forvar1641,
                 reg1640,
                 reg1639,
                 forvar1638,
                 reg1637,
                 reg1631,
                 forvar1628,
                 reg1627,
                 reg1635,
                 reg1634,
                 reg1632,
                 forvar1631,
                 reg1629,
                 forvar1627,
                 reg1622,
                 reg1620,
                 reg1619,
                 reg1616,
                 reg1615,
                 reg1614,
                 reg1613,
                 reg1612,
                 reg1610,
                 forvar1609,
                 reg1607,
                 forvar1606,
                 reg1605,
                 reg1604,
                 forvar1603,
                 reg1598,
                 reg1597,
                 reg1595,
                 reg1591,
                 reg1590,
                 reg1589,
                 reg1588,
                 reg1586,
                 reg1583,
                 forvar1577,
                 reg1580,
                 reg1579,
                 reg1577,
                 reg1575,
                 reg1574,
                 reg1573,
                 reg1571,
                 reg1570,
                 forvar1567,
                 reg1563,
                 reg1562,
                 reg1560,
                 reg1558,
                 reg1556,
                 reg1555,
                 forvar1553,
                 forvar1552,
                 reg1547,
                 forvar1544,
                 reg1543,
                 reg1542,
                 reg1540,
                 reg1535,
                 reg1534,
                 reg1532,
                 reg1531,
                 reg1529,
                 reg1527,
                 reg1526,
                 reg1525,
                 reg1524,
                 reg1523,
                 reg1520,
                 reg1519,
                 reg1518,
                 reg1516,
                 reg1515,
                 reg1514,
                 forvar1513,
                 reg1511,
                 reg1509,
                 forvar1507,
                 reg1506,
                 reg1504,
                 reg1500,
                 reg1497,
                 reg1493,
                 reg1490,
                 forvar1488,
                 reg1487,
                 reg1485,
                 reg1483,
                 reg1482,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1478,
                 reg1475,
                 reg1474,
                 reg1471,
                 forvar1468,
                 reg1467,
                 forvar1466,
                 reg1465,
                 reg1462,
                 reg1461,
                 reg1458,
                 reg1454,
                 reg1453,
                 reg1451,
                 forvar1448,
                 reg1443,
                 forvar1440,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1440 = (1'h0); (forvar1440 < (2'h3)); forvar1440 = (forvar1440 + (1'h1)))
        begin
          reg1441 <= $signed($unsigned(wire1435));
          if ($unsigned((wire1434[(4'h9):(3'h7)] ?
              {{(wire1434 ? wire1436 : wire1434)},
                  wire1437[(4'h9):(3'h5)],
                  ((wire1439 ? wire1439 : wire1439) ?
                      forvar1440[(3'h7):(2'h3)] : (7'h50))} : {(forvar1440 ?
                      {reg1441} : (wire1435 << wire1438)),
                  (^~((8'ha9) ? wire1436 : wire1436))})))
            begin
              reg1442 <= (-(^(-((wire1435 ~^ (8'haa)) & wire1436))));
            end
          else
            begin
              reg1443 = $signed($unsigned($signed(wire1434[(5'h19):(3'h7)])));
              reg1444 <= (7'h51);
              reg1445 <= $unsigned(((((wire1437 <= wire1436) < $signed(reg1444)) ?
                  $unsigned((~^wire1439)) : wire1436[(5'h18):(5'h17)]) <<< {(wire1437[(1'h1):(1'h1)] < (reg1443 ?
                      (8'hba) : reg1441))}));
              reg1446 <= (~&(|$unsigned({forvar1440,
                  $signed(wire1436),
                  reg1443})));
              reg1447 <= $unsigned(($signed((~&(+reg1446))) ?
                  reg1442[(2'h3):(2'h3)] : $signed($signed((reg1446 ?
                      wire1438 : forvar1440)))));
            end
          for (forvar1448 = (1'h0); (forvar1448 < (1'h1)); forvar1448 = (forvar1448 + (1'h1)))
            begin
              reg1449 <= $signed($signed({(+wire1434),
                  ({reg1443, wire1434} ? (~^(8'hb2)) : (!reg1445))}));
              reg1450 <= ($signed(wire1435[(4'h9):(3'h6)]) ?
                  {$unsigned(forvar1440[(3'h7):(2'h3)]),
                      reg1445} : reg1442[(4'ha):(1'h1)]);
              reg1451 = reg1441[(2'h2):(1'h0)];
              reg1452 <= (8'ha0);
              reg1453 = (~&({$unsigned((~|reg1442)),
                  reg1451,
                  (!reg1449)} >= {$signed(((7'h4d) ? wire1437 : forvar1448)),
                  reg1451,
                  (!(7'h53))}));
              reg1454 = $unsigned({(forvar1448 ?
                      (forvar1448 ?
                          reg1451[(4'ha):(4'h8)] : (^~(7'h45))) : ((forvar1440 || wire1435) & (~|reg1453))),
                  (reg1451[(2'h3):(2'h3)] ~^ reg1442)});
            end
          if (forvar1440[(5'h12):(4'hc)])
            begin
              reg1455 <= {(^$unsigned($unsigned(reg1454[(4'h8):(2'h3)]))),
                  ((+(wire1435 ? forvar1448 : reg1447[(4'ha):(1'h0)])) ?
                      $signed({((8'hbd) ?
                              wire1439 : reg1442)}) : (+($signed(reg1452) ?
                          $signed(reg1444) : $unsigned((8'hb7))))),
                  ($unsigned(({(8'h9d)} - reg1454[(2'h3):(1'h1)])) << wire1437)};
              reg1456 <= (-(!$signed(reg1442)));
              reg1457 <= wire1434;
            end
          else
            begin
              reg1455 <= {{$signed(($signed(reg1457) ?
                          (reg1447 ~^ wire1436) : reg1454[(4'h9):(3'h6)])),
                      $unsigned(wire1437[(4'h9):(1'h1)]),
                      $signed(reg1443)},
                  reg1454[(2'h3):(1'h0)],
                  $unsigned(reg1455[(4'hd):(2'h3)])};
              reg1458 = wire1436;
              reg1459 <= (8'hbd);
              reg1460 <= ({((wire1439[(5'h11):(1'h0)] || {reg1459}) | (reg1447 ?
                      $signed((8'hb5)) : (reg1459 ? reg1453 : reg1444))),
                  $signed((wire1438[(4'h9):(3'h5)] != reg1457[(4'h8):(1'h1)]))} * (reg1441 != reg1450[(4'hd):(3'h4)]));
              reg1461 = ((reg1450[(3'h5):(1'h0)] ?
                      $signed((~^(reg1444 ?
                          reg1452 : reg1445))) : $unsigned(((wire1438 ?
                              wire1437 : reg1458) ?
                          reg1454 : $unsigned(forvar1440)))) ?
                  (-reg1442[(3'h5):(2'h3)]) : reg1444[(4'hd):(1'h1)]);
              reg1462 = ((reg1454 >= ((8'hba) >>> ($unsigned(reg1460) ^~ (forvar1448 || reg1459)))) > ($signed(reg1459[(4'h8):(1'h0)]) ?
                  {(wire1435[(5'h1e):(5'h16)] ?
                          ((7'h42) ? reg1452 : reg1461) : reg1445),
                      (reg1454[(3'h5):(3'h5)] ?
                          reg1458[(3'h7):(1'h0)] : $unsigned(wire1434))} : reg1443));
              reg1463 <= reg1447[(4'h8):(3'h5)];
            end
          reg1464 <= $signed((reg1463[(3'h4):(2'h2)] ^~ ($signed((^(8'hb4))) ?
              $signed({reg1463}) : $signed(reg1458))));
          reg1465 = wire1435[(4'hf):(4'hd)];
        end
      for (forvar1466 = (1'h0); (forvar1466 < (1'h0)); forvar1466 = (forvar1466 + (1'h1)))
        begin
          reg1467 = reg1452;
        end
      for (forvar1468 = (1'h0); (forvar1468 < (2'h3)); forvar1468 = (forvar1468 + (1'h1)))
        begin
          reg1469 <= ((&wire1438[(5'h19):(4'hd)]) ?
              {(8'h9e),
                  ($signed($unsigned(reg1456)) ?
                      (^~$unsigned(reg1451)) : $unsigned((8'haf))),
                  ($unsigned((forvar1440 || (7'h55))) ?
                      (|reg1459[(3'h4):(1'h0)]) : (^~reg1467))} : reg1453);
          if (reg1450)
            begin
              reg1470 <= reg1445;
              reg1471 = reg1465;
              reg1472 <= (^~$unsigned((reg1446 >= (forvar1468[(5'h19):(5'h13)] ?
                  reg1471 : (wire1439 ? reg1445 : reg1457)))));
              reg1473 <= $signed(reg1445);
              reg1474 = ($signed($signed(reg1453)) ^ $signed((($signed(reg1461) ?
                      (!reg1450) : ((7'h55) < (8'hbb))) ?
                  $unsigned((reg1470 ?
                      reg1458 : (7'h54))) : forvar1466[(2'h3):(2'h3)])));
            end
          else
            begin
              reg1470 <= (reg1464[(5'h1b):(4'hc)] ?
                  (((((7'h44) > (8'hb8)) ?
                          (wire1435 ? reg1446 : wire1438) : (reg1458 ?
                              reg1474 : reg1445)) ?
                      $signed((+wire1436)) : $signed((reg1471 ~^ reg1461))) > ($signed($signed(reg1474)) ?
                      {$unsigned(reg1464),
                          $signed((7'h4a)),
                          (reg1472 ?
                              reg1453 : reg1445)} : $unsigned($signed((8'hb7))))) : ({reg1458} - $signed(((8'hb4) >= reg1465))));
              reg1471 = reg1464;
              reg1474 = reg1442;
              reg1475 = reg1441[(3'h6):(2'h2)];
            end
          reg1476 <= {((reg1470 ? (~|reg1450) : {(reg1464 <<< reg1441)}) ?
                  reg1456[(2'h2):(1'h1)] : (reg1454[(4'h9):(1'h0)] * (reg1474[(2'h3):(2'h2)] ?
                      (&reg1464) : $signed(reg1460)))),
              $signed(reg1462[(5'h12):(4'h9)]),
              $unsigned((^(8'had)))};
          reg1477 <= ($signed(reg1442[(1'h0):(1'h0)]) > ((~^reg1467[(2'h3):(1'h0)]) ?
              reg1441[(3'h6):(1'h0)] : $signed($signed($signed(reg1450)))));
          reg1478 = {(reg1453[(3'h6):(2'h3)] ?
                  (~|{(reg1458 ? reg1470 : reg1441),
                      reg1443,
                      $signed(reg1477)}) : (^($unsigned(forvar1466) ?
                      reg1462 : (reg1463 <= forvar1448))))};
          if ({$unsigned(wire1436[(4'hd):(4'hc)]),
              (~$signed((8'hb1))),
              reg1460})
            begin
              reg1479 = {((-($signed(wire1437) || (8'hac))) ?
                      reg1464 : reg1449[(4'ha):(1'h1)])};
              reg1480 = $signed(($unsigned((((8'h9c) >= forvar1448) ?
                      (8'haf) : (reg1469 ? reg1454 : (8'hbf)))) ?
                  (~&{(8'hb8), {forvar1448}}) : {reg1477[(5'h10):(5'h10)],
                      ((~|reg1464) ~^ (7'h40)),
                      $signed($signed(reg1457))}));
              reg1481 = (!($signed((~{wire1436})) ^~ $unsigned(reg1451)));
              reg1482 = ((-reg1452[(1'h0):(1'h0)]) ?
                  (~^forvar1440[(4'hd):(1'h0)]) : {((reg1450[(5'h10):(3'h6)] > reg1470) ?
                          (|(^~reg1456)) : reg1445),
                      $unsigned(((reg1457 ? reg1455 : reg1447) ?
                          reg1449 : $signed(reg1462)))});
              reg1483 = (forvar1468 <= (reg1479[(4'hb):(1'h0)] <= {(reg1481 ?
                      reg1453 : (!(7'h46)))}));
              reg1484 <= reg1464[(5'h1e):(4'h9)];
              reg1485 = (&reg1443[(3'h5):(3'h5)]);
            end
          else
            begin
              reg1479 = $unsigned(reg1469);
              reg1484 <= reg1458;
              reg1486 <= (!(~^(reg1447[(3'h6):(3'h4)] ?
                  ($unsigned(reg1485) & (reg1483 ?
                      (8'ha1) : reg1449)) : (~^(reg1453 ?
                      reg1453 : reg1477)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg1487 = ((wire1437[(3'h5):(3'h4)] ?
          reg1447[(3'h5):(3'h4)] : (({wire1436, wire1434, reg1464} ?
                  $unsigned(reg1472) : (reg1455 ? wire1439 : reg1460)) ?
              (-$signed(reg1459)) : ((~wire1435) ?
                  $signed(reg1442) : (wire1435 ?
                      reg1473 : reg1447)))) >>> ($signed(((~^(8'hb9)) ?
              $signed(reg1447) : reg1455[(4'hd):(3'h7)])) ?
          (reg1456 ?
              $unsigned((reg1486 ?
                  (7'h53) : reg1472)) : {(-reg1486)}) : $unsigned(reg1446[(3'h4):(2'h2)])));
      for (forvar1488 = (1'h0); (forvar1488 < (3'h4)); forvar1488 = (forvar1488 + (1'h1)))
        begin
          reg1489 <= (^reg1487[(3'h5):(1'h0)]);
          if ({{$unsigned($signed((7'h50)))},
              (($unsigned(((8'hbf) ?
                  wire1436 : reg1457)) && reg1469[(2'h2):(2'h2)]) > ($signed(reg1445[(4'ha):(1'h1)]) ?
                  (reg1444[(5'h19):(5'h15)] ?
                      (^wire1438) : (forvar1488 != wire1438)) : (reg1442[(3'h4):(1'h1)] ?
                      $unsigned(reg1484) : (-reg1456))))})
            begin
              reg1490 = $unsigned($unsigned(reg1446[(3'h5):(3'h4)]));
              reg1491 <= (wire1437[(3'h6):(2'h3)] & ((+((~|reg1459) ?
                  $signed(wire1435) : (^~wire1439))) == {((reg1457 ^~ reg1484) <<< ((7'h47) ?
                      reg1472 : (7'h43)))}));
              reg1492 <= (-((!($unsigned(reg1484) > {reg1490, reg1486})) ?
                  (reg1446[(1'h0):(1'h0)] ?
                      $unsigned(reg1490[(2'h2):(1'h1)]) : (8'hb6)) : reg1464));
              reg1493 = $signed(reg1456[(2'h2):(2'h2)]);
              reg1494 <= ((7'h4b) ?
                  reg1492[(3'h7):(1'h1)] : $signed((reg1487[(1'h1):(1'h1)] <<< {reg1484})));
            end
          else
            begin
              reg1490 = ((reg1457[(1'h0):(1'h0)] != (((8'hb7) ?
                      reg1490[(1'h0):(1'h0)] : $signed(reg1491)) ?
                  ((reg1442 > (7'h4d)) ?
                      $unsigned(wire1436) : (reg1455 ?
                          reg1441 : reg1476)) : {(|(8'ha8)),
                      $unsigned(reg1476)})) | reg1472[(3'h7):(3'h4)]);
              reg1493 = ($unsigned(({reg1492, (reg1446 - reg1494)} ?
                  {$signed(reg1492),
                      reg1441,
                      $unsigned(reg1459)} : ((&reg1476) ?
                      reg1456[(1'h0):(1'h0)] : (reg1452 ~^ reg1455)))) <= {$signed($signed($signed(reg1491)))});
            end
          reg1495 <= $unsigned(wire1439[(3'h7):(3'h7)]);
          reg1496 <= $signed($unsigned($unsigned(($signed(reg1494) ?
              (|(7'h42)) : {reg1444, wire1434, reg1455}))));
        end
      if ($signed(reg1494))
        begin
          reg1497 = ($unsigned({(~&$unsigned(reg1496)),
              (7'h55)}) > (~&(((7'h51) ~^ $unsigned(reg1441)) & (reg1442[(4'hd):(4'hc)] ?
              (reg1490 >>> reg1470) : reg1476[(2'h2):(1'h1)]))));
        end
      else
        begin
          reg1498 <= (~(wire1439 < $signed(({wire1434} ~^ $unsigned((8'had))))));
          if (reg1469)
            begin
              reg1499 <= reg1486;
              reg1500 = $unsigned($unsigned({$signed({reg1493, reg1447}),
                  $signed($signed(reg1442)),
                  (^(^reg1470))}));
              reg1501 <= (^(8'ha3));
              reg1502 <= $signed((&$unsigned($signed((+reg1492)))));
              reg1503 <= $unsigned((reg1441 ?
                  (!reg1460) : {(reg1469 ^~ $signed((8'hb9))),
                      ({wire1439, (7'h45)} ? $unsigned(reg1498) : reg1459)}));
              reg1504 = (&$unsigned($signed(((reg1477 ? reg1495 : reg1464) ?
                  (^~reg1446) : $unsigned(reg1502)))));
              reg1505 <= $signed(((reg1472[(5'h11):(3'h7)] && (^~{reg1464})) ?
                  reg1487[(1'h0):(1'h0)] : $unsigned($unsigned($signed(reg1504)))));
            end
          else
            begin
              reg1500 = $signed({reg1486, (~|$signed($unsigned(reg1457)))});
              reg1501 <= (-$signed($signed($unsigned(reg1497))));
              reg1502 <= $signed($unsigned(reg1472));
              reg1504 = reg1505;
              reg1506 = ($signed($unsigned(($signed(reg1459) ^ $signed(reg1469)))) ?
                  {(((|(7'h47)) ? $unsigned(reg1442) : reg1489) ?
                          {reg1496, {(8'ha2)}} : (7'h56)),
                      reg1493} : reg1470[(5'h16):(5'h14)]);
            end
          for (forvar1507 = (1'h0); (forvar1507 < (2'h3)); forvar1507 = (forvar1507 + (1'h1)))
            begin
              reg1508 <= reg1494;
              reg1509 = reg1484[(3'h4):(1'h0)];
              reg1510 <= ($signed(reg1486[(1'h0):(1'h0)]) ?
                  $unsigned(($unsigned((reg1504 ?
                      wire1438 : reg1456)) || reg1505[(5'h19):(4'hd)])) : ($unsigned(reg1489) ?
                      ((^$signed((8'hbb))) ?
                          $unsigned(reg1477) : ((reg1477 - (8'hb9)) ?
                              (reg1509 <<< reg1445) : $unsigned(reg1503))) : ({wire1437,
                          (~|(8'hb9))} * $signed((!reg1442)))));
              reg1511 = (7'h4a);
              reg1512 <= $signed({$signed(((-reg1503) ?
                      $signed(reg1504) : (reg1442 ? reg1441 : reg1455))),
                  reg1470[(5'h10):(1'h1)]});
            end
          for (forvar1513 = (1'h0); (forvar1513 < (1'h1)); forvar1513 = (forvar1513 + (1'h1)))
            begin
              reg1514 = wire1437[(3'h5):(1'h1)];
              reg1515 = $signed((8'had));
              reg1516 = reg1484[(4'h9):(3'h4)];
            end
          if ({$signed(((!((8'hac) ?
                  reg1484 : reg1441)) <= reg1514[(4'h8):(3'h4)]))})
            begin
              reg1517 <= ((reg1486[(4'h9):(3'h4)] << (~^$unsigned($signed(reg1505)))) + $signed(reg1505[(5'h12):(4'hb)]));
              reg1518 = reg1450;
              reg1519 = $signed((^~reg1464[(4'hf):(4'hf)]));
              reg1520 = (^$signed({({reg1464,
                      (8'hab),
                      reg1515} <= (~^reg1477))}));
            end
          else
            begin
              reg1517 <= $signed($signed(reg1514));
              reg1521 <= reg1496[(3'h6):(3'h4)];
              reg1522 <= (8'ha1);
              reg1523 = reg1515;
              reg1524 = ($signed($unsigned(($signed(reg1519) - $signed(reg1512)))) ?
                  $signed($unsigned(({reg1508, reg1506, reg1442} ?
                      (8'ha6) : reg1520[(1'h1):(1'h1)]))) : ((8'hb4) ?
                      (8'hae) : $unsigned(reg1494[(2'h2):(1'h0)])));
              reg1525 = $signed(($signed($unsigned((reg1464 ?
                      forvar1513 : reg1489))) ?
                  $unsigned(reg1502[(4'ha):(4'ha)]) : ($signed(reg1457) ?
                      $unsigned((wire1436 == reg1512)) : reg1441[(2'h3):(2'h3)])));
              reg1526 = reg1494[(2'h2):(2'h2)];
            end
          if ({($unsigned($unsigned(reg1442)) ?
                  $signed(reg1502[(5'h11):(4'h8)]) : {$signed((reg1521 <= reg1441))}),
              $signed(reg1469),
              reg1455[(4'h8):(1'h1)]})
            begin
              reg1527 = (($signed(($unsigned((8'ha5)) != (reg1487 || reg1495))) < $unsigned((((8'hb8) ?
                          reg1469 : reg1518) ?
                      {reg1486} : (reg1515 ? reg1512 : reg1446)))) ?
                  $signed($signed($signed((&reg1442)))) : $signed(((|((8'hb7) ?
                      reg1519 : reg1446)) != $signed((reg1489 << reg1473)))));
              reg1528 <= reg1491;
              reg1529 = {reg1506[(4'hb):(3'h7)]};
            end
          else
            begin
              reg1527 = $unsigned(((7'h4d) >> (((reg1505 >> reg1521) ?
                      (~^(7'h4a)) : {reg1452}) ?
                  {$unsigned(reg1497)} : (!reg1487))));
              reg1528 <= {$unsigned({wire1436, reg1508[(4'h8):(1'h1)]}),
                  ($unsigned($signed($unsigned(reg1464))) ?
                      {(8'hb9),
                          {(reg1499 ? wire1436 : reg1490),
                              {reg1469}}} : (reg1527[(4'h9):(2'h2)] <= (|(!reg1493)))),
                  reg1514};
              reg1530 <= reg1508[(4'hd):(3'h6)];
              reg1531 = $unsigned(reg1490);
              reg1532 = ((~&reg1460) + $unsigned((-$unsigned(reg1460))));
            end
          if (reg1463)
            begin
              reg1533 <= reg1457;
              reg1534 = $signed(reg1519[(5'h13):(5'h13)]);
              reg1535 = {reg1459};
              reg1536 <= $unsigned(reg1497);
              reg1537 <= ({($unsigned(((8'ha6) ^ reg1506)) && ($signed(reg1476) >= reg1452[(1'h1):(1'h1)])),
                      ((reg1525[(5'h18):(4'h8)] >>> $unsigned(reg1442)) ?
                          wire1439 : $unsigned(reg1446))} ?
                  (^~(~&reg1490)) : reg1504[(4'hf):(4'hb)]);
              reg1538 <= ((^($signed(reg1464) ?
                      ((wire1439 >> wire1434) ?
                          reg1509[(5'h10):(4'ha)] : forvar1488[(3'h5):(2'h2)]) : ($unsigned(reg1457) ?
                          {(8'h9f), reg1444, reg1533} : (!reg1524)))) ?
                  $unsigned((((^~reg1510) ^ (^reg1516)) ?
                      ((~&reg1501) ?
                          (7'h53) : reg1449) : reg1533)) : $signed({(reg1493[(4'hb):(2'h3)] <<< $unsigned(reg1473)),
                      reg1460[(5'h13):(1'h1)],
                      reg1498}));
              reg1539 <= $signed($signed((((~|reg1503) ?
                  $signed((8'hb0)) : (|reg1450)) & $unsigned(reg1522[(2'h3):(2'h3)]))));
            end
          else
            begin
              reg1533 <= $signed({(reg1509 >> wire1437),
                  reg1529[(3'h4):(1'h1)],
                  (&$unsigned(reg1516[(4'hc):(3'h6)]))});
              reg1536 <= (7'h54);
              reg1540 = reg1498;
              reg1541 <= $signed((+$unsigned((reg1456 * (|reg1486)))));
            end
        end
      reg1542 = $unsigned($unsigned(((reg1489 ?
              $unsigned((8'ha0)) : $signed(reg1501)) ?
          $unsigned((reg1490 || reg1477)) : reg1449)));
    end
  always
    @(posedge clk) begin
      reg1543 = ((^$unsigned($unsigned($signed(reg1537)))) >> ($unsigned($unsigned(reg1498[(1'h0):(1'h0)])) ?
          (^~$unsigned(((7'h58) ~^ (8'hb6)))) : (~reg1528)));
      for (forvar1544 = (1'h0); (forvar1544 < (3'h5)); forvar1544 = (forvar1544 + (1'h1)))
        begin
          reg1545 <= (({reg1539[(5'h13):(4'hc)]} >> $signed(reg1464[(5'h14):(2'h2)])) ?
              (reg1445 ?
                  ((((8'hbc) << (7'h55)) < (reg1484 ?
                      (8'ha1) : reg1456)) * (reg1539[(5'h19):(3'h4)] | $signed(wire1438))) : {reg1469,
                      (7'h44)}) : reg1442[(4'hf):(4'h8)]);
          reg1546 <= reg1464[(4'he):(3'h4)];
          reg1547 = $signed($unsigned($unsigned((~^(reg1457 && reg1546)))));
          reg1548 <= $unsigned($signed($signed($unsigned(reg1450[(4'h8):(3'h4)]))));
          reg1549 <= (-reg1463);
          reg1550 <= (~|{reg1456[(2'h2):(2'h2)],
              {(((8'haa) ~^ reg1452) - reg1512)},
              {reg1457[(3'h4):(3'h4)],
                  reg1447[(4'ha):(4'ha)],
                  ($unsigned(reg1522) != $signed(reg1510))}});
          reg1551 <= $unsigned(reg1502);
        end
      for (forvar1552 = (1'h0); (forvar1552 < (3'h6)); forvar1552 = (forvar1552 + (1'h1)))
        begin
          for (forvar1553 = (1'h0); (forvar1553 < (3'h6)); forvar1553 = (forvar1553 + (1'h1)))
            begin
              reg1554 <= $signed((reg1469[(2'h2):(1'h1)] ?
                  $signed($unsigned($signed(reg1496))) : reg1457[(4'hf):(4'hf)]));
              reg1555 = ($signed(($signed((&reg1446)) ?
                      $signed($signed(reg1528)) : $signed(wire1436[(3'h4):(2'h2)]))) ?
                  (((!(wire1435 ? (8'hbe) : reg1501)) ?
                      (^$signed(reg1445)) : reg1469) ~^ (({reg1473,
                              (7'h55),
                              reg1486} ?
                          reg1484 : reg1441[(2'h3):(1'h1)]) ?
                      $unsigned({reg1444,
                          reg1543}) : {reg1455[(4'h8):(3'h4)]})) : reg1537[(2'h3):(1'h0)]);
              reg1556 = ($signed($unsigned($unsigned((reg1496 ?
                  reg1505 : wire1438)))) >= (&(($signed(reg1522) > (~reg1537)) ?
                  (8'haf) : reg1464)));
              reg1557 <= (8'h9e);
              reg1558 = (((reg1536[(2'h2):(1'h0)] >>> (((8'ha1) == reg1508) >>> (reg1554 ?
                      (7'h4e) : reg1441))) ?
                  reg1555[(4'h8):(1'h0)] : (~|($signed(forvar1544) | reg1442))) ~^ reg1452[(2'h3):(1'h1)]);
              reg1559 <= reg1551;
              reg1560 = $signed($signed(reg1489[(2'h2):(1'h0)]));
            end
        end
      reg1561 <= {$unsigned($signed((~^reg1548[(4'ha):(4'h9)]))),
          $unsigned((~((|reg1510) ? ((8'hb6) != reg1486) : reg1503))),
          reg1558[(3'h6):(1'h0)]};
      reg1562 = reg1459;
      reg1563 = reg1459;
    end
  always
    @(posedge clk) begin
      reg1564 <= $unsigned(reg1459[(4'ha):(3'h4)]);
    end
  assign wire1565 = ((reg1505[(4'h8):(3'h7)] ~^ (^((8'hb8) >= ((8'hb0) ?
                        wire1434 : reg1498)))) > ({($unsigned(reg1469) ?
                            wire1435[(5'h17):(3'h6)] : wire1438[(5'h11):(3'h7)]),
                        ($unsigned(reg1442) <= (reg1557 ? reg1442 : reg1528)),
                        ((reg1441 && reg1476) ?
                            $signed(reg1538) : reg1530[(5'h12):(4'hc)])} & $signed(reg1551)));
  assign wire1566 = (((((reg1521 ? reg1521 : reg1539) ^ (reg1491 >> reg1550)) ?
                        reg1521 : (reg1548 == reg1495)) - reg1491) <<< (((~&$unsigned((8'hb7))) && reg1545) ?
                        $signed(reg1517[(5'h10):(1'h1)]) : wire1438[(3'h6):(2'h2)]));
  always
    @(posedge clk) begin
      if (reg1460[(4'hb):(3'h6)])
        begin
          for (forvar1567 = (1'h0); (forvar1567 < (3'h6)); forvar1567 = (forvar1567 + (1'h1)))
            begin
              reg1568 <= (^{{reg1536},
                  ($signed({reg1470, reg1551}) ? reg1545 : wire1437)});
              reg1569 <= reg1537[(1'h0):(1'h0)];
            end
          if (($signed($unsigned($unsigned(reg1463))) ?
              $signed((&(8'ha7))) : reg1473))
            begin
              reg1570 = ($signed(reg1512) ~^ reg1537);
            end
          else
            begin
              reg1570 = $signed((+((~$signed(reg1470)) ?
                  (wire1438[(5'h15):(3'h7)] ?
                      wire1566 : $signed(reg1521)) : forvar1567[(1'h0):(1'h0)])));
              reg1571 = $unsigned(((({wire1434} > (reg1554 <= (8'hb6))) ?
                      reg1517 : ((-reg1486) ?
                          (reg1528 ? reg1457 : (8'h9f)) : (wire1436 ?
                              wire1566 : reg1550))) ?
                  $unsigned(($unsigned(reg1536) ?
                      ((8'hb4) ?
                          reg1496 : (7'h4d)) : (8'haa))) : (~&reg1491[(2'h2):(1'h1)])));
            end
          reg1572 <= $unsigned($signed((^~reg1549[(4'hc):(4'h8)])));
          reg1573 = ($unsigned($unsigned((~$unsigned(reg1522)))) ?
              $signed({$signed(reg1550[(5'h11):(4'h8)]),
                  $unsigned(reg1449)}) : (~^$unsigned(($signed(reg1447) ?
                  $signed(wire1436) : reg1501))));
          if ((-$signed((reg1494 ?
              (^~reg1452) : ($signed(reg1450) <= (reg1457 >> (8'hb5)))))))
            begin
              reg1574 = (^~$signed((^~{reg1470[(4'he):(1'h0)]})));
              reg1575 = (($unsigned({(-reg1445)}) ?
                  $signed({reg1559}) : $unsigned(reg1559)) | reg1447);
              reg1576 <= $unsigned(({((reg1533 < reg1501) ?
                          $signed(reg1536) : (reg1446 ? reg1541 : reg1557)),
                      ($signed(reg1477) && $unsigned(reg1494))} ?
                  (-((reg1533 && reg1545) >>> {reg1463,
                      wire1566,
                      reg1537})) : {{$unsigned(reg1503)}}));
              reg1577 = (~&((({reg1469, (8'hbd)} | (^reg1546)) ?
                  (|(reg1561 ?
                      (8'hb9) : reg1492)) : (!((8'hba) != reg1533))) <<< (~|wire1435[(2'h3):(1'h0)])));
              reg1578 <= ({(((reg1492 < (8'ha2)) ^ (wire1566 ?
                          reg1549 : reg1539)) ?
                      {(~&reg1503)} : reg1564)} << (reg1551[(5'h14):(3'h6)] ?
                  reg1495[(5'h14):(4'hf)] : ((!(reg1530 ? (8'hb9) : reg1510)) ?
                      $signed({wire1566,
                          (7'h54),
                          reg1551}) : ($unsigned(reg1548) <<< $unsigned(reg1539)))));
              reg1579 = $unsigned(reg1578[(2'h2):(1'h0)]);
              reg1580 = $unsigned((((!(~reg1455)) ?
                      $unsigned((~&reg1576)) : reg1561[(4'hc):(4'h9)]) ?
                  reg1561[(5'h14):(4'hd)] : {$unsigned(((8'haf) ?
                          reg1449 : reg1578))}));
            end
          else
            begin
              reg1574 = reg1464;
              reg1576 <= reg1444[(5'h1b):(5'h15)];
              reg1578 <= {reg1457[(3'h7):(2'h2)]};
              reg1581 <= $signed({(reg1442[(1'h1):(1'h1)] ?
                      (-reg1569) : reg1470[(1'h0):(1'h0)]),
                  $signed((!$unsigned(reg1546))),
                  $signed((reg1477 ^~ $signed(wire1566)))});
              reg1582 <= $signed(reg1472[(4'hc):(3'h5)]);
            end
        end
      else
        begin
          reg1567 <= reg1573;
          reg1570 = (-$signed((wire1435 ?
              reg1444 : ($unsigned(reg1464) * reg1503))));
          if (((reg1486 ? reg1551 : reg1495[(5'h14):(5'h11)]) ?
              (reg1579 ?
                  reg1472[(1'h1):(1'h1)] : reg1486) : ((reg1580 * (reg1464 >> reg1498)) ?
                  reg1457 : (^~($unsigned((8'hbc)) ?
                      (reg1557 ? reg1579 : reg1492) : $signed(reg1445))))))
            begin
              reg1572 <= $signed($signed(($signed($unsigned((8'hb9))) - (~^reg1548))));
              reg1573 = $signed((~|$signed($signed($unsigned(reg1460)))));
              reg1576 <= ({reg1455[(3'h5):(1'h0)],
                      $signed(reg1459),
                      ($signed((~(7'h52))) ?
                          reg1445[(1'h1):(1'h1)] : $signed((^~(8'ha2))))} ?
                  {(reg1456[(1'h0):(1'h0)] ?
                          ((8'ha1) ~^ (reg1469 ?
                              reg1517 : reg1491)) : $signed($unsigned(wire1437))),
                      $unsigned($unsigned(reg1546))} : $unsigned($signed(((~|reg1573) >> $unsigned(reg1445)))));
            end
          else
            begin
              reg1572 <= reg1503;
            end
          for (forvar1577 = (1'h0); (forvar1577 < (2'h2)); forvar1577 = (forvar1577 + (1'h1)))
            begin
              reg1578 <= $unsigned((reg1557[(4'h9):(4'h8)] <<< $signed(reg1575)));
              reg1579 = reg1476[(4'hc):(4'ha)];
              reg1581 <= ($signed((^~(+$unsigned(reg1503)))) ?
                  (($unsigned(reg1492) < (7'h41)) | (^$signed($signed((8'h9c))))) : (($unsigned((reg1561 && reg1445)) ?
                      $signed($signed(reg1578)) : $unsigned($unsigned(reg1472))) * (+reg1554[(5'h11):(4'hb)])));
            end
          reg1582 <= $unsigned((7'h41));
          if ((($unsigned((wire1435 ^~ $unsigned(reg1517))) ?
                  $signed(reg1557) : reg1536) ?
              ((~|((+reg1484) ?
                  reg1577[(3'h4):(2'h3)] : $signed(reg1469))) >>> reg1473) : (reg1502 >>> $signed(($signed((8'had)) ?
                  reg1559 : {reg1559, reg1581, (8'ha2)})))))
            begin
              reg1583 = reg1501[(1'h1):(1'h0)];
              reg1584 <= $unsigned((+((reg1486[(3'h6):(3'h5)] ?
                  (reg1447 && reg1557) : reg1521) >>> (!(!reg1554)))));
              reg1585 <= (7'h58);
              reg1586 = ($unsigned(reg1484) ? (~$unsigned(wire1434)) : reg1584);
            end
          else
            begin
              reg1583 = reg1557;
              reg1584 <= $unsigned($signed(wire1566));
              reg1585 <= ((reg1472 ?
                      (reg1559[(2'h2):(2'h2)] - (reg1470 ?
                          reg1446 : $signed(reg1445))) : (reg1581[(5'h10):(4'ha)] > $unsigned((reg1442 ?
                          (8'haf) : reg1568)))) ?
                  $signed(reg1456[(2'h2):(1'h0)]) : reg1444);
              reg1587 <= $unsigned((({(reg1489 ~^ (8'hbc))} ^~ $signed($unsigned((7'h51)))) ?
                  ({((7'h50) ? reg1495 : (8'hbf)),
                      (~&(7'h44)),
                      $unsigned(wire1436)} & $unsigned((^~(8'ha2)))) : ($signed(wire1436) ^~ $signed((reg1570 ?
                      reg1559 : (8'hb5))))));
              reg1588 = (reg1459[(4'h8):(4'h8)] ?
                  {reg1530,
                      $unsigned(((~|reg1569) < (reg1473 ? reg1564 : reg1545))),
                      (reg1505[(1'h0):(1'h0)] >> reg1496[(4'h8):(3'h5)])} : wire1565);
              reg1589 = $signed(((reg1530[(2'h2):(1'h0)] == $unsigned((reg1477 <<< reg1522))) ?
                  (~^$unsigned(forvar1567[(4'hf):(4'h9)])) : {{reg1486}}));
              reg1590 = ($signed(reg1517) != {$signed($signed($signed(forvar1567))),
                  $unsigned($unsigned({reg1484, reg1530, reg1470})),
                  $unsigned($signed((8'h9c)))});
            end
          if ($signed($signed((|reg1545[(4'hb):(1'h0)]))))
            begin
              reg1591 = $signed(reg1551);
              reg1592 <= {(reg1510[(2'h3):(2'h3)] ?
                      reg1530 : reg1545[(1'h0):(1'h0)])};
              reg1593 <= $unsigned(($signed((^reg1510[(3'h6):(3'h6)])) ?
                  reg1442[(2'h3):(2'h3)] : {$signed({reg1536})}));
              reg1594 <= reg1573;
              reg1595 = ($signed({$unsigned({reg1570}),
                      (&$unsigned(forvar1567))}) ?
                  reg1573 : $unsigned(reg1491));
              reg1596 <= ((reg1476 ?
                  {reg1568[(1'h0):(1'h0)]} : (~(~$unsigned(reg1581)))) || $unsigned(reg1541[(3'h4):(1'h1)]));
            end
          else
            begin
              reg1591 = reg1463;
              reg1595 = reg1444;
              reg1597 = $signed({reg1484[(5'h18):(4'h8)],
                  (~&$unsigned((^reg1596)))});
              reg1598 = (~|$unsigned(reg1559));
              reg1599 <= $unsigned(wire1566[(1'h1):(1'h0)]);
              reg1600 <= {$unsigned((~|reg1541))};
              reg1601 <= reg1554;
            end
        end
      reg1602 <= forvar1567;
      for (forvar1603 = (1'h0); (forvar1603 < (2'h3)); forvar1603 = (forvar1603 + (1'h1)))
        begin
          reg1604 = (~&((reg1583[(1'h0):(1'h0)] ~^ reg1491) + ((~reg1457) ?
              (8'hbd) : ($signed(reg1587) >>> {reg1592, reg1598, wire1434}))));
          reg1605 = (+reg1522);
          for (forvar1606 = (1'h0); (forvar1606 < (2'h3)); forvar1606 = (forvar1606 + (1'h1)))
            begin
              reg1607 = $signed(($signed(reg1492) ~^ forvar1603));
              reg1608 <= {((-reg1595) ?
                      (reg1541 * reg1441[(3'h4):(1'h0)]) : ($signed(reg1597[(3'h5):(3'h4)]) ?
                          reg1452 : {((7'h43) >= wire1566),
                              $signed(reg1546)}))};
            end
          for (forvar1609 = (1'h0); (forvar1609 < (1'h0)); forvar1609 = (forvar1609 + (1'h1)))
            begin
              reg1610 = (+{(!{(reg1607 ? (7'h4b) : reg1486),
                      (~|reg1502),
                      (reg1596 != reg1508)}),
                  ((8'hab) ? reg1546 : $signed($unsigned(reg1583))),
                  (reg1472[(3'h5):(3'h5)] && $unsigned({(8'hae), reg1512}))});
              reg1611 <= (~|($unsigned(((reg1588 ? reg1596 : wire1565) ?
                      reg1452 : $signed(reg1587))) ?
                  wire1438[(5'h11):(5'h10)] : {((reg1548 ? (8'hb2) : reg1580) ?
                          (reg1530 & reg1486) : ((7'h43) ?
                              wire1439 : reg1449))}));
              reg1612 = $unsigned($signed(reg1442[(3'h5):(1'h0)]));
              reg1613 = $signed(reg1608[(2'h2):(1'h1)]);
              reg1614 = (reg1590 ?
                  ($unsigned(reg1505[(2'h3):(1'h0)]) && ((&((7'h4c) ?
                      reg1599 : reg1463)) ~^ ($unsigned(reg1489) >>> (reg1517 << reg1589)))) : (~^($signed(reg1489[(3'h6):(2'h3)]) ?
                      ((reg1569 ? reg1601 : reg1587) ?
                          ((8'hb0) >>> reg1502) : ((7'h58) >= wire1439)) : (reg1476 ?
                          (reg1470 <<< (7'h58)) : $signed(reg1477)))));
              reg1615 = (reg1571[(2'h2):(2'h2)] ?
                  (!((reg1594[(3'h4):(2'h3)] || (reg1592 >>> (8'ha1))) ?
                      reg1611 : $unsigned(reg1455))) : $unsigned(($signed(reg1496[(4'h8):(3'h7)]) <<< ($unsigned(wire1436) + (reg1599 ~^ reg1586)))));
            end
          if (reg1489[(4'hc):(1'h0)])
            begin
              reg1616 = (reg1446[(2'h3):(1'h1)] ?
                  reg1600[(5'h10):(5'h10)] : reg1569);
              reg1617 <= (~^$unsigned({reg1539[(5'h1c):(3'h7)],
                  wire1439,
                  reg1456[(1'h1):(1'h1)]}));
              reg1618 <= ($unsigned(reg1498) << $unsigned(reg1484));
              reg1619 = (-reg1614[(5'h10):(4'h8)]);
            end
          else
            begin
              reg1616 = reg1548;
              reg1619 = ((7'h4f) ?
                  (&$unsigned(reg1588)) : (((8'hb0) || ($unsigned(reg1598) ?
                          reg1455[(3'h4):(2'h2)] : {reg1598, (7'h45)})) ?
                      ($signed((~^(8'h9c))) ?
                          ((8'hbf) << (~|reg1586)) : (+wire1439)) : (^~(((8'hb8) < reg1577) && reg1444[(5'h15):(4'he)]))));
              reg1620 = reg1477[(1'h0):(1'h0)];
              reg1621 <= ({(8'hb4),
                  ((!{forvar1606, reg1568}) ?
                      $unsigned(reg1573[(5'h18):(5'h11)]) : wire1438),
                  reg1573} & (^~$signed(reg1611[(3'h6):(2'h3)])));
              reg1622 = $signed((((~&$unsigned(reg1459)) ?
                      wire1437[(2'h3):(2'h2)] : ($signed(reg1460) ?
                          (wire1436 ? (8'haa) : reg1473) : (reg1616 ?
                              reg1470 : reg1551))) ?
                  (|(reg1559 >> (reg1442 || reg1538))) : ($unsigned(reg1577[(1'h1):(1'h1)]) || (|$unsigned((7'h45))))));
              reg1623 <= $signed((($signed(wire1437[(2'h2):(1'h1)]) == reg1445) ^~ (reg1607 ?
                  {((8'h9d) <<< reg1582),
                      $unsigned((8'hb0))} : (&$unsigned(reg1608)))));
              reg1624 <= $signed((reg1567 >> {reg1569,
                  $unsigned({(8'haa), reg1600, reg1571}),
                  {$signed(reg1442),
                      (reg1598 ? reg1574 : wire1566),
                      ((8'hae) ? reg1499 : reg1614)}}));
            end
          reg1625 <= $unsigned(((reg1460[(4'ha):(3'h5)] << reg1528[(3'h5):(3'h4)]) * $unsigned($unsigned((reg1591 | reg1477)))));
        end
      reg1626 <= reg1449;
      if ((($signed($signed($signed((8'hb5)))) ?
              {reg1580[(2'h2):(2'h2)],
                  reg1444[(4'h9):(2'h2)],
                  reg1489[(4'hb):(2'h3)]} : reg1572[(3'h5):(3'h4)]) ?
          (reg1442[(1'h0):(1'h0)] ^~ reg1575) : $signed((~&((~|reg1585) <<< (~^reg1574))))))
        begin
          for (forvar1627 = (1'h0); (forvar1627 < (3'h6)); forvar1627 = (forvar1627 + (1'h1)))
            begin
              reg1628 <= (($unsigned($unsigned($unsigned(reg1581))) ?
                  reg1442[(2'h3):(2'h3)] : reg1546[(5'h15):(4'h8)]) >>> $signed((|(|$signed((8'hb0))))));
              reg1629 = $signed(wire1439);
              reg1630 <= ($unsigned(reg1505) ? (8'h9f) : $unsigned({(7'h4e)}));
            end
          for (forvar1631 = (1'h0); (forvar1631 < (2'h2)); forvar1631 = (forvar1631 + (1'h1)))
            begin
              reg1632 = reg1528;
              reg1633 <= reg1528;
              reg1634 = ($unsigned((($unsigned((8'had)) ?
                          ((8'hb3) >>> reg1594) : $signed(reg1564)) ?
                      (~^reg1537[(4'h8):(2'h3)]) : reg1586[(3'h4):(1'h0)])) ?
                  (((~|reg1573) << $unsigned((reg1608 ^ reg1604))) ?
                      $signed((|(reg1594 ^~ reg1548))) : ((^~(~^reg1501)) ?
                          ($signed(reg1442) ^ (+reg1496)) : ($signed((8'h9d)) | reg1550[(5'h1a):(5'h10)]))) : wire1435);
              reg1635 = (($signed(reg1571[(2'h3):(1'h1)]) ?
                      (((&reg1564) ?
                              {reg1476, reg1605} : (reg1588 ?
                                  forvar1609 : reg1469)) ?
                          (-$signed(reg1613)) : (~&{reg1473,
                              reg1551})) : reg1472) ?
                  $unsigned(($signed((~|reg1594)) & (&(forvar1567 >>> reg1550)))) : ($unsigned($signed(reg1494)) << reg1624[(5'h17):(2'h2)]));
            end
        end
      else
        begin
          reg1627 = reg1598[(3'h7):(2'h2)];
          for (forvar1628 = (1'h0); (forvar1628 < (2'h2)); forvar1628 = (forvar1628 + (1'h1)))
            begin
              reg1630 <= reg1589[(2'h3):(2'h2)];
              reg1631 = $unsigned($signed($unsigned(reg1626)));
            end
          reg1633 <= $unsigned($signed(((reg1546 < ((8'haf) ?
              reg1554 : (7'h44))) - $unsigned(((8'hb9) ? (8'hbf) : (8'hb1))))));
          reg1636 <= $signed({{((reg1464 ^~ reg1628) ~^ (reg1588 <= reg1598)),
                  ($unsigned((7'h40)) | $unsigned((8'ha0))),
                  reg1618[(4'h8):(2'h3)]},
              $signed(reg1473[(5'h17):(4'he)]),
              (reg1629 ? $unsigned($signed((8'ha5))) : $unsigned((^reg1627)))});
          reg1637 = (reg1447[(4'h8):(1'h0)] ?
              ((^~reg1632) ^~ $signed((8'ha4))) : {(($unsigned(reg1568) + $signed((8'h9f))) ~^ (((8'hba) ?
                          reg1627 : reg1634) ?
                      reg1633 : ((7'h54) - reg1622))),
                  (^~$unsigned($unsigned((8'hb0))))});
          for (forvar1638 = (1'h0); (forvar1638 < (2'h3)); forvar1638 = (forvar1638 + (1'h1)))
            begin
              reg1639 = (8'hae);
            end
          reg1640 = (&(~^reg1486[(3'h4):(2'h2)]));
        end
      for (forvar1641 = (1'h0); (forvar1641 < (3'h4)); forvar1641 = (forvar1641 + (1'h1)))
        begin
          reg1642 <= reg1594;
        end
    end
  always
    @(posedge clk) begin
      for (forvar1643 = (1'h0); (forvar1643 < (3'h6)); forvar1643 = (forvar1643 + (1'h1)))
        begin
          if (reg1568)
            begin
              reg1644 <= (reg1557[(1'h0):(1'h0)] ?
                  reg1554[(5'h19):(5'h16)] : $signed($signed(reg1456[(1'h1):(1'h1)])));
              reg1645 <= (7'h41);
              reg1646 = (~((reg1496 <= (^(7'h49))) ?
                  (^((reg1567 ? reg1494 : wire1437) ?
                      ((8'ha3) >= reg1602) : $unsigned(reg1582))) : reg1539));
              reg1647 <= reg1444[(5'h19):(5'h17)];
              reg1648 = $unsigned($unsigned(($signed($signed(reg1572)) ?
                  reg1576[(4'he):(3'h5)] : ((~|wire1434) ~^ reg1546))));
            end
          else
            begin
              reg1646 = ((~(-reg1601[(2'h2):(1'h1)])) ?
                  reg1592 : $unsigned(((!$signed(reg1546)) == {{reg1494,
                          reg1533}})));
            end
          if ($unsigned(reg1647))
            begin
              reg1649 = (reg1464 >>> reg1569[(3'h6):(1'h0)]);
              reg1650 = (reg1572[(2'h2):(2'h2)] ?
                  (+reg1501) : (reg1450[(4'h9):(3'h6)] || (7'h48)));
              reg1651 <= reg1559;
              reg1652 = reg1530;
            end
          else
            begin
              reg1651 <= $unsigned(reg1572);
              reg1652 = {reg1441, reg1498[(4'h9):(3'h4)], $signed(reg1625)};
              reg1653 = reg1548;
            end
          for (forvar1654 = (1'h0); (forvar1654 < (1'h0)); forvar1654 = (forvar1654 + (1'h1)))
            begin
              reg1655 = $unsigned($unsigned(($signed((reg1626 ?
                  reg1559 : reg1457)) + $unsigned(reg1498[(4'h9):(4'h8)]))));
              reg1656 = reg1592[(3'h7):(2'h2)];
              reg1657 <= $unsigned(({(!(reg1630 - (8'hbb))),
                      reg1633[(1'h1):(1'h0)],
                      $signed(reg1554[(5'h1a):(2'h3)])} ?
                  (+$signed((reg1476 + reg1476))) : (~(reg1510 ?
                      (~^reg1446) : ((7'h46) ? reg1445 : reg1646)))));
              reg1658 <= ((~&reg1528[(3'h6):(2'h3)]) ?
                  (-((~^((8'hbb) ?
                      reg1450 : (8'hb2))) >= wire1435[(4'hf):(4'hf)])) : reg1499[(1'h0):(1'h0)]);
              reg1659 <= $unsigned({(reg1582 ^ (&reg1496)),
                  (-reg1486),
                  {$unsigned((+reg1564))}});
            end
          reg1660 = $unsigned(reg1611);
          reg1661 <= reg1559[(2'h2):(1'h0)];
          reg1662 = {reg1564[(4'hb):(3'h6)],
              (($unsigned($signed(reg1508)) ^ (~^$unsigned(reg1551))) * ($unsigned((7'h55)) ?
                  (|reg1455[(4'hc):(4'h9)]) : reg1492[(5'h11):(4'hd)])),
              ($unsigned(reg1611[(2'h2):(1'h0)]) ^ ($signed((reg1645 ?
                      reg1621 : reg1658)) ?
                  reg1449 : $signed({reg1650})))};
          reg1663 <= ($unsigned($signed((~&$unsigned(reg1537)))) ~^ (&$unsigned(reg1554)));
        end
      for (forvar1664 = (1'h0); (forvar1664 < (1'h1)); forvar1664 = (forvar1664 + (1'h1)))
        begin
          for (forvar1665 = (1'h0); (forvar1665 < (1'h0)); forvar1665 = (forvar1665 + (1'h1)))
            begin
              reg1666 <= reg1656[(4'he):(3'h4)];
              reg1667 <= (reg1494[(1'h1):(1'h1)] ?
                  (reg1489[(4'hd):(4'h9)] == $signed($signed((~^forvar1643)))) : $signed({(&(^reg1624)),
                      reg1494,
                      reg1650[(4'hd):(3'h7)]}));
              reg1668 <= $signed((^~reg1559[(1'h1):(1'h1)]));
            end
          for (forvar1669 = (1'h0); (forvar1669 < (1'h1)); forvar1669 = (forvar1669 + (1'h1)))
            begin
              reg1670 <= reg1624;
              reg1671 = reg1569;
              reg1672 <= ($signed({(((8'ha8) ? (8'ha2) : reg1594) ?
                          (reg1541 ? reg1456 : reg1528) : reg1576)}) ?
                  reg1649[(3'h6):(3'h6)] : $unsigned($signed(reg1447[(4'h8):(2'h3)])));
              reg1673 <= (8'ha7);
              reg1674 <= {(~^(((~|reg1649) ?
                      reg1549[(5'h1b):(5'h19)] : $unsigned(reg1528)) != reg1473[(4'hf):(4'h8)])),
                  ((reg1459 & wire1435) ?
                      (reg1559[(1'h1):(1'h1)] ^~ reg1569) : (((8'hb2) >= (reg1657 ?
                              wire1434 : reg1549)) ?
                          wire1439[(5'h10):(3'h7)] : wire1566)),
                  (~&(^{forvar1643, (reg1456 ? reg1533 : (8'ha4))}))};
              reg1675 <= (8'h9c);
              reg1676 <= reg1626;
            end
          for (forvar1677 = (1'h0); (forvar1677 < (2'h2)); forvar1677 = (forvar1677 + (1'h1)))
            begin
              reg1678 = {wire1566,
                  (~(&((reg1592 ? reg1517 : (7'h4f)) ?
                      ((7'h46) ? reg1582 : reg1587) : $signed(reg1653)))),
                  $signed($signed(reg1447[(3'h5):(3'h5)]))};
              reg1679 = $unsigned((forvar1669 > $unsigned((reg1554[(2'h2):(1'h0)] ?
                  (reg1600 != (7'h4f)) : (reg1646 ? (7'h52) : reg1646)))));
              reg1680 = $signed($unsigned(wire1435));
              reg1681 <= ($unsigned((~^forvar1669)) != reg1444[(3'h5):(1'h1)]);
              reg1682 = (reg1667[(3'h5):(2'h3)] ?
                  (reg1449[(3'h7):(1'h1)] & {(~forvar1669[(4'hd):(4'ha)]),
                      (~^(reg1599 ? (7'h55) : reg1671)),
                      {((7'h45) && reg1530)}}) : $signed((-(^~wire1435[(5'h10):(4'h8)]))));
              reg1683 = (reg1668[(3'h7):(3'h6)] * reg1621);
            end
        end
    end
  assign wire1684 = (reg1675 >= reg1585);
  assign wire1685 = (reg1623 | reg1651);
  module1686 #() modinst1907 (.wire1687(reg1498), .wire1690(reg1502), .wire1689(reg1473), .clk(clk), .wire1688(reg1501), .wire1691(reg1658), .y(wire1906));
  always
    @(posedge clk) begin
      for (forvar1908 = (1'h0); (forvar1908 < (2'h3)); forvar1908 = (forvar1908 + (1'h1)))
        begin
          reg1909 = reg1666;
          if (wire1566[(1'h1):(1'h0)])
            begin
              reg1910 <= $unsigned(reg1503);
              reg1911 <= $unsigned(reg1608);
              reg1912 = $signed((~^$signed(reg1674[(1'h0):(1'h0)])));
              reg1913 = $signed($signed({((~|reg1670) ?
                      $unsigned(reg1681) : $signed(reg1909))}));
              reg1914 = $signed(reg1659);
              reg1915 <= $signed(reg1633);
            end
          else
            begin
              reg1910 <= $unsigned($unsigned(reg1472[(5'h10):(4'hf)]));
              reg1912 = $signed((({$unsigned(reg1647),
                  (~&reg1564),
                  reg1596} << ({reg1668, reg1460, reg1528} ?
                  (reg1486 ?
                      reg1447 : reg1915) : {reg1661})) >= wire1566[(1'h1):(1'h0)]));
              reg1915 <= ($signed(($unsigned((reg1541 * (7'h57))) <= reg1596)) ^ ($unsigned({(reg1447 ?
                          wire1439 : reg1522),
                      $unsigned(forvar1908)}) ?
                  $unsigned(($signed(reg1528) ?
                      $signed(reg1557) : $signed(reg1911))) : reg1456));
              reg1916 <= ((reg1502[(5'h13):(3'h7)] ^ ((~&$unsigned(reg1592)) ?
                      reg1642[(4'hf):(4'hc)] : ((reg1663 >= reg1608) << $signed(forvar1908)))) ?
                  $unsigned((-reg1642[(4'he):(4'h8)])) : ($unsigned(($signed(reg1663) ?
                      $unsigned(reg1602) : reg1676[(4'h9):(1'h1)])) * reg1564));
              reg1917 = $unsigned(($signed(((~|reg1472) * $unsigned(reg1913))) == wire1438[(2'h2):(1'h0)]));
            end
          reg1918 <= reg1470;
          reg1919 <= ($signed({(~&$unsigned((8'ha5))),
              $unsigned((~&reg1548)),
              reg1666}) ^~ $signed(wire1436[(5'h1d):(5'h13)]));
        end
      reg1920 <= $unsigned(reg1621[(4'he):(4'ha)]);
      reg1921 = (8'had);
      reg1922 = reg1916[(1'h0):(1'h0)];
      if (reg1557[(4'ha):(1'h1)])
        begin
          reg1923 = (reg1600[(4'hc):(3'h7)] & $signed((reg1521 <= (reg1491 ?
              (reg1593 ^ reg1557) : reg1672))));
          reg1924 = $signed(reg1594);
          reg1925 <= reg1922;
          if (reg1530)
            begin
              reg1926 = (^(&(reg1548[(3'h4):(1'h0)] ^~ reg1585)));
              reg1927 <= $unsigned(((~^(~|(|wire1436))) ?
                  (|$unsigned($unsigned(reg1545))) : (+(8'hb0))));
              reg1928 <= ((7'h46) ?
                  $unsigned(($signed($unsigned((8'hab))) ?
                      ((^reg1539) << (reg1457 ?
                          reg1626 : (8'hae))) : $signed((reg1599 ?
                          reg1496 : reg1920)))) : (reg1494 ?
                      $signed($unsigned($signed(reg1600))) : (reg1568 ?
                          reg1924[(4'hd):(4'ha)] : (~&(reg1444 || reg1503)))));
            end
          else
            begin
              reg1926 = (~&$signed((reg1501[(1'h1):(1'h1)] ?
                  (reg1927[(3'h6):(1'h1)] & ((8'hbd) ?
                      reg1512 : reg1611)) : ((~^reg1673) ?
                      $signed((8'h9c)) : {reg1484}))));
              reg1929 = {reg1927,
                  ($unsigned((&reg1923)) ?
                      ((~&$signed(reg1494)) ?
                          ({wire1565} ?
                              reg1536 : $signed(reg1549)) : reg1633[(5'h15):(1'h1)]) : (|(&(-reg1572))))};
              reg1930 <= {$unsigned(wire1436),
                  ((8'ha0) ?
                      reg1442 : ({$signed((8'hbc))} ?
                          $signed($unsigned(reg1667)) : (8'ha1)))};
              reg1931 = $signed(reg1657);
            end
          if ($signed($signed(reg1564[(1'h1):(1'h1)])))
            begin
              reg1932 <= (~^($unsigned((~{reg1658,
                  reg1675})) < (reg1494[(1'h1):(1'h1)] ?
                  $unsigned(reg1517[(5'h12):(5'h10)]) : reg1569)));
              reg1933 = $unsigned((reg1441 ~^ $unsigned((((7'h4c) ?
                      wire1685 : (7'h4c)) ?
                  $signed(reg1495) : {(7'h55), reg1484, wire1906}))));
              reg1934 = {$signed(((+$signed((7'h4f))) >= reg1661[(3'h5):(2'h2)]))};
              reg1935 <= $unsigned(reg1549);
              reg1936 <= {{{$signed({(7'h4a), reg1672, wire1436}), reg1578},
                      {(&(reg1446 ? (7'h54) : reg1672)), {{(7'h42), reg1599}}},
                      (&(reg1621 ? {reg1636, reg1674} : $signed(reg1926)))},
                  $unsigned((^~$signed($unsigned((7'h45)))))};
            end
          else
            begin
              reg1933 = {reg1455,
                  (($signed({reg1917}) >= (^reg1521[(1'h0):(1'h0)])) >>> {$unsigned((reg1927 ?
                          reg1473 : reg1582))})};
            end
          for (forvar1937 = (1'h0); (forvar1937 < (3'h5)); forvar1937 = (forvar1937 + (1'h1)))
            begin
              reg1938 <= wire1906[(5'h15):(4'h8)];
              reg1939 = ($unsigned((^reg1925)) ?
                  $signed((+(^reg1636))) : reg1537[(3'h4):(2'h2)]);
            end
          reg1940 <= ($signed($unsigned(($unsigned(wire1684) | (reg1663 == reg1469)))) & $signed($unsigned($unsigned((reg1657 <<< reg1914)))));
        end
      else
        begin
          if ($unsigned(wire1439[(3'h6):(3'h5)]))
            begin
              reg1925 <= reg1919;
              reg1927 <= $signed($signed($signed((reg1934[(1'h0):(1'h0)] ?
                  $unsigned((7'h43)) : (reg1935 && reg1939)))));
              reg1928 <= (!reg1537[(4'h8):(1'h1)]);
            end
          else
            begin
              reg1923 = forvar1908;
              reg1924 = $unsigned(reg1912);
              reg1925 <= (+$signed(((~^(^~reg1449)) && $signed(reg1932[(4'h8):(3'h6)]))));
              reg1926 = $unsigned((reg1576 <<< (7'h48)));
            end
          for (forvar1929 = (1'h0); (forvar1929 < (2'h3)); forvar1929 = (forvar1929 + (1'h1)))
            begin
              reg1931 = reg1549;
              reg1932 <= reg1926;
              reg1935 <= ({((7'h54) && ($signed(reg1624) ?
                          reg1936 : $signed(wire1906)))} ?
                  reg1554[(4'hf):(2'h2)] : reg1538[(2'h3):(2'h2)]);
              reg1937 = (!reg1564);
            end
          if ($signed(reg1668[(1'h1):(1'h1)]))
            begin
              reg1938 <= reg1578[(2'h2):(2'h2)];
              reg1940 <= $unsigned($signed(reg1545));
              reg1941 = {$unsigned(({$signed(reg1621),
                          (reg1625 ? reg1470 : reg1486),
                          ((7'h52) ? reg1549 : reg1594)} ?
                      ($unsigned((8'hbf)) <<< reg1909[(1'h0):(1'h0)]) : ((wire1439 ?
                              reg1572 : reg1593) ?
                          wire1439 : reg1499))),
                  $unsigned($unsigned(((reg1578 - reg1628) == $signed(reg1938))))};
              reg1942 <= $unsigned((~{($signed(reg1910) ?
                      (reg1676 << reg1666) : $unsigned(reg1636)),
                  reg1572,
                  (7'h53)}));
              reg1943 = reg1473;
            end
          else
            begin
              reg1939 = (&reg1472[(4'hf):(1'h0)]);
              reg1940 <= reg1456;
              reg1941 = $unsigned(((8'hbf) ?
                  {$unsigned(reg1913[(4'hf):(3'h7)]),
                      $unsigned(wire1437)} : $unsigned($signed((7'h45)))));
            end
          reg1944 = $unsigned((~reg1548));
          if ($unsigned(reg1593))
            begin
              reg1945 = ($signed($signed($unsigned($signed(reg1675)))) << $signed((^reg1522[(4'hf):(4'hf)])));
              reg1946 = (reg1944[(1'h1):(1'h0)] >> $signed({$unsigned($unsigned(reg1642))}));
              reg1947 = ({$signed(reg1492[(5'h15):(4'h8)]),
                      ((reg1549 != {reg1935, wire1437, (8'ha8)}) ?
                          ((~^reg1572) ?
                              {reg1628} : (reg1539 << (8'ha8))) : wire1565)} ?
                  {$unsigned($signed(reg1533[(4'ha):(3'h5)])),
                      ($unsigned($unsigned((8'ha4))) >= reg1498[(1'h0):(1'h0)]),
                      $unsigned(($signed(reg1581) ?
                          reg1657 : $signed((8'hb7))))} : reg1495[(4'h9):(3'h4)]);
            end
          else
            begin
              reg1948 <= reg1486[(1'h0):(1'h0)];
              reg1949 <= reg1675[(4'he):(4'h8)];
              reg1950 = (~^$unsigned((&(!(~&reg1505)))));
            end
          if ($unsigned({({(reg1651 ? (8'hbe) : (7'h48)),
                      (-(8'h9f)),
                      {reg1926}} ?
                  ((+forvar1929) >> reg1914) : (reg1675 && (reg1929 ?
                      reg1668 : reg1926))),
              $unsigned($unsigned((7'h52))),
              $unsigned($unsigned(reg1594))}))
            begin
              reg1951 <= {reg1557[(3'h4):(2'h3)],
                  $unsigned($unsigned((~reg1663))),
                  $signed(((((8'hbe) ? reg1505 : reg1909) ~^ {reg1510,
                      reg1623}) * (~|{reg1647})))};
              reg1952 <= $unsigned(reg1911);
              reg1953 <= (((^~(~&(7'h54))) ?
                      {$unsigned(((8'hae) <<< reg1922)),
                          $unsigned((8'ha1))} : reg1582) ?
                  (^~((reg1668[(4'hb):(2'h2)] ?
                      $unsigned(reg1935) : {(7'h55)}) << ({reg1572,
                      reg1942,
                      reg1441} & (reg1594 ?
                      reg1498 : reg1645)))) : reg1469[(2'h2):(1'h1)]);
              reg1954 = reg1645[(4'h8):(1'h1)];
            end
          else
            begin
              reg1954 = reg1623;
              reg1955 = $signed(reg1505[(3'h4):(3'h4)]);
              reg1956 = reg1581[(5'h11):(3'h6)];
              reg1957 <= reg1672[(4'ha):(4'h8)];
              reg1958 <= $unsigned((^(($signed(reg1469) >> ((8'hb1) ^ reg1499)) ?
                  reg1625[(4'hd):(4'ha)] : $signed((-reg1492)))));
              reg1959 <= (&reg1642[(4'hd):(4'hc)]);
              reg1960 <= $unsigned(reg1539);
            end
        end
    end
  module1961 #() modinst2322 (wire2321, clk, reg1460, reg1484, reg1495, reg1568, reg1681);
  assign wire2323 = $unsigned($signed(reg1444[(5'h1b):(5'h16)]));
  assign wire2324 = (reg1596 < ((reg1549[(5'h12):(2'h3)] << (((8'h9d) ?
                                reg1630 : reg1441) ?
                            {reg1587,
                                wire1439,
                                reg1464} : reg1463[(3'h4):(2'h3)])) ?
                        ($unsigned($signed(reg1557)) >= {{reg1636,
                                reg1546,
                                (8'hac)},
                            (reg1533 * reg1545)}) : reg1545[(5'h18):(5'h15)]));
  always
    @(posedge clk) begin
      reg2325 <= reg1910[(5'h16):(4'h8)];
    end
  assign wire2326 = $signed(($signed($signed($unsigned((8'hb7)))) ?
                        {$signed($unsigned(wire1566)),
                            ((reg1498 & reg1444) ?
                                (&reg1940) : (reg1617 >>> reg1626)),
                            reg1442} : (^reg1911)));
  always
    @(posedge clk) begin
      if ((-((($unsigned(reg1916) > reg1470) && reg1663[(1'h0):(1'h0)]) | reg1533[(4'hb):(2'h2)])))
        begin
          if (((8'h9d) - (reg1495 ? (^(~^{reg1442, reg1564})) : reg1522)))
            begin
              reg2327 <= (~^$signed({((~&(7'h43)) ?
                      $signed(reg1545) : $signed((8'ha8)))}));
              reg2328 <= (7'h43);
              reg2329 = $signed($unsigned($unsigned(reg1919[(1'h0):(1'h0)])));
              reg2330 <= reg1932;
              reg2331 = reg1636[(2'h2):(2'h2)];
            end
          else
            begin
              reg2329 = $unsigned((^~reg1469));
            end
        end
      else
        begin
          for (forvar2327 = (1'h0); (forvar2327 < (1'h1)); forvar2327 = (forvar2327 + (1'h1)))
            begin
              reg2329 = reg1510;
              reg2331 = $signed($signed(((reg1495[(3'h5):(1'h0)] ?
                      reg1528 : $signed(wire2323)) ?
                  reg1608 : reg1951[(3'h7):(3'h5)])));
              reg2332 = $unsigned(reg1916[(3'h5):(2'h3)]);
              reg2333 = (+reg1915);
            end
          reg2334 = $unsigned((reg1568 ?
              (({reg1920, reg1666} ?
                  (reg1594 ?
                      wire1566 : (8'hb0)) : {(7'h4c)}) != reg1584[(4'he):(4'hd)]) : ($unsigned((reg1578 ?
                  reg1549 : wire1437)) <<< (+$unsigned(reg1538)))));
          for (forvar2335 = (1'h0); (forvar2335 < (2'h3)); forvar2335 = (forvar2335 + (1'h1)))
            begin
              reg2336 = ((~^(reg1545[(3'h5):(3'h4)] ?
                      reg1581[(4'hb):(1'h0)] : ((~^forvar2335) ?
                          {(8'hb0), wire1438, reg2325} : $signed((7'h45))))) ?
                  (^reg1530) : $unsigned($unsigned($signed(reg1559[(1'h1):(1'h0)]))));
              reg2337 <= {(|reg1582),
                  (-{($unsigned((7'h4f)) ? reg1676 : $unsigned(reg1601)),
                      reg1911}),
                  reg2336};
              reg2338 = reg1441[(3'h4):(1'h0)];
              reg2339 = $unsigned(reg1456[(1'h0):(1'h0)]);
              reg2340 <= $unsigned(wire2321);
            end
          reg2341 <= reg1658[(5'h12):(4'hc)];
        end
    end
  always
    @(posedge clk) begin
      reg2342 = (($signed(wire1435[(5'h18):(4'he)]) ?
              ((reg1522[(4'hd):(4'hd)] ?
                      (reg1621 ? (8'h9c) : reg1494) : reg1596) ?
                  $unsigned($signed(reg1536)) : {reg1621,
                      (reg1447 ?
                          reg1505 : reg1441)}) : {($signed(reg1601) ^ reg1460[(4'he):(4'hb)])}) ?
          {(($unsigned(wire2321) << $signed(wire1439)) ?
                  ((7'h4f) ?
                      reg1925[(3'h6):(2'h3)] : reg1473) : (&reg1568[(5'h13):(4'h9)]))} : {$unsigned($signed(reg1444)),
              {($signed(reg1476) ?
                      (reg1512 - reg1567) : {wire1685, wire2324, reg1521})},
              ((!$signed((8'hb9))) ^ ((reg1445 ?
                  (7'h4d) : reg1484) <<< $unsigned(reg1953)))});
      for (forvar2343 = (1'h0); (forvar2343 < (2'h2)); forvar2343 = (forvar2343 + (1'h1)))
        begin
          if ((~|{$signed($signed(reg1594[(3'h4):(1'h0)]))}))
            begin
              reg2344 = ($signed(($unsigned($unsigned(reg1548)) || $unsigned((-(8'h9d))))) || reg1489[(4'he):(1'h1)]);
              reg2345 <= reg1522[(2'h3):(1'h1)];
              reg2346 = reg1949[(5'h11):(2'h3)];
              reg2347 = ($signed($signed((-(|reg1602)))) ?
                  $signed((~^(&{reg1633, reg1442, reg1464}))) : (|(~|reg2325)));
            end
          else
            begin
              reg2345 <= reg1600[(5'h12):(3'h4)];
              reg2346 = {$unsigned(((((8'hb0) ? reg1446 : reg1536) ?
                      wire2324[(5'h17):(5'h11)] : (8'hac)) << (forvar2343 & wire1436[(3'h5):(3'h4)]))),
                  (+(~wire1906[(4'he):(3'h5)])),
                  $signed((|((reg1486 ^~ (8'ha0)) ?
                      (reg1960 < reg1919) : wire1436)))};
              reg2347 = $signed($unsigned((reg1663 ?
                  $unsigned($signed(reg1608)) : ((reg1596 & reg1508) * (wire2326 != reg1587)))));
            end
        end
      reg2348 <= {((^~reg1594) ?
              $signed((-reg1510[(4'h8):(3'h5)])) : $unsigned($unsigned((~&reg2345)))),
          wire2324};
      reg2349 <= $signed(($signed({$signed(reg1576)}) | (reg1948 > reg1602)));
      for (forvar2350 = (1'h0); (forvar2350 < (1'h0)); forvar2350 = (forvar2350 + (1'h1)))
        begin
          if ($unsigned({$signed(wire1439[(1'h1):(1'h1)])}))
            begin
              reg2351 <= (~^reg1659);
              reg2352 = wire1565[(5'h17):(3'h4)];
              reg2353 = $signed(reg1550);
              reg2354 = reg1463[(2'h3):(2'h3)];
            end
          else
            begin
              reg2351 <= ((-(wire2324 ?
                  ({reg1469} ?
                      ((8'hbb) ?
                          reg1473 : reg1674) : $signed(wire1438)) : ($unsigned(reg1681) >>> (reg1463 << forvar2350)))) | reg1621);
              reg2352 = reg1938[(4'he):(3'h4)];
              reg2355 <= $unsigned({$unsigned((^{reg1460}))});
              reg2356 = $unsigned($signed(reg1617[(1'h0):(1'h0)]));
              reg2357 <= $signed((-reg1441[(2'h3):(1'h1)]));
              reg2358 = reg1476[(2'h2):(1'h1)];
              reg2359 = reg1463;
            end
          reg2360 = reg2327;
          reg2361 <= reg1469;
          if ((^(~|((reg1447 < (reg1676 > reg1561)) ?
              $unsigned((reg1510 ?
                  reg1647 : reg2330)) : reg1936[(2'h2):(1'h0)]))))
            begin
              reg2362 = $unsigned((&(reg1486[(4'h8):(4'h8)] ?
                  ((reg1960 ? (7'h46) : wire1437) ?
                      $unsigned(reg1561) : (^reg1476)) : $signed($signed(reg1561)))));
            end
          else
            begin
              reg2363 <= reg1647;
              reg2364 = $unsigned(((reg1636 ?
                  (~|(reg1495 ^ (8'hbb))) : reg1492) > reg1486[(1'h1):(1'h0)]));
              reg2365 <= $unsigned((reg2330 ?
                  (|$signed((~&reg1502))) : (~&reg1486)));
              reg2366 = {reg1633[(4'he):(3'h4)]};
            end
          reg2367 = ($signed($unsigned($unsigned({(7'h43)}))) ?
              {$signed((~|$unsigned(reg1667))),
                  wire1565[(4'h9):(3'h6)]} : $signed((^~($signed(wire2323) >= $signed(reg1930)))));
          reg2368 = reg2346;
          reg2369 = {(reg1533 | reg1626[(4'he):(3'h7)]),
              (($unsigned((reg1444 ? reg1476 : reg1551)) ?
                      reg1455[(4'he):(4'ha)] : ($signed(reg1952) < reg1536)) ?
                  $unsigned($unsigned(reg1596)) : {(^$signed(reg1651)),
                      reg1663}),
              $unsigned(reg2340)};
        end
      reg2370 = $signed($signed(((&$unsigned(reg1644)) > {{reg1623, reg1596},
          (~wire2324)})));
      reg2371 <= (((8'ha4) ^ (reg2325[(4'hb):(4'h8)] >= {{reg2347,
                  reg1911,
                  reg1668},
              $unsigned(reg1444),
              (reg2369 ? reg2352 : (8'ha0))})) ?
          $unsigned((~|$unsigned((reg1675 ?
              (7'h45) : reg1584)))) : $unsigned(({(!(7'h4e))} ?
              ({(8'h9d),
                  reg2364,
                  reg1935} ~^ (reg1561 | reg2328)) : {(^reg1521),
                  reg1578[(2'h2):(1'h0)]})));
    end
  always
    @(posedge clk) begin
      if (reg1953)
        begin
          reg2372 = (-(reg1601 != {$signed((~|(8'ha3))),
              {(8'ha1), reg1644[(4'h8):(4'h8)]},
              reg1473[(1'h1):(1'h1)]}));
          reg2373 = (({(&reg1910[(5'h11):(1'h1)]),
                  wire1437[(1'h0):(1'h0)]} >= $unsigned(($signed((8'ha0)) != (reg1576 ?
                  reg1572 : wire1566)))) ?
              (reg1444 | ((~|reg1508[(3'h7):(1'h1)]) ?
                  reg1477[(2'h3):(2'h3)] : reg1960[(5'h13):(4'h9)])) : (reg1958[(4'he):(1'h1)] ?
                  (&reg1472[(2'h2):(1'h0)]) : {(+(^reg1930)),
                      (((8'hb2) != reg1925) != $signed((8'haf))),
                      ((8'hb8) << (-(7'h54)))}));
          reg2374 <= reg1642;
        end
      else
        begin
          if (((^~(reg1942 ? {(reg1601 ? reg1630 : (7'h47))} : reg1932)) ?
              $unsigned($unsigned($signed((reg1452 ?
                  reg1587 : reg1587)))) : reg1936))
            begin
              reg2372 = ($unsigned({$unsigned((~|reg2327))}) ?
                  {$signed((reg1600[(5'h15):(4'ha)] <<< $unsigned(reg1661))),
                      $unsigned((^~(-wire1436))),
                      (-$signed({reg1675,
                          wire1436}))} : reg1957[(4'h8):(3'h7)]);
            end
          else
            begin
              reg2372 = $unsigned(($signed(({reg1601} ?
                      (reg1647 ? reg1505 : reg1541) : reg1587[(3'h5):(1'h0)])) ?
                  reg1567 : wire2324));
              reg2374 <= reg1494[(2'h2):(2'h2)];
            end
          reg2375 <= $unsigned((~|(&reg1512)));
          reg2376 = (^$unsigned($unsigned((~reg1958[(4'h8):(4'h8)]))));
          reg2377 = reg1587;
          for (forvar2378 = (1'h0); (forvar2378 < (1'h0)); forvar2378 = (forvar2378 + (1'h1)))
            begin
              reg2379 = $signed(($signed(reg1958) ?
                  ($signed(wire2321) > ((-reg1587) > (reg1502 ?
                      reg1469 : reg1545))) : $signed(reg1935)));
              reg2380 = ((reg1930 ?
                  $signed({(reg1645 == reg2337)}) : $unsigned({(wire1438 ?
                          reg1667 : reg2377),
                      (reg1651 > reg1959),
                      (reg2375 ?
                          (7'h43) : reg1600)})) >>> $unsigned(reg2327[(1'h0):(1'h0)]));
              reg2381 = $unsigned(($unsigned((~{reg1508, reg2371, reg2376})) ?
                  $signed({(^~reg1592)}) : reg1911[(1'h1):(1'h1)]));
              reg2382 <= (~|reg1611);
              reg2383 = $unsigned(reg1551);
            end
        end
      reg2384 <= {reg2371};
      if (($unsigned($signed(reg1911)) ?
          reg1460[(4'h9):(3'h7)] : $unsigned((|{reg1559,
              {reg1495, reg1911},
              {reg1657, reg1608, reg2381}}))))
        begin
          reg2385 <= forvar2378;
          reg2386 = $signed(({((^~reg2348) >> (reg1659 ? (8'hb8) : (8'hb8))),
              $unsigned($signed(reg1681))} << ((7'h4c) ?
              reg2384 : reg1625[(3'h5):(3'h5)])));
          if (reg1546)
            begin
              reg2387 = reg1582[(5'h16):(2'h2)];
              reg2388 <= reg1676[(3'h5):(1'h1)];
              reg2389 <= (((reg1618[(4'h9):(3'h7)] - reg1623[(3'h4):(2'h2)]) ?
                  reg1559 : (~|wire1438)) == reg1617[(3'h4):(1'h1)]);
              reg2390 = reg1621[(1'h0):(1'h0)];
            end
          else
            begin
              reg2387 = (|{(^~$signed(reg1960[(5'h19):(1'h1)])),
                  (+{(reg1470 >>> reg1938)})});
              reg2390 = $signed(reg1569[(3'h6):(3'h4)]);
              reg2391 <= ((reg1576 ?
                      reg1495 : (reg1910 ?
                          $signed((reg1644 ?
                              reg1578 : reg1541)) : reg1508[(4'hf):(4'hd)])) ?
                  {($signed($unsigned((8'ha6))) ?
                          reg2389[(3'h5):(2'h3)] : $signed((wire1685 != reg1548)))} : ($signed($unsigned(reg2372[(1'h1):(1'h0)])) || reg1958));
              reg2392 = $unsigned({{$signed((8'ha2)),
                      $unsigned(reg1958[(4'h9):(3'h5)]),
                      reg2351[(1'h1):(1'h0)]}});
              reg2393 = (wire1437 ^~ (reg2390 || reg1626[(1'h1):(1'h0)]));
              reg2394 = reg1668[(2'h2):(1'h0)];
            end
        end
      else
        begin
          reg2385 <= reg1608;
          if ($unsigned($unsigned(reg1569[(4'h8):(3'h5)])))
            begin
              reg2386 = (|$unsigned((+({reg1911, (8'ha5)} | (reg1472 ?
                  reg2380 : wire1437)))));
              reg2388 <= (((8'h9f) > $signed(((reg1486 << (7'h51)) ?
                  reg1537 : (~&wire1438)))) ~^ $signed(($signed(((8'hb6) <= reg1499)) ?
                  $unsigned($unsigned(reg1545)) : ($signed(reg1581) == (reg1948 << reg1625)))));
              reg2389 <= $unsigned((wire1438[(4'hc):(4'ha)] ?
                  ($unsigned((reg1561 & reg2380)) <= {$signed((7'h40))}) : wire1565));
            end
          else
            begin
              reg2386 = $signed((7'h4f));
              reg2388 <= {{(reg1491[(3'h6):(3'h4)] ~^ (reg1441 <<< $signed(wire1685))),
                      (($signed(reg1658) | (~|reg1492)) ?
                          {$signed(reg1508),
                              {reg1621},
                              reg2341[(4'h8):(1'h1)]} : $unsigned($unsigned(wire2323)))}};
              reg2389 <= {{$unsigned(reg1601[(2'h2):(2'h2)])},
                  (((~(-reg1456)) ?
                      $unsigned({(7'h48),
                          (8'ha2),
                          reg1495}) : $signed((reg1486 ?
                          (7'h4b) : (8'hbc)))) - $unsigned($unsigned($unsigned(reg1476))))};
              reg2390 = $signed((~|(|$signed(reg1676))));
              reg2392 = reg1676;
            end
          if (($unsigned($unsigned(($unsigned(reg1675) ?
              (reg1495 ? reg1449 : (8'ha6)) : $unsigned(reg2325)))) << reg2345))
            begin
              reg2393 = reg1594[(1'h0):(1'h0)];
              reg2395 <= (reg1567[(4'hb):(1'h1)] ?
                  $signed((~^reg1476)) : (((8'hbf) && ((^wire2323) > reg1958[(5'h10):(4'he)])) ?
                      $unsigned((~&$unsigned(reg1449))) : reg1667));
              reg2396 <= reg1676[(3'h7):(1'h0)];
              reg2397 <= {(reg1949 ?
                      reg1469[(2'h2):(1'h0)] : ($unsigned(reg1910[(4'he):(3'h4)]) ?
                          reg1572[(4'h9):(3'h4)] : $signed($unsigned(reg1444)))),
                  reg1599,
                  (!reg1919[(1'h0):(1'h0)])};
              reg2398 = $unsigned(($signed(reg2375) ?
                  (reg1486 ^ reg1663) : reg1608[(1'h0):(1'h0)]));
              reg2399 <= {reg2340};
              reg2400 = (reg1512 == (($signed((|reg2373)) ?
                      (8'hb0) : ((reg1645 ?
                          (8'h9c) : reg2363) >> reg1911[(1'h1):(1'h1)])) ?
                  reg1557[(3'h4):(3'h4)] : reg2361[(4'h9):(2'h2)]));
            end
          else
            begin
              reg2393 = $signed(($unsigned(($unsigned(reg1494) ~^ ((8'hab) ?
                  reg1600 : (7'h47)))) | (-($unsigned(reg1582) ?
                  reg1503 : ((8'ha0) >> reg1559)))));
              reg2394 = ((&($unsigned((reg1477 ? reg1919 : (7'h50))) ?
                      reg1936[(4'hd):(4'h8)] : (~&$signed(reg2381)))) ?
                  {(((reg2372 != wire2326) ?
                              $unsigned(reg1592) : reg1958[(2'h2):(1'h0)]) ?
                          $unsigned((~reg1927)) : (wire2326[(3'h5):(2'h2)] + reg1602)),
                      $unsigned($unsigned(reg2376[(3'h7):(3'h7)]))} : reg2389);
              reg2398 = reg1569[(3'h5):(2'h3)];
              reg2400 = reg1624;
            end
          for (forvar2401 = (1'h0); (forvar2401 < (2'h2)); forvar2401 = (forvar2401 + (1'h1)))
            begin
              reg2402 <= $signed(({($unsigned(reg1952) < (reg2392 ?
                          (8'ha5) : wire1685))} ?
                  reg1470[(3'h7):(3'h6)] : $unsigned($unsigned((reg1593 ?
                      (7'h58) : reg1541)))));
              reg2403 <= $unsigned(((8'ha6) ?
                  (~^$signed((reg1584 ?
                      reg2325 : reg1492))) : (~|{reg2385[(4'hd):(4'ha)],
                      (reg2389 ^ reg1601),
                      $unsigned(reg1940)})));
              reg2404 = reg1666[(4'hc):(4'h9)];
              reg2405 = (((({reg1672, reg2388} >> {reg1503,
                          reg1484}) - (&wire2324)) ?
                      $unsigned((^~$signed(reg1668))) : $unsigned($unsigned((wire1906 ?
                          reg1549 : (7'h50))))) ?
                  {((&$unsigned(reg1958)) ^ $unsigned((!(8'hb6)))),
                      {(reg2365[(4'h8):(2'h3)] ?
                              reg2384[(1'h0):(1'h0)] : reg1958),
                          reg1567},
                      reg1464[(3'h5):(2'h3)]} : ($signed(reg1663) << wire1438[(4'ha):(2'h3)]));
            end
          for (forvar2406 = (1'h0); (forvar2406 < (3'h6)); forvar2406 = (forvar2406 + (1'h1)))
            begin
              reg2407 <= reg1935[(1'h0):(1'h0)];
              reg2408 <= reg1587;
              reg2409 = reg1528[(5'h13):(2'h3)];
              reg2410 = $unsigned($signed(((reg1958[(5'h1c):(5'h14)] ?
                  $signed(wire2326) : (7'h47)) & ({wire2326,
                  (7'h56)} <<< ((7'h43) ? reg1517 : reg1935)))));
              reg2411 = reg1935[(3'h7):(3'h5)];
              reg2412 <= (reg2348 && {$signed(reg1486[(3'h4):(3'h4)])});
              reg2413 <= reg1512[(1'h0):(1'h0)];
            end
          for (forvar2414 = (1'h0); (forvar2414 < (2'h2)); forvar2414 = (forvar2414 + (1'h1)))
            begin
              reg2415 = $unsigned(({{$unsigned(reg2384),
                      reg1617[(1'h1):(1'h1)],
                      reg2392[(4'hb):(2'h2)]},
                  $unsigned((^reg1675)),
                  (~^$signed(reg1477))} < (8'hbb)));
              reg2416 <= (~reg1633);
              reg2417 <= $signed(reg1675[(4'hb):(3'h6)]);
              reg2418 <= ($signed(($signed(reg2377[(4'hb):(4'h8)]) ?
                  $unsigned((+wire1439)) : forvar2378[(1'h1):(1'h0)])) < ((~(reg2395[(1'h0):(1'h0)] >>> (reg2412 ?
                      forvar2406 : reg1447))) ?
                  ((~&reg1919) ?
                      $unsigned($signed(reg1930)) : (-reg1910[(1'h0):(1'h0)])) : reg2380));
            end
          if (($unsigned((reg1645 ?
              reg1668[(4'h9):(4'h8)] : wire1906[(5'h16):(5'h16)])) | reg2373[(1'h0):(1'h0)]))
            begin
              reg2419 = {(^reg1596[(3'h4):(1'h1)]),
                  ($unsigned(reg1623) | {({reg1469,
                          reg1936} | ((8'ha9) >> forvar2378)),
                      ((reg1578 ? reg2383 : reg2330) ?
                          reg1499 : reg2385[(4'hc):(3'h4)])}),
                  ((!((~|reg2409) <<< reg1538)) >= $unsigned((|{wire1685,
                      reg2383})))};
              reg2420 = {(|((^~(|wire1906)) - (reg1617[(2'h2):(1'h1)] ?
                      $unsigned(reg1928) : $signed(reg2394)))),
                  $signed($signed(((reg1528 * reg1446) ^ $unsigned(reg1447)))),
                  (($signed($unsigned(reg1510)) ?
                      $unsigned(wire1439) : wire2323[(2'h2):(2'h2)]) >> reg1623[(5'h11):(4'hc)])};
            end
          else
            begin
              reg2421 <= {reg1633, reg2373};
              reg2422 <= ({$signed(reg1495),
                      (reg1596[(4'hc):(3'h5)] << $signed(reg1621))} ?
                  $unsigned(reg1915[(4'hc):(4'hc)]) : reg1486);
            end
        end
      reg2423 <= wire2324[(4'he):(2'h2)];
      for (forvar2424 = (1'h0); (forvar2424 < (1'h1)); forvar2424 = (forvar2424 + (1'h1)))
        begin
          reg2425 = (reg1936 & (reg2410[(2'h3):(1'h0)] ?
              (reg1633 ?
                  ($unsigned(reg1602) ?
                      reg1659 : {reg1668,
                          reg1549,
                          (7'h43)}) : $signed(reg1559)) : (+$unsigned($unsigned((7'h43))))));
          for (forvar2426 = (1'h0); (forvar2426 < (1'h0)); forvar2426 = (forvar2426 + (1'h1)))
            begin
              reg2427 <= (wire1685[(4'hc):(3'h7)] + $signed((reg2337 ?
                  reg2349[(4'he):(3'h5)] : $signed(reg1633))));
              reg2428 = $unsigned({reg1449[(4'ha):(3'h7)], reg1450});
              reg2429 = $unsigned({$signed(reg1659[(5'h1c):(1'h1)])});
              reg2430 = ((reg2413 || $unsigned((^~reg1942[(5'h13):(4'ha)]))) | (-$unsigned($unsigned(reg1498))));
              reg2431 <= $signed(($signed({reg2417[(5'h15):(5'h15)],
                  $signed(reg1457)}) == $signed($unsigned($signed((7'h42))))));
              reg2432 <= (+wire2321);
              reg2433 = reg2377[(4'hc):(2'h2)];
            end
          reg2434 = reg2428[(5'h16):(3'h6)];
          reg2435 = $signed(($unsigned(((reg1608 > (7'h54)) >= (reg1441 << (7'h4e)))) <<< $signed($unsigned((reg1554 ?
              reg1460 : reg1953)))));
        end
    end
  assign wire2436 = reg1916[(3'h7):(1'h0)];
  assign wire2437 = (reg1569 ?
                        $unsigned($signed($unsigned(reg1551))) : ((reg1642 ?
                            $signed((reg1611 ?
                                reg1916 : reg1502)) : (-$signed(reg2337))) != (((wire1435 ?
                                (8'h9d) : reg2355) ?
                            (reg2427 ?
                                reg2412 : reg1585) : $signed(reg2427)) >> (reg1647 ?
                            (reg1568 << reg1675) : reg2395))));
  assign wire2438 = ({($unsigned($unsigned(reg1633)) < ({reg2361, reg1501} ?
                            (|reg1618) : reg1505)),
                        wire1684[(5'h10):(5'h10)]} >> (8'hbe));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module52  (y, clk, wire57, wire56, wire55, wire54, wire53);
  output wire [(32'hfa0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire57;
  input wire [(4'he):(1'h0)] wire56;
  input wire [(5'h18):(1'h0)] wire55;
  input wire [(5'h13):(1'h0)] wire54;
  input wire signed [(3'h7):(1'h0)] wire53;
  wire [(3'h6):(1'h0)] wire1272;
  wire signed [(3'h5):(1'h0)] wire1271;
  wire signed [(5'h10):(1'h0)] wire1269;
  wire [(5'h13):(1'h0)] wire350;
  wire signed [(5'h11):(1'h0)] wire349;
  wire signed [(4'hf):(1'h0)] wire348;
  wire signed [(5'h1b):(1'h0)] wire313;
  wire [(5'h16):(1'h0)] wire157;
  wire signed [(4'hb):(1'h0)] wire156;
  wire [(4'hd):(1'h0)] wire155;
  wire [(5'h10):(1'h0)] wire154;
  wire [(5'h13):(1'h0)] wire87;
  wire signed [(4'hf):(1'h0)] wire58;
  reg [(5'h14):(1'h0)] reg422 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg421 = (1'h0);
  reg [(5'h1d):(1'h0)] reg419 = (1'h0);
  reg [(3'h5):(1'h0)] reg417 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg415 = (1'h0);
  reg [(3'h7):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg410 = (1'h0);
  reg [(3'h5):(1'h0)] reg409 = (1'h0);
  reg [(2'h2):(1'h0)] reg408 = (1'h0);
  reg [(5'h1c):(1'h0)] reg406 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg402 = (1'h0);
  reg [(5'h16):(1'h0)] reg401 = (1'h0);
  reg [(5'h1a):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg398 = (1'h0);
  reg [(5'h11):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg390 = (1'h0);
  reg [(3'h6):(1'h0)] reg389 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg387 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg385 = (1'h0);
  reg [(5'h1e):(1'h0)] reg384 = (1'h0);
  reg [(4'hb):(1'h0)] reg383 = (1'h0);
  reg [(4'hd):(1'h0)] reg379 = (1'h0);
  reg [(5'h1a):(1'h0)] reg378 = (1'h0);
  reg [(5'h1e):(1'h0)] reg373 = (1'h0);
  reg [(5'h14):(1'h0)] reg372 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg370 = (1'h0);
  reg [(2'h3):(1'h0)] reg368 = (1'h0);
  reg [(4'hd):(1'h0)] reg367 = (1'h0);
  reg [(5'h1b):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg363 = (1'h0);
  reg [(4'hf):(1'h0)] reg357 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg355 = (1'h0);
  reg [(5'h1c):(1'h0)] reg347 = (1'h0);
  reg [(4'hc):(1'h0)] reg346 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg345 = (1'h0);
  reg [(5'h16):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg338 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg337 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg326 = (1'h0);
  reg [(4'he):(1'h0)] reg325 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg178 = (1'h0);
  reg [(4'he):(1'h0)] reg177 = (1'h0);
  reg [(5'h1f):(1'h0)] reg175 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg174 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg167 = (1'h0);
  reg [(2'h2):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg160 = (1'h0);
  reg [(3'h4):(1'h0)] reg159 = (1'h0);
  reg [(5'h1f):(1'h0)] reg148 = (1'h0);
  reg [(3'h5):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg146 = (1'h0);
  reg [(5'h1d):(1'h0)] reg143 = (1'h0);
  reg [(5'h1b):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg136 = (1'h0);
  reg [(5'h16):(1'h0)] reg134 = (1'h0);
  reg [(5'h18):(1'h0)] reg132 = (1'h0);
  reg [(5'h12):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg124 = (1'h0);
  reg signed [(4'he):(1'h0)] reg123 = (1'h0);
  reg [(5'h1d):(1'h0)] reg121 = (1'h0);
  reg [(5'h15):(1'h0)] reg119 = (1'h0);
  reg [(5'h1a):(1'h0)] reg118 = (1'h0);
  reg [(5'h14):(1'h0)] reg116 = (1'h0);
  reg [(5'h1d):(1'h0)] reg115 = (1'h0);
  reg [(3'h7):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg112 = (1'h0);
  reg [(5'h1b):(1'h0)] reg111 = (1'h0);
  reg [(3'h7):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg103 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg101 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg98 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg97 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg93 = (1'h0);
  reg [(5'h18):(1'h0)] reg92 = (1'h0);
  reg [(4'ha):(1'h0)] reg91 = (1'h0);
  reg [(3'h4):(1'h0)] reg90 = (1'h0);
  reg [(5'h15):(1'h0)] reg85 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg78 = (1'h0);
  reg [(5'h1a):(1'h0)] reg73 = (1'h0);
  reg [(5'h1f):(1'h0)] reg72 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg65 = (1'h0);
  reg [(2'h2):(1'h0)] reg63 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg60 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg423 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg420 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg418 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg416 = (1'h0);
  reg [(2'h2):(1'h0)] reg413 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg412 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg411 = (1'h0);
  reg [(5'h1e):(1'h0)] reg407 = (1'h0);
  reg [(5'h13):(1'h0)] reg404 = (1'h0);
  reg signed [(4'he):(1'h0)] reg400 = (1'h0);
  reg [(5'h18):(1'h0)] reg397 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar396 = (1'h0);
  reg [(5'h1e):(1'h0)] reg394 = (1'h0);
  reg [(3'h4):(1'h0)] reg393 = (1'h0);
  reg [(2'h2):(1'h0)] reg392 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg391 = (1'h0);
  reg [(4'ha):(1'h0)] reg386 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg382 = (1'h0);
  reg [(3'h4):(1'h0)] reg381 = (1'h0);
  reg [(5'h1f):(1'h0)] reg380 = (1'h0);
  reg [(5'h1a):(1'h0)] reg377 = (1'h0);
  reg [(4'hf):(1'h0)] reg376 = (1'h0);
  reg [(5'h13):(1'h0)] reg375 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg371 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg369 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg365 = (1'h0);
  reg [(5'h12):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg362 = (1'h0);
  reg [(5'h15):(1'h0)] reg361 = (1'h0);
  reg [(5'h12):(1'h0)] reg360 = (1'h0);
  reg [(5'h1f):(1'h0)] reg359 = (1'h0);
  reg [(5'h1e):(1'h0)] reg358 = (1'h0);
  reg [(4'h8):(1'h0)] forvar356 = (1'h0);
  reg [(4'he):(1'h0)] reg354 = (1'h0);
  reg [(5'h13):(1'h0)] forvar353 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar352 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg351 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg341 = (1'h0);
  reg [(5'h18):(1'h0)] forvar340 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg339 = (1'h0);
  reg [(5'h1f):(1'h0)] reg336 = (1'h0);
  reg [(3'h4):(1'h0)] forvar335 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg333 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg332 = (1'h0);
  reg [(3'h4):(1'h0)] reg329 = (1'h0);
  reg [(5'h1c):(1'h0)] reg328 = (1'h0);
  reg [(5'h1c):(1'h0)] reg324 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg323 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg321 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg320 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar319 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg317 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar316 = (1'h0);
  reg [(3'h7):(1'h0)] reg315 = (1'h0);
  reg [(5'h18):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar171 = (1'h0);
  reg [(3'h4):(1'h0)] reg170 = (1'h0);
  reg [(5'h1a):(1'h0)] reg169 = (1'h0);
  reg [(2'h3):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg165 = (1'h0);
  reg [(4'ha):(1'h0)] reg164 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg163 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg162 = (1'h0);
  reg [(4'he):(1'h0)] forvar161 = (1'h0);
  reg [(3'h7):(1'h0)] reg158 = (1'h0);
  reg signed [(4'he):(1'h0)] reg153 = (1'h0);
  reg [(3'h6):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg151 = (1'h0);
  reg [(5'h1f):(1'h0)] reg150 = (1'h0);
  reg [(3'h7):(1'h0)] reg149 = (1'h0);
  reg [(5'h13):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar144 = (1'h0);
  reg [(3'h5):(1'h0)] reg141 = (1'h0);
  reg [(4'hf):(1'h0)] reg140 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg137 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg135 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar130 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar129 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg127 = (1'h0);
  reg [(3'h7):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg122 = (1'h0);
  reg [(5'h15):(1'h0)] forvar120 = (1'h0);
  reg [(5'h18):(1'h0)] forvar105 = (1'h0);
  reg [(4'he):(1'h0)] reg117 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg114 = (1'h0);
  reg [(3'h7):(1'h0)] reg109 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg107 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg106 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg102 = (1'h0);
  reg [(4'h9):(1'h0)] reg96 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar93 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg89 = (1'h0);
  reg [(3'h7):(1'h0)] forvar88 = (1'h0);
  reg [(4'ha):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar82 = (1'h0);
  reg [(5'h15):(1'h0)] reg81 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg79 = (1'h0);
  reg [(5'h1d):(1'h0)] reg77 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg76 = (1'h0);
  reg [(5'h1a):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg71 = (1'h0);
  reg [(5'h1d):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg69 = (1'h0);
  reg [(4'hf):(1'h0)] reg68 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg67 = (1'h0);
  reg [(5'h1f):(1'h0)] reg64 = (1'h0);
  reg [(5'h12):(1'h0)] reg62 = (1'h0);
  reg [(3'h4):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar59 = (1'h0);
  assign y = {wire1272,
                 wire1271,
                 wire1269,
                 wire350,
                 wire349,
                 wire348,
                 wire313,
                 wire157,
                 wire156,
                 wire155,
                 wire154,
                 wire87,
                 wire58,
                 reg422,
                 reg421,
                 reg419,
                 reg417,
                 reg415,
                 reg414,
                 reg410,
                 reg409,
                 reg408,
                 reg406,
                 reg405,
                 reg403,
                 reg402,
                 reg401,
                 reg399,
                 reg398,
                 reg395,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg385,
                 reg384,
                 reg383,
                 reg379,
                 reg378,
                 reg373,
                 reg372,
                 reg370,
                 reg368,
                 reg367,
                 reg366,
                 reg363,
                 reg357,
                 reg355,
                 reg347,
                 reg346,
                 reg345,
                 reg342,
                 reg338,
                 reg337,
                 reg331,
                 reg330,
                 reg327,
                 reg326,
                 reg325,
                 reg322,
                 reg178,
                 reg177,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg167,
                 reg166,
                 reg160,
                 reg159,
                 reg148,
                 reg147,
                 reg146,
                 reg143,
                 reg142,
                 reg138,
                 reg136,
                 reg134,
                 reg132,
                 reg131,
                 reg126,
                 reg124,
                 reg123,
                 reg121,
                 reg119,
                 reg118,
                 reg116,
                 reg115,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg105,
                 reg104,
                 reg103,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg85,
                 reg84,
                 reg83,
                 reg78,
                 reg73,
                 reg72,
                 reg66,
                 reg65,
                 reg63,
                 reg60,
                 reg423,
                 reg420,
                 reg418,
                 reg416,
                 reg413,
                 reg412,
                 reg411,
                 reg407,
                 reg404,
                 reg400,
                 reg397,
                 forvar396,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg386,
                 reg382,
                 reg381,
                 reg380,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg371,
                 reg369,
                 reg365,
                 reg364,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 forvar356,
                 reg354,
                 forvar353,
                 forvar352,
                 reg351,
                 reg344,
                 reg343,
                 reg341,
                 forvar340,
                 reg339,
                 reg336,
                 forvar335,
                 reg334,
                 reg333,
                 reg332,
                 reg329,
                 reg328,
                 reg324,
                 reg323,
                 reg321,
                 reg320,
                 forvar319,
                 reg318,
                 reg317,
                 forvar316,
                 reg315,
                 reg176,
                 forvar171,
                 reg170,
                 reg169,
                 reg168,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 forvar161,
                 reg158,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg145,
                 forvar144,
                 reg141,
                 reg140,
                 reg139,
                 reg137,
                 reg135,
                 reg133,
                 forvar130,
                 forvar129,
                 reg128,
                 reg127,
                 reg125,
                 reg122,
                 forvar120,
                 forvar105,
                 reg117,
                 reg114,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg102,
                 reg96,
                 reg95,
                 forvar93,
                 reg89,
                 forvar88,
                 reg86,
                 forvar82,
                 reg81,
                 reg80,
                 reg79,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg64,
                 reg62,
                 reg61,
                 forvar59,
                 (1'h0)};
  assign wire58 = $signed((wire53 ^ $unsigned(wire53)));
  always
    @(posedge clk) begin
      for (forvar59 = (1'h0); (forvar59 < (3'h6)); forvar59 = (forvar59 + (1'h1)))
        begin
          reg60 <= {$signed((^~($unsigned(wire57) ?
                  $signed(wire54) : $signed(forvar59)))),
              $signed((($unsigned(wire57) & $signed(wire53)) == (((7'h56) != wire55) || ((8'hb6) ^ forvar59))))};
          if (((wire58[(4'h8):(2'h2)] ?
                  ({$unsigned(wire57), $unsigned(wire55)} ?
                      (~^wire54) : forvar59[(2'h3):(2'h3)]) : (&((&reg60) > ((7'h4d) ?
                      wire56 : wire57)))) ?
              (($signed((~&forvar59)) <<< ({reg60} ?
                  $signed(wire58) : (reg60 ?
                      wire58 : wire55))) <= $unsigned(reg60[(4'h8):(3'h4)])) : wire56))
            begin
              reg61 = ($unsigned(wire55) ?
                  wire58 : (&($signed((forvar59 >> (8'ha7))) ?
                      (wire56 <<< (wire56 <= wire55)) : {wire58[(3'h6):(1'h1)],
                          $signed((7'h43)),
                          {wire57, forvar59, forvar59}})));
              reg62 = wire55[(3'h5):(3'h5)];
              reg63 <= wire53[(1'h0):(1'h0)];
              reg64 = $unsigned({(((wire58 ? wire55 : wire55) ?
                          wire53[(1'h1):(1'h1)] : (7'h50)) ?
                      (|$signed(wire54)) : $signed({wire53, (7'h41)})),
                  wire55[(3'h4):(2'h2)],
                  (~$unsigned(reg60))});
            end
          else
            begin
              reg61 = wire54;
              reg63 <= ($unsigned((wire55[(4'ha):(4'h8)] ?
                  $unsigned($unsigned(wire56)) : (wire58[(3'h7):(2'h3)] ~^ (wire53 && wire53)))) ^ ((forvar59 ?
                  $signed((wire56 <= wire58)) : $signed((reg60 + wire58))) ^ {(((8'hbc) ?
                          wire55 : reg64) ?
                      $unsigned(reg64) : $signed(wire56)),
                  (~^((7'h4b) ? (7'h4d) : wire57))}));
              reg65 <= reg63;
              reg66 <= wire58[(3'h5):(3'h4)];
              reg67 = ((+(~^(~&reg60))) && (&(!{(8'ha9), wire57, reg63})));
              reg68 = $unsigned($signed(({(&reg65)} ?
                  (wire56 >> reg65) : $signed($signed(wire54)))));
            end
          if ((!($unsigned($signed(((8'hb6) & wire55))) ?
              wire56[(3'h5):(1'h0)] : reg62)))
            begin
              reg69 = (reg60[(4'h8):(2'h2)] <= ((((~reg64) ?
                  (wire54 ?
                      (7'h50) : wire58) : $signed(wire54)) > $signed({reg68})) ^ (((~reg60) <<< wire55) ?
                  $signed((reg68 ? reg68 : wire53)) : (~$signed(wire57)))));
              reg70 = (~^reg63);
              reg71 = ((reg65 || (~^{(reg60 + reg61),
                      $unsigned((8'haf)),
                      (wire53 ? reg60 : reg66)})) ?
                  ($signed((8'hbe)) ?
                      forvar59 : $signed($unsigned({reg60,
                          (7'h51),
                          wire55}))) : $unsigned({(reg65[(1'h0):(1'h0)] > {wire56,
                          (8'hb0)})}));
              reg72 <= (^~{reg68[(4'ha):(1'h0)],
                  ((~^reg64) ?
                      $unsigned($signed(reg69)) : reg67[(3'h5):(3'h5)])});
              reg73 <= wire55[(4'hf):(4'hc)];
              reg74 = $unsigned(wire53);
            end
          else
            begin
              reg72 <= (^reg68);
              reg74 = $unsigned((reg71 ?
                  {(~&(&reg72)),
                      {(reg64 ? reg66 : reg66),
                          wire55[(4'hd):(3'h5)],
                          ((8'hb3) != reg73)},
                      ($unsigned((8'h9f)) & ((8'hbd) ?
                          wire57 : wire55))} : ((-(~^reg74)) ?
                      ($unsigned(reg67) ?
                          $signed(forvar59) : $signed(reg64)) : reg72[(5'h15):(5'h13)])));
              reg75 = (~$unsigned({(-$unsigned((7'h53)))}));
              reg76 = reg65[(2'h2):(2'h2)];
              reg77 = reg64[(5'h11):(5'h10)];
              reg78 <= {reg62[(4'hd):(4'h8)]};
              reg79 = (wire54 ?
                  $signed((($signed(reg76) >> (^wire56)) < reg72)) : ($signed(wire57) ?
                      (~&$unsigned($unsigned(reg72))) : ($unsigned(reg60) ?
                          $signed(reg72) : ((reg69 > reg67) <= reg60))));
            end
          reg80 = {(((^~(reg66 ?
                      reg66 : wire54)) * ($unsigned((8'ha8)) - (~&reg64))) ?
                  (~(reg65 ?
                      $signed(reg79) : $unsigned(reg68))) : $unsigned(wire55)),
              reg65};
          reg81 = $unsigned(($signed($signed(reg66[(1'h1):(1'h0)])) ?
              ({reg66} != wire53[(3'h5):(2'h2)]) : ((-(reg74 ?
                  wire53 : (7'h46))) * ((reg79 ? reg65 : wire56) ?
                  $unsigned(reg66) : (reg64 >= (7'h47))))));
          for (forvar82 = (1'h0); (forvar82 < (3'h4)); forvar82 = (forvar82 + (1'h1)))
            begin
              reg83 <= $signed($unsigned(reg76));
              reg84 <= (reg76 ?
                  $signed((reg74 <<< ((reg69 ?
                      reg79 : wire58) + reg60))) : ((+(+reg79[(3'h4):(2'h2)])) ?
                      ($signed((reg65 ?
                          reg63 : wire53)) ^~ $signed(reg75)) : reg78));
            end
          reg85 <= (&$signed({$unsigned(reg79[(2'h3):(1'h1)]),
              {((8'hbb) + (7'h42))}}));
        end
      reg86 = (~reg63[(1'h1):(1'h0)]);
    end
  assign wire87 = ({$signed((-reg72)),
                          reg73,
                          ($unsigned($signed(reg63)) ?
                              (8'hb7) : (|(reg72 ? wire58 : wire54)))} ?
                      $unsigned($signed(((reg60 ~^ reg65) ^ $unsigned(reg72)))) : {reg84[(3'h4):(1'h1)],
                          reg60});
  always
    @(posedge clk) begin
      for (forvar88 = (1'h0); (forvar88 < (2'h2)); forvar88 = (forvar88 + (1'h1)))
        begin
          reg89 = ({(~$unsigned(reg78))} ?
              ($unsigned($signed((wire54 - reg72))) != (reg72 >= ((wire57 ^ reg63) >> (wire57 ?
                  reg63 : reg83)))) : ((({(8'hab)} <= $signed(reg63)) ?
                  (((7'h57) ?
                      wire54 : wire58) == $signed(wire58)) : reg60[(3'h6):(1'h0)]) * (wire53 >>> $unsigned((wire57 ?
                  reg72 : wire55)))));
          reg90 <= reg84;
          reg91 <= (~|($signed((reg78[(4'hf):(1'h1)] ?
                  (^reg84) : $unsigned(reg63))) ?
              $unsigned(({reg63, wire57, wire56} ?
                  (8'hb6) : (reg90 ? reg60 : wire57))) : $signed(reg73)));
          reg92 <= (((8'h9c) ?
              $unsigned(((+wire58) - {(8'ha0),
                  reg90})) : wire58[(4'h9):(4'h8)]) > wire53);
        end
      if ((reg85 || reg83[(5'h1a):(4'hc)]))
        begin
          reg93 <= {(~&(reg84[(3'h7):(3'h7)] | ((reg85 << wire54) ?
                  (reg60 > (8'hbb)) : ((8'hab) - reg65))))};
        end
      else
        begin
          for (forvar93 = (1'h0); (forvar93 < (3'h6)); forvar93 = (forvar93 + (1'h1)))
            begin
              reg94 <= (wire57 & (-$signed(reg91)));
              reg95 = $unsigned((reg78[(4'he):(4'hb)] ?
                  {($unsigned(reg90) ? (|reg65) : ((7'h40) != (7'h41))),
                      $unsigned(wire87),
                      $unsigned($unsigned(reg66))} : reg90[(1'h1):(1'h0)]));
              reg96 = wire56[(4'hc):(3'h7)];
              reg97 <= {((reg72 + reg60[(2'h2):(1'h0)]) < $unsigned(((reg60 ^~ (7'h53)) ?
                      $unsigned(reg72) : reg73))),
                  $unsigned(reg94)};
              reg98 <= (~|(reg94 ?
                  $signed(($signed(reg95) * $signed((7'h4b)))) : $unsigned((8'ha5))));
              reg99 <= (reg73 ? $signed(reg89) : reg94[(3'h5):(2'h3)]);
              reg100 <= $signed(reg98);
            end
        end
      if ((~&$unsigned(($signed(reg99[(4'h8):(1'h1)]) <= $unsigned($signed(reg92))))))
        begin
          if ($unsigned($unsigned((+reg93))))
            begin
              reg101 <= {reg96[(2'h3):(1'h1)]};
              reg102 = {reg98};
            end
          else
            begin
              reg101 <= $signed(($unsigned(($unsigned(reg91) + (reg100 ?
                  wire56 : reg65))) || reg65));
              reg103 <= (wire54 ? reg89 : reg95);
            end
          if ($signed($unsigned($unsigned((reg94[(1'h1):(1'h1)] ~^ (reg91 - reg93))))))
            begin
              reg104 <= (reg99 ?
                  ($unsigned(reg66) ^~ (|$unsigned(reg100[(1'h1):(1'h0)]))) : $unsigned((+(reg78 ?
                      {(8'hab), wire55, (8'haf)} : (|forvar88)))));
              reg105 <= reg60;
              reg106 = reg101[(3'h7):(2'h2)];
            end
          else
            begin
              reg104 <= (-{(~|((forvar93 ?
                      forvar93 : wire57) == $unsigned(wire58)))});
              reg106 = $unsigned(forvar93);
              reg107 = forvar88[(3'h6):(3'h6)];
              reg108 = $signed(reg78[(4'hb):(2'h2)]);
              reg109 = $signed(reg99[(4'hc):(3'h7)]);
            end
          reg110 <= (^$signed(wire57[(1'h1):(1'h0)]));
          reg111 <= wire57[(4'h8):(2'h2)];
          if ((~reg95[(3'h6):(3'h6)]))
            begin
              reg112 <= reg94;
              reg113 <= (($signed((~&(wire53 != reg112))) ?
                      reg65[(2'h3):(2'h2)] : ((&$signed(reg65)) >= {(reg103 ?
                              (7'h52) : reg108)})) ?
                  reg99 : reg66[(3'h4):(1'h0)]);
              reg114 = $unsigned((^~wire56));
              reg115 <= reg98;
              reg116 <= {reg78[(4'hd):(2'h3)], reg109, reg97[(2'h2):(2'h2)]};
            end
          else
            begin
              reg114 = ($signed(reg101[(1'h1):(1'h0)]) ?
                  reg73 : (wire55[(3'h4):(2'h2)] ?
                      (~&$unsigned((~&reg94))) : (-$unsigned((reg98 ?
                          reg105 : (7'h52))))));
              reg117 = reg78;
            end
        end
      else
        begin
          if (reg115[(4'hd):(4'h8)])
            begin
              reg101 <= reg94[(4'hf):(4'hb)];
            end
          else
            begin
              reg102 = $signed(reg89);
              reg103 <= reg111[(5'h18):(1'h0)];
              reg104 <= ($unsigned(reg115[(5'h15):(1'h1)]) ?
                  reg107 : $unsigned(wire58));
            end
          for (forvar105 = (1'h0); (forvar105 < (2'h3)); forvar105 = (forvar105 + (1'h1)))
            begin
              reg106 = (({({reg107, reg103} - $unsigned(reg96))} ^ reg89) ?
                  ($signed($unsigned((reg116 << reg83))) ?
                      (!{{reg89, (8'hb4)},
                          $signed((8'hac)),
                          $unsigned(reg93)}) : ((^$signed(reg115)) ?
                          reg78[(4'hb):(1'h1)] : {$signed(reg85)})) : (reg84 < (8'hba)));
              reg110 <= ($unsigned((8'h9c)) ?
                  (~^$unsigned(($signed(reg111) ?
                      reg94 : reg111))) : reg109[(3'h7):(3'h5)]);
              reg114 = reg101;
              reg117 = ($signed($signed(reg93)) ?
                  ((reg96 ?
                      ({wire87, reg110} ?
                          reg110 : (8'hb4)) : reg108[(4'h9):(2'h2)]) >= reg93[(5'h10):(3'h6)]) : $unsigned(reg109));
            end
          reg118 <= ((reg65[(2'h2):(1'h0)] ?
              $signed(($unsigned((7'h4c)) ?
                  reg94 : $signed(reg116))) : $unsigned((~&reg94))) != (~^forvar88[(2'h3):(2'h2)]));
          reg119 <= reg104;
          for (forvar120 = (1'h0); (forvar120 < (1'h0)); forvar120 = (forvar120 + (1'h1)))
            begin
              reg121 <= ((~^$unsigned(reg118[(2'h2):(1'h0)])) ?
                  ((reg83[(3'h6):(1'h0)] | (7'h52)) >>> reg91[(2'h3):(2'h2)]) : $signed($unsigned(reg63)));
              reg122 = $signed(reg66[(3'h6):(1'h1)]);
              reg123 <= $signed($unsigned((wire57[(4'h9):(1'h0)] ?
                  reg60[(3'h5):(3'h5)] : reg119[(5'h14):(3'h6)])));
              reg124 <= (8'ha9);
              reg125 = (~|reg110);
              reg126 <= $unsigned($unsigned(($unsigned(reg122[(1'h1):(1'h1)]) ?
                  ((reg92 ? reg83 : reg107) ?
                      ((7'h47) & reg96) : (reg97 ? reg102 : reg93)) : wire53)));
              reg127 = (8'h9d);
            end
        end
      reg128 = reg126;
      for (forvar129 = (1'h0); (forvar129 < (3'h6)); forvar129 = (forvar129 + (1'h1)))
        begin
          for (forvar130 = (1'h0); (forvar130 < (3'h4)); forvar130 = (forvar130 + (1'h1)))
            begin
              reg131 <= $signed($signed(reg90[(1'h0):(1'h0)]));
              reg132 <= forvar129;
              reg133 = ($unsigned(reg102[(3'h6):(3'h6)]) ?
                  reg83 : {$signed({(reg78 ? forvar88 : reg92)}), (7'h43)});
              reg134 <= reg99[(4'hc):(3'h7)];
              reg135 = (($unsigned($unsigned(((7'h51) == reg103))) ?
                  ($signed(reg101) > ((8'ha5) <= reg131[(3'h4):(3'h4)])) : reg124) == ($signed($unsigned((~^forvar105))) + (^~$unsigned((~|reg104)))));
            end
          reg136 <= reg92;
          if ({$unsigned(reg113[(1'h1):(1'h1)]),
              reg66,
              {($signed((reg106 ? reg65 : reg110)) ?
                      $unsigned($unsigned(wire55)) : $unsigned((reg136 ?
                          reg108 : reg65)))}})
            begin
              reg137 = ({(~|$unsigned($signed(reg98))),
                      {(~&forvar129[(2'h2):(1'h0)])},
                      $signed((reg91 - (&reg102)))} ?
                  wire54[(4'hb):(4'ha)] : $unsigned(((reg92 <<< reg109) ?
                      {$signed(reg60)} : ($signed(reg119) & reg92))));
            end
          else
            begin
              reg138 <= forvar120[(2'h3):(1'h1)];
              reg139 = $signed((($signed(reg100[(1'h0):(1'h0)]) ?
                  reg117[(4'hb):(3'h7)] : (|(~&reg98))) <<< (~&((~reg103) ?
                  reg107 : (reg73 == reg89)))));
              reg140 = (~&$signed({(!$signed(reg114))}));
              reg141 = (reg110[(3'h5):(1'h1)] ?
                  (reg83[(5'h1a):(3'h7)] ^ reg63[(1'h0):(1'h0)]) : ($signed(reg105) ?
                      reg99[(4'hd):(1'h0)] : (+reg90)));
              reg142 <= (~&{(|($signed(reg108) >= (reg96 ? reg124 : reg137))),
                  reg121[(4'hc):(4'h8)],
                  (|$unsigned((reg124 >>> reg104)))});
              reg143 <= (($unsigned((-reg60[(1'h1):(1'h0)])) * ((reg65[(1'h1):(1'h1)] < reg92) ?
                  $unsigned(reg126) : reg103)) ^ $unsigned(((~(reg84 ^ reg94)) ?
                  reg89 : ((7'h41) < $signed(wire56)))));
            end
          for (forvar144 = (1'h0); (forvar144 < (3'h4)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 = ((($signed(reg138[(3'h4):(2'h2)]) || (+(forvar88 << reg92))) | $unsigned($signed($unsigned(reg138)))) || reg98[(5'h19):(1'h1)]);
              reg146 <= (&(((+(~&reg126)) ?
                  ($signed(wire54) - $signed(reg121)) : {$unsigned(reg119)}) - (wire87 ?
                  (~^(reg117 ?
                      forvar105 : reg135)) : $signed(reg124[(4'hb):(3'h4)]))));
              reg147 <= (~&($unsigned((^~$unsigned((8'hbe)))) ?
                  $unsigned($unsigned(reg142[(1'h1):(1'h1)])) : (~&(7'h49))));
              reg148 <= ($signed((reg141 & wire56)) || ((((reg73 ?
                      reg117 : reg96) ?
                  reg93[(1'h0):(1'h0)] : $signed(forvar120)) && $signed($unsigned(reg65))) == reg116));
              reg149 = (^~reg73);
              reg150 = ($signed({{reg60, (8'hac), reg149}}) ?
                  ($signed(reg140) ?
                      $unsigned(((reg91 ?
                          reg96 : reg136) && (^(7'h54)))) : forvar120[(3'h7):(3'h6)]) : ((reg121[(5'h1a):(5'h14)] & reg83) ?
                      $unsigned(reg91) : (7'h57)));
              reg151 = (+((8'hb1) >>> reg100));
            end
          reg152 = $signed($unsigned(forvar93[(4'ha):(3'h7)]));
        end
      reg153 = ($unsigned(reg115) ?
          ((8'hb2) >> (+($unsigned(reg90) << reg89[(4'he):(1'h1)]))) : ((((reg105 + reg139) ?
                  (reg142 ?
                      (8'hb0) : reg65) : (reg149 + reg126)) == (~|((7'h52) ?
                  reg85 : reg102))) ?
              (+reg127[(4'hb):(4'h9)]) : (+((reg78 ? reg111 : forvar144) ?
                  (8'h9f) : wire87))));
    end
  assign wire154 = reg146;
  assign wire155 = $unsigned($unsigned((((reg72 | (8'h9c)) ?
                       $signed(reg138) : (-(8'h9c))) <= (^~$unsigned(reg92)))));
  assign wire156 = (!{$unsigned((!((7'h45) ? reg147 : reg99)))});
  assign wire157 = (|reg132[(4'hf):(4'hb)]);
  always
    @(posedge clk) begin
      reg158 = ((!($signed((^(7'h54))) ?
          (reg85[(5'h13):(5'h12)] * {reg111,
              wire87,
              (7'h40)}) : (~&$unsigned((7'h50))))) * reg101);
      reg159 <= reg91[(4'ha):(3'h7)];
      reg160 <= $unsigned(({$signed($unsigned(reg118)),
          $unsigned($signed((7'h41)))} >> reg158[(3'h6):(3'h4)]));
      for (forvar161 = (1'h0); (forvar161 < (3'h4)); forvar161 = (forvar161 + (1'h1)))
        begin
          if ((~^$unsigned($unsigned($signed(wire55)))))
            begin
              reg162 = $unsigned(((+(^(8'hbe))) ?
                  reg148[(4'he):(2'h3)] : wire53));
              reg163 = $signed($signed(($signed(reg159) + ((-reg138) ?
                  {(7'h4a), reg84} : (~^reg84)))));
              reg164 = {(~(~wire57))};
              reg165 = {(((reg92[(4'hc):(4'h9)] ~^ wire87[(4'hc):(4'ha)]) ?
                          ($signed((8'h9c)) == reg134[(4'hb):(1'h0)]) : $unsigned(((7'h54) * (8'hbd)))) ?
                      $unsigned(wire56[(4'h8):(3'h4)]) : ($unsigned((!reg78)) >> ((|reg105) ?
                          (wire155 ? reg63 : reg136) : ((7'h42) ?
                              reg85 : reg90)))),
                  $unsigned(wire156[(3'h7):(1'h1)])};
              reg166 <= $unsigned({reg73, {$unsigned(reg159)}});
              reg167 <= $signed(reg143);
              reg168 = {{((reg90 | (reg126 && forvar161)) ?
                          (^wire155[(3'h7):(1'h1)]) : wire157),
                      (reg90 ^~ ({(8'hb1),
                          reg158,
                          reg121} & $unsigned((8'ha3)))),
                      (&({wire156, reg116} ?
                          $unsigned(reg90) : $signed(reg142)))}};
            end
          else
            begin
              reg166 <= (~|reg148);
              reg167 <= (reg118 || (reg132[(2'h2):(1'h1)] ?
                  {reg136,
                      $unsigned($unsigned(reg92))} : $signed($unsigned($signed(reg124)))));
              reg168 = $unsigned(reg163);
            end
          reg169 = wire53;
          reg170 = (reg112 > ((((reg134 ? reg93 : reg121) <<< (~(8'ha4))) ?
              (!(reg100 ?
                  reg60 : reg65)) : ($unsigned(reg72) <= (~&reg159))) <<< $unsigned((|$signed(wire53)))));
          for (forvar171 = (1'h0); (forvar171 < (3'h6)); forvar171 = (forvar171 + (1'h1)))
            begin
              reg172 <= reg124;
              reg173 <= reg132[(3'h5):(1'h1)];
              reg174 <= reg148;
              reg175 <= $unsigned(reg72[(5'h19):(3'h6)]);
              reg176 = $unsigned(((reg65 >> ((~|wire56) == $signed(wire157))) ?
                  {({(7'h48)} + wire57[(3'h5):(1'h0)])} : reg170[(1'h1):(1'h0)]));
              reg177 <= reg136;
            end
          reg178 <= $signed((+wire155[(2'h3):(1'h0)]));
        end
    end
  module179 #() modinst314 (.wire180(wire155), .wire181(reg78), .wire182(reg103), .wire183(reg126), .y(wire313), .wire185(reg110), .clk(clk), .wire184(wire157));
  always
    @(posedge clk) begin
      reg315 = reg138[(1'h0):(1'h0)];
      for (forvar316 = (1'h0); (forvar316 < (3'h6)); forvar316 = (forvar316 + (1'h1)))
        begin
          reg317 = reg104[(5'h10):(4'h8)];
        end
      if ($signed($signed($unsigned((wire58 ~^ reg315)))))
        begin
          reg318 = (($unsigned({(reg159 != (8'ha6)), reg174}) ?
                  reg105[(4'he):(3'h4)] : reg92) ?
              ((|($unsigned(reg65) ? reg101 : wire57)) ?
                  (((wire87 ? reg112 : wire56) & (reg103 >= reg148)) ?
                      {$signed(reg178),
                          {reg99,
                              wire56}} : (^~(!reg99))) : {reg126[(4'hd):(3'h6)],
                      ($signed(reg110) & $signed(reg94)),
                      ($signed(reg126) - reg148[(5'h18):(4'ha)])}) : ((reg91[(1'h0):(1'h0)] ^ {$signed((8'h9f)),
                  (~(8'ha3))}) - (~|(~$unsigned(reg116)))));
          for (forvar319 = (1'h0); (forvar319 < (3'h4)); forvar319 = (forvar319 + (1'h1)))
            begin
              reg320 = ($signed($signed(reg105[(4'hc):(2'h2)])) ?
                  reg147 : ($signed({wire58[(4'ha):(3'h4)], $signed(reg65)}) ?
                      (~(+$unsigned(wire54))) : {((wire313 <= wire58) ?
                              (~|reg160) : $unsigned(reg91))}));
              reg321 = ((&($unsigned(reg92[(4'h8):(3'h7)]) ?
                  ((reg124 ? reg146 : reg147) ?
                      reg318[(5'h15):(1'h1)] : (~&reg100)) : $unsigned((reg175 & (7'h4f))))) ~^ reg118[(4'he):(4'hb)]);
              reg322 <= (~&reg101);
              reg323 = reg132[(1'h1):(1'h0)];
              reg324 = ({(~$signed((reg90 ? reg166 : forvar316))),
                      $unsigned((~|$signed(reg177))),
                      reg174} ?
                  ((+(+(8'ha9))) * (reg110[(3'h5):(3'h4)] ?
                      ((reg60 + reg174) ?
                          $signed((7'h55)) : (-(8'ha1))) : $unsigned((wire56 ?
                          reg85 : wire57)))) : $unsigned($signed(reg63)));
            end
          if ($unsigned(reg94))
            begin
              reg325 <= {(reg101[(3'h6):(1'h1)] & {reg100, wire56}),
                  reg172,
                  (+$unsigned({(~^reg72), ((8'ha9) ? reg94 : reg142), reg85}))};
              reg326 <= ({reg115[(3'h6):(2'h3)],
                      $unsigned($signed({forvar319}))} ?
                  ({(^(wire56 + (8'haa)))} * ((|reg112) * (^(|(7'h42))))) : {{(((8'hba) ?
                              reg103 : forvar316) || $signed(reg142))},
                      (~&reg113),
                      $unsigned(reg132[(4'h8):(1'h1)])});
              reg327 <= ($unsigned((^$unsigned((reg178 ?
                  reg104 : reg175)))) - wire55[(1'h0):(1'h0)]);
              reg328 = {(+($unsigned({reg101}) ?
                      reg327[(4'hb):(2'h3)] : (reg119 ?
                          $unsigned(reg98) : reg116))),
                  $signed((~^$signed($unsigned(wire156))))};
              reg329 = ($signed($unsigned($signed($unsigned((8'ha9))))) < reg324);
              reg330 <= $signed({((reg90[(1'h0):(1'h0)] ?
                      (reg111 != reg147) : $unsigned(reg103)) ^~ ((~&(8'hb4)) ^~ wire55[(4'hd):(4'h8)])),
                  {((reg112 ? reg123 : reg147) ? (~^wire58) : (+reg112)),
                      (&(wire55 | forvar319))}});
            end
          else
            begin
              reg325 <= $signed($signed({reg167[(5'h10):(4'hb)],
                  (reg329[(2'h3):(1'h1)] ?
                      $signed(reg85) : $signed((8'ha1)))}));
              reg326 <= $signed(({$unsigned((wire55 ? reg72 : wire154)),
                      $unsigned($signed(reg142)),
                      $signed($unsigned(reg103))} ?
                  reg116[(5'h10):(4'h8)] : $signed(reg323)));
              reg327 <= reg315;
            end
        end
      else
        begin
          reg318 = ((($signed(wire155[(1'h0):(1'h0)]) ^~ {$unsigned(reg325)}) ?
              {((~^(8'hbd)) >> ((8'haf) ~^ reg325))} : $signed(($signed(wire53) + ((7'h41) && reg111)))) && (reg63 <= $signed(((~^reg321) ^~ (reg173 * (7'h56))))));
          for (forvar319 = (1'h0); (forvar319 < (3'h4)); forvar319 = (forvar319 + (1'h1)))
            begin
              reg320 = $unsigned(((&(&(wire53 ? reg110 : reg100))) ?
                  (wire55[(1'h1):(1'h1)] <= $unsigned((7'h4a))) : (reg132 >> reg85)));
              reg322 <= (((reg113[(2'h3):(1'h0)] & $signed(reg78[(4'hf):(1'h1)])) ?
                  reg124[(3'h6):(3'h6)] : {(^~((7'h4f) >>> reg105)),
                      ((reg84 ? (8'hae) : reg148) ?
                          $unsigned(reg66) : (reg167 <<< reg113)),
                      reg167}) ^ $unsigned($unsigned((wire57 ?
                  reg60 : reg93))));
              reg325 <= reg330[(5'h10):(3'h5)];
              reg328 = (&wire157);
              reg329 = {{(~{(~|reg116)}), reg132}, reg330[(5'h1c):(5'h1b)]};
            end
          if (((reg113 << $unsigned($unsigned({reg321, (7'h4c)}))) ?
              (&$unsigned(reg315[(3'h5):(1'h1)])) : ((-$signed(reg166[(2'h2):(1'h1)])) | $signed(reg167[(3'h4):(1'h0)]))))
            begin
              reg330 <= $unsigned($unsigned(reg147[(3'h4):(1'h0)]));
              reg331 <= ($signed({$signed((reg328 ? (8'hba) : (8'ha7))),
                  reg105[(4'h8):(3'h7)],
                  reg63[(1'h0):(1'h0)]}) == reg126[(3'h4):(2'h2)]);
              reg332 = (|((reg112[(5'h10):(3'h6)] >> $signed((reg177 ?
                      reg111 : (8'ha6)))) ?
                  (-((reg83 == reg330) ?
                      (~reg85) : (reg177 != reg98))) : (wire155 ?
                      (!(7'h4e)) : $signed($signed(reg124)))));
            end
          else
            begin
              reg330 <= (^~$signed(((((8'hb3) - reg118) > $signed(reg119)) + (+reg325[(1'h0):(1'h0)]))));
              reg331 <= ({(^(8'h9d))} >>> reg105);
              reg332 = wire154[(4'he):(3'h6)];
              reg333 = (reg85[(4'hf):(2'h3)] ^ reg330);
            end
          reg334 = $unsigned(reg172);
          for (forvar335 = (1'h0); (forvar335 < (3'h6)); forvar335 = (forvar335 + (1'h1)))
            begin
              reg336 = (~^{reg334[(5'h10):(3'h4)]});
            end
          reg337 <= $unsigned((reg332[(2'h2):(1'h1)] | $signed($signed(reg110))));
        end
      if (reg110)
        begin
          reg338 <= (^$signed((((~^reg332) * (reg174 ? reg119 : (8'hba))) ?
              forvar335 : (+$signed(reg72)))));
          reg339 = (reg325 ?
              {(~&wire57[(5'h12):(4'ha)]),
                  reg78,
                  {(~$unsigned(wire56)), (7'h51)}} : reg175[(4'he):(4'h9)]);
          for (forvar340 = (1'h0); (forvar340 < (3'h4)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 = reg123[(4'h9):(3'h5)];
              reg342 <= $signed((~|reg167[(5'h17):(3'h7)]));
              reg343 = ((-$unsigned($unsigned(forvar335[(2'h2):(1'h1)]))) || (wire313[(5'h12):(4'h8)] ~^ reg103[(5'h12):(1'h0)]));
              reg344 = ({$signed(((reg142 ? reg327 : reg322) ?
                      $unsigned(reg341) : $unsigned((8'hab)))),
                  (|reg160)} << $signed(reg73[(1'h1):(1'h1)]));
              reg345 <= $signed(wire313);
            end
          reg346 <= reg83;
          reg347 <= reg143[(3'h5):(1'h0)];
        end
      else
        begin
          reg339 = reg321;
        end
    end
  assign wire348 = $unsigned(reg85[(1'h0):(1'h0)]);
  assign wire349 = {(reg142[(5'h12):(3'h7)] ? reg175 : reg326[(4'h9):(1'h0)]),
                       (wire53[(2'h3):(2'h2)] & ($unsigned((reg84 ?
                           reg97 : wire156)) <<< ((~reg91) ?
                           (7'h4e) : $unsigned(reg118)))),
                       reg110};
  assign wire350 = $unsigned(reg103[(4'hd):(4'hc)]);
  always
    @(posedge clk) begin
      reg351 = (((((wire55 >> reg138) ? reg178 : reg112[(4'hb):(2'h2)]) ?
                  wire156 : reg118[(3'h7):(3'h7)]) ?
              $unsigned(reg85) : (!reg91[(3'h5):(3'h4)])) ?
          ((reg136 ?
              (((8'ha5) < wire154) ? reg90 : wire349) : $unsigned((reg330 ?
                  reg93 : reg345))) > (($signed((7'h54)) & (reg166 ?
              reg126 : reg84)) != (+(reg173 >> reg325)))) : ((^reg119) ^~ {reg138,
              (!wire348)}));
      for (forvar352 = (1'h0); (forvar352 < (1'h1)); forvar352 = (forvar352 + (1'h1)))
        begin
          for (forvar353 = (1'h0); (forvar353 < (1'h1)); forvar353 = (forvar353 + (1'h1)))
            begin
              reg354 = $signed(wire350);
              reg355 <= wire55[(4'h8):(3'h5)];
            end
          for (forvar356 = (1'h0); (forvar356 < (3'h6)); forvar356 = (forvar356 + (1'h1)))
            begin
              reg357 <= $unsigned($signed((-($signed(reg73) ?
                  (!reg92) : (+(8'ha8))))));
              reg358 = $unsigned($signed(((8'hb6) ?
                  wire157 : (|(wire57 ^ reg119)))));
              reg359 = $unsigned(((!((7'h54) ?
                      $signed(reg131) : (wire55 ? reg84 : reg146))) ?
                  $unsigned({(reg103 & reg159)}) : (($unsigned(reg354) ?
                      $signed((8'hbc)) : (wire53 ?
                          (7'h45) : reg113)) >>> reg111[(5'h13):(2'h3)])));
              reg360 = {reg346[(4'hb):(2'h2)]};
              reg361 = ($unsigned($signed(($signed(wire157) < $unsigned(reg115)))) >> $signed(reg116));
              reg362 = reg97;
            end
          if ((($signed($signed(reg345)) ?
                  (reg351 ?
                      (&{reg159,
                          reg142,
                          reg136}) : ($unsigned(reg166) << reg143)) : reg178[(4'hb):(3'h7)]) ?
              (~^$unsigned({reg326})) : reg60[(3'h5):(1'h0)]))
            begin
              reg363 <= reg331[(1'h1):(1'h0)];
              reg364 = (!($signed({(reg72 ? (7'h55) : reg160), wire55}) ?
                  reg78 : $signed(((~&(8'hba)) ? reg147 : forvar352))));
              reg365 = {((8'hbc) ?
                      $signed(reg83) : ($unsigned((reg72 ^ reg66)) ?
                          $unsigned((wire350 ? wire87 : reg177)) : reg99)),
                  reg354,
                  ({(~^(reg73 ?
                          forvar356 : reg142))} >= (wire157 + $unsigned((reg103 ?
                      (8'ha4) : wire349))))};
            end
          else
            begin
              reg364 = reg100[(1'h1):(1'h1)];
              reg366 <= ($signed((($unsigned(reg322) ?
                      reg360[(1'h0):(1'h0)] : $signed(reg90)) && reg115)) ?
                  $unsigned(reg123[(3'h7):(3'h7)]) : $unsigned(($signed(reg360[(1'h1):(1'h1)]) ?
                      ({reg146} < (reg99 & wire58)) : (reg121[(4'h9):(3'h6)] ^~ reg178))));
              reg367 <= $signed(reg104[(4'he):(3'h4)]);
            end
          if (($unsigned(reg357) - (8'haa)))
            begin
              reg368 <= ((7'h55) >>> $signed($unsigned(($unsigned((8'ha1)) ?
                  reg337 : reg327))));
              reg369 = ($signed($unsigned($unsigned((reg175 ?
                      reg63 : reg330)))) ?
                  (~^reg368) : (|(($signed(reg325) ^ reg363[(5'h13):(5'h12)]) ?
                      ($signed(reg366) ^~ reg78[(4'hb):(4'h8)]) : (^~(wire87 & wire349)))));
            end
          else
            begin
              reg369 = reg359[(5'h17):(3'h6)];
              reg370 <= reg90;
            end
          reg371 = (reg359 & ($unsigned($signed($signed(reg134))) ?
              $signed($signed((wire53 ? reg115 : reg177))) : ((~^((8'hb4) ?
                  reg347 : reg360)) ^ (~^(reg126 & reg65)))));
          if ($unsigned(wire349))
            begin
              reg372 <= $signed($unsigned(reg174[(3'h5):(3'h4)]));
              reg373 <= $signed($signed(reg83));
              reg374 = {reg342[(3'h4):(1'h1)],
                  {($unsigned((reg105 ? reg351 : reg138)) >>> (reg126 ?
                          $signed((7'h43)) : $signed(reg85))),
                      reg355}};
            end
          else
            begin
              reg374 = {(&wire154[(2'h2):(1'h1)])};
              reg375 = $signed((|$signed($signed(reg372[(5'h13):(3'h7)]))));
              reg376 = $unsigned(reg119[(5'h15):(3'h4)]);
              reg377 = $signed($signed($unsigned($unsigned($unsigned(reg374)))));
              reg378 <= (~&($signed(({(8'haf), (8'h9d)} ?
                      $unsigned(reg361) : ((8'ha5) ? reg85 : reg173))) ?
                  reg331[(2'h2):(2'h2)] : reg159[(2'h2):(1'h0)]));
              reg379 <= ($signed(reg126[(4'ha):(3'h6)]) ?
                  $signed($unsigned((^~(wire313 >= reg100)))) : ((^~(!reg78)) ?
                      reg93 : (((wire156 ? (7'h49) : reg112) ?
                          (-reg358) : reg131) >> (|(reg97 != wire87)))));
              reg380 = $signed(((wire155[(4'hd):(3'h5)] ?
                  reg358[(4'h9):(3'h5)] : $signed($unsigned(forvar356))) && {reg111[(5'h13):(3'h7)],
                  (reg147[(3'h5):(3'h4)] ?
                      (reg142 >>> reg126) : $signed(wire58))}));
            end
        end
      reg381 = reg177;
      if (($unsigned((^$unsigned((|reg367)))) ?
          $unsigned(reg92[(4'hc):(4'hb)]) : reg72[(2'h3):(2'h3)]))
        begin
          reg382 = (((|(reg72[(4'hd):(2'h3)] ?
                  (^(8'ha0)) : $unsigned(reg134))) * reg138) ?
              ((~|((7'h42) ? $unsigned(reg378) : $unsigned(reg121))) ?
                  reg101 : $signed($signed((reg355 ?
                      reg104 : reg94)))) : $signed($unsigned($unsigned(forvar353))));
          reg383 <= ((~|(&($signed(reg322) + (reg351 <= reg105)))) >> (~($signed($signed(reg358)) >>> (-reg105[(3'h6):(2'h2)]))));
          if ($signed((($unsigned($signed(forvar353)) ^~ ({reg347} < (reg94 ?
                  forvar352 : wire54))) ?
              $unsigned((8'h9c)) : ((^(reg121 & wire350)) ?
                  {$unsigned(reg142)} : reg121))))
            begin
              reg384 <= (reg357 + ($unsigned((8'ha1)) ?
                  ((reg377 ? {reg331, wire58} : {(7'h40)}) ?
                      ((reg174 ?
                          (7'h53) : reg136) * $unsigned(wire350)) : (7'h4c)) : reg361[(4'hd):(4'hd)]));
              reg385 <= (($signed(reg381[(1'h0):(1'h0)]) < reg146[(4'hb):(1'h1)]) <= $signed(((reg358 | (reg342 <= reg355)) ?
                  $signed(reg147[(3'h5):(1'h0)]) : (&{reg379}))));
              reg386 = $signed(($unsigned(reg148) ^~ (reg66 ?
                  reg85[(5'h13):(4'h9)] : (-(reg65 >> reg91)))));
              reg387 <= $signed((~|$signed(((8'hbc) ^ (8'ha8)))));
              reg388 <= (($unsigned(reg131) <= ((&reg124) * ((~|(8'hb0)) < (~reg138)))) ~^ ((7'h49) >= $signed((reg167[(1'h1):(1'h0)] - $signed(reg364)))));
              reg389 <= reg103[(4'hd):(4'h8)];
              reg390 <= (^(~&(reg364 >> $unsigned({(8'hbd)}))));
            end
          else
            begin
              reg386 = $unsigned((^{$signed((~&wire157)),
                  ((reg390 * reg354) ? $signed((8'hb6)) : wire348),
                  $signed(reg66)}));
              reg387 <= wire313[(5'h10):(4'hc)];
              reg391 = (&$signed((|$unsigned($signed(reg177)))));
              reg392 = (8'ha5);
              reg393 = $unsigned((reg388[(3'h6):(3'h4)] ?
                  ($unsigned({reg377}) ?
                      ($signed((7'h55)) ?
                          reg373[(1'h1):(1'h0)] : wire57) : ((reg73 ?
                          reg378 : reg100) != (wire154 != reg101))) : (^$signed(((8'ha2) || wire54)))));
              reg394 = $signed((((~|$unsigned((7'h49))) * $signed({(7'h48)})) ?
                  (^{reg100[(1'h1):(1'h0)]}) : (($signed(reg384) ?
                          reg327 : (8'hb1)) ?
                      (~reg91) : $signed($unsigned(reg391)))));
            end
          reg395 <= $unsigned(((&{$signed(reg373)}) ^ wire58));
          for (forvar396 = (1'h0); (forvar396 < (1'h1)); forvar396 = (forvar396 + (1'h1)))
            begin
              reg397 = (^reg374);
              reg398 <= (($signed($signed($unsigned(reg63))) ?
                  $signed(reg110[(1'h1):(1'h1)]) : (!reg347[(5'h12):(3'h5)])) * $signed(forvar356));
              reg399 <= reg99[(4'hc):(4'ha)];
              reg400 = reg112;
              reg401 <= reg65;
              reg402 <= ($signed((~(^~$signed(reg361)))) ^ reg390);
            end
          reg403 <= $unsigned((+$unsigned({(reg326 == reg90)})));
        end
      else
        begin
          if (reg374)
            begin
              reg383 <= wire57[(5'h10):(2'h3)];
              reg384 <= (wire87[(1'h0):(1'h0)] < (((|{reg78,
                      (8'hb9)}) ~^ reg372[(4'hf):(3'h6)]) ?
                  reg327 : (reg401[(4'hd):(4'h9)] ?
                      ((reg363 ? wire53 : reg98) ?
                          $signed(reg100) : (+(8'ha7))) : ((~forvar396) ?
                          (^~reg375) : ((8'ha0) ? reg138 : (7'h4a))))));
            end
          else
            begin
              reg383 <= ((-((reg115[(4'hc):(1'h0)] <= $unsigned(reg174)) ?
                  reg384[(5'h13):(3'h7)] : $unsigned((reg322 ~^ reg369)))) || ({($unsigned(reg368) ?
                      (reg379 ? (8'h9c) : wire57) : (^reg83)),
                  (^~$signed(reg403)),
                  reg369} || (($signed(reg369) ?
                  $signed(reg372) : reg134[(5'h12):(4'hb)]) ~^ ($signed(reg374) ?
                  (reg175 ? reg337 : reg142) : {reg386, reg166}))));
              reg386 = ((reg367[(3'h7):(2'h3)] ?
                  (reg367 ?
                      reg402[(4'h9):(4'h9)] : reg364[(1'h0):(1'h0)]) : $unsigned(((reg355 ?
                      reg394 : (8'hb8)) == (~&reg111)))) >> reg346);
              reg387 <= reg375;
              reg391 = (8'ha5);
              reg392 = $unsigned(({$unsigned({reg91})} == $signed(reg373[(5'h1e):(5'h18)])));
            end
          reg395 <= reg84;
          for (forvar396 = (1'h0); (forvar396 < (3'h6)); forvar396 = (forvar396 + (1'h1)))
            begin
              reg398 <= (wire57 ?
                  reg402[(1'h0):(1'h0)] : (&$signed(((reg338 ?
                          (7'h55) : reg104) ?
                      (reg65 ? (8'haa) : reg326) : $unsigned(wire156)))));
              reg400 = $signed((reg355[(4'h9):(2'h2)] ?
                  wire156 : (reg177[(3'h5):(2'h3)] << wire55)));
            end
          if (reg342)
            begin
              reg401 <= (|$unsigned($signed($unsigned((reg101 ^~ reg113)))));
              reg404 = $unsigned((+(^$signed($signed(reg98)))));
              reg405 <= reg354[(4'hc):(3'h6)];
              reg406 <= (((7'h46) ?
                  reg345 : reg325) || {$signed($unsigned($unsigned(reg118))),
                  $unsigned((&(~^reg175))),
                  ((&{(8'h9e), reg372, reg388}) ^~ {((8'ha7) ?
                          (7'h45) : reg345),
                      ((7'h44) != reg364),
                      {wire87, reg85, reg397}})});
              reg407 = (~|((reg175 ?
                      (~(reg105 && reg380)) : ($unsigned(reg382) ?
                          $unsigned(reg351) : (8'hbb))) ?
                  ($unsigned(reg94) & reg113[(3'h4):(1'h0)]) : (8'hbe)));
            end
          else
            begin
              reg401 <= wire348[(4'h9):(1'h1)];
              reg404 = $unsigned(reg136);
              reg407 = $unsigned($signed(wire349));
              reg408 <= (^(reg104 | wire350[(4'h8):(4'h8)]));
              reg409 <= reg338[(4'h8):(1'h1)];
              reg410 <= reg361[(4'hb):(4'h8)];
              reg411 = $signed({reg124});
            end
          if ($unsigned($signed($unsigned($unsigned({reg377,
              reg368,
              reg103})))))
            begin
              reg412 = (&(~&(&$signed((-wire154)))));
              reg413 = (^~({{{wire87, reg90, reg338},
                      (&reg121),
                      reg377[(4'hb):(3'h4)]},
                  ({reg112, reg357, reg387} >= (8'hb8))} - ($unsigned({(8'haa),
                      reg405,
                      reg338}) ?
                  ((~&reg390) || reg111[(5'h16):(3'h6)]) : reg121[(5'h15):(1'h0)])));
              reg414 <= $signed(reg331[(2'h2):(1'h0)]);
              reg415 <= {((~&{((8'hbb) * reg84)}) < $unsigned((|$signed(reg73)))),
                  reg126,
                  $signed($unsigned(((^~(7'h55)) ?
                      reg60[(3'h5):(1'h0)] : (reg72 * reg136))))};
              reg416 = ($unsigned((+((reg146 | reg392) ?
                  $unsigned((8'hab)) : wire156))) >> (reg412[(3'h7):(3'h4)] & $signed(reg366[(4'he):(4'hc)])));
              reg417 <= (wire157 ^ ((&$signed($signed(reg405))) ?
                  ($signed((reg345 & reg78)) ?
                      ($signed(reg85) >> (7'h43)) : $unsigned((reg338 ?
                          wire349 : reg105))) : ((&reg358) ?
                      (!{reg361,
                          reg363,
                          (7'h47)}) : $signed((reg410 * reg132)))));
            end
          else
            begin
              reg414 <= $signed(($unsigned($unsigned(reg121[(5'h18):(5'h11)])) ?
                  (reg394[(4'hc):(1'h0)] < reg365[(4'h9):(3'h7)]) : reg357));
              reg416 = $signed(((-((reg110 >= reg415) <= $unsigned((8'hb4)))) == reg131));
              reg417 <= {reg97[(2'h3):(1'h1)], reg138[(3'h5):(3'h5)]};
              reg418 = $signed(((+(wire87[(2'h3):(1'h1)] != $unsigned((8'ha5)))) ?
                  $signed({$signed(reg115)}) : (reg118[(5'h11):(3'h6)] ?
                      {(reg354 && reg394),
                          (reg63 >= (8'hae))} : {$unsigned((7'h56))})));
              reg419 <= $unsigned((reg414 ?
                  $unsigned(reg382) : (((wire56 ? reg358 : (7'h4e)) ?
                      (wire55 ?
                          reg366 : reg121) : reg90[(1'h0):(1'h0)]) < ($unsigned(reg413) ?
                      $signed(reg131) : (wire349 ? reg365 : reg105)))));
              reg420 = ($unsigned({reg85,
                      {(reg414 ? reg388 : (8'hb9)), (~|reg419)}}) ?
                  (^~(reg345 ?
                      $signed(((8'h9c) ?
                          (8'had) : (8'hb0))) : (~^(+reg375)))) : $unsigned({{(reg116 ?
                              reg389 : reg98),
                          $unsigned((7'h57))},
                      (reg398 < (wire54 ? reg173 : reg105)),
                      wire57}));
              reg421 <= ($unsigned((reg345[(2'h2):(2'h2)] ?
                  (~&(reg72 ?
                      reg399 : reg401)) : wire157[(2'h3):(2'h2)])) == (~($unsigned({reg338,
                  (8'ha7)}) != (|$unsigned(reg388)))));
            end
          reg422 <= $unsigned(reg60);
          reg423 = $unsigned({(&wire155[(3'h7):(2'h2)]),
              reg134[(5'h15):(4'h8)]});
        end
    end
  module424 #() modinst1270 (wire1269, clk, reg104, reg398, reg112, reg403, reg111, reg103);
  assign wire1271 = ((~reg178[(5'h13):(4'h9)]) ?
                        $unsigned((&$signed((+wire87)))) : ($unsigned(reg123) - ($signed((reg132 ?
                            reg131 : reg322)) * ($unsigned(wire55) ?
                            (reg327 <<< wire350) : (8'ha9)))));
  assign wire1272 = (+$unsigned((reg85 ?
                        ((reg123 ?
                            reg415 : wire1271) + reg373[(5'h1a):(5'h19)]) : (^~reg405[(3'h4):(1'h0)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module424
#(parameter param1266 = ({(!(((7'h4f) << (8'hbb)) ? ((7'h42) ? (8'hae) : (8'haa)) : ((8'h9d) != (8'ha3)))), {((7'h4d) ? ((8'h9e) ? (7'h56) : (7'h4e)) : ((7'h49) ? (7'h4b) : (8'hb0))), ((8'hbd) ? ((8'h9d) ? (7'h4c) : (8'ha0)) : ((8'ha2) ? (7'h44) : (8'hb0))), ((7'h47) ? ((7'h4e) >= (8'ha8)) : {(7'h4e), (7'h43)})}} >>> (7'h45)), 
parameter param1267 = ({{({param1266} | (param1266 << (8'ha9))), (|(param1266 && param1266)), ((~param1266) | (param1266 == (8'h9c)))}, {(&{(7'h57), (8'hbc)}), (param1266 * (param1266 <= param1266))}} + param1266), 
parameter param1268 = (&((param1266 ? ((~^param1266) & param1266) : (7'h52)) & param1266)))
(y, clk, wire430, wire429, wire428, wire427, wire426, wire425);
  output wire [(32'h37e9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire430;
  input wire signed [(5'h1e):(1'h0)] wire429;
  input wire [(4'h8):(1'h0)] wire428;
  input wire [(2'h3):(1'h0)] wire427;
  input wire [(5'h19):(1'h0)] wire426;
  input wire signed [(2'h2):(1'h0)] wire425;
  wire [(5'h1f):(1'h0)] wire1265;
  wire signed [(5'h1a):(1'h0)] wire1215;
  wire [(4'h9):(1'h0)] wire1089;
  wire [(5'h1f):(1'h0)] wire678;
  wire [(2'h2):(1'h0)] wire670;
  wire [(4'hc):(1'h0)] wire594;
  wire signed [(4'hb):(1'h0)] wire564;
  wire [(5'h18):(1'h0)] wire431;
  reg signed [(2'h2):(1'h0)] reg1261 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1260 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1255 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1254 = (1'h0);
  reg [(5'h17):(1'h0)] reg1253 = (1'h0);
  reg [(5'h13):(1'h0)] reg1252 = (1'h0);
  reg [(5'h15):(1'h0)] reg1251 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1247 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1246 = (1'h0);
  reg [(3'h5):(1'h0)] reg1243 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1239 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1238 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1235 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1231 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1230 = (1'h0);
  reg [(5'h19):(1'h0)] reg1229 = (1'h0);
  reg [(3'h4):(1'h0)] reg1228 = (1'h0);
  reg [(4'h8):(1'h0)] reg1225 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1224 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1222 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1221 = (1'h0);
  reg [(3'h4):(1'h0)] reg1218 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1214 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1213 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1211 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1210 = (1'h0);
  reg [(3'h5):(1'h0)] reg1207 = (1'h0);
  reg [(5'h11):(1'h0)] reg1204 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1200 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1194 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1191 = (1'h0);
  reg [(3'h4):(1'h0)] reg1190 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1187 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1186 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1181 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1180 = (1'h0);
  reg [(5'h14):(1'h0)] reg1179 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1178 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1177 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1175 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1172 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1171 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1169 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1167 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1164 = (1'h0);
  reg [(4'hb):(1'h0)] reg1160 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1159 = (1'h0);
  reg [(5'h10):(1'h0)] reg1155 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1154 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1151 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1150 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1148 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1147 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1146 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1144 = (1'h0);
  reg [(5'h19):(1'h0)] reg1142 = (1'h0);
  reg [(4'hd):(1'h0)] reg1131 = (1'h0);
  reg [(3'h5):(1'h0)] reg1138 = (1'h0);
  reg [(5'h17):(1'h0)] reg1137 = (1'h0);
  reg [(3'h4):(1'h0)] reg1134 = (1'h0);
  reg [(4'hc):(1'h0)] reg1129 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1126 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1123 = (1'h0);
  reg [(4'h9):(1'h0)] reg1120 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1119 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1117 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1114 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1108 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1106 = (1'h0);
  reg [(4'h9):(1'h0)] reg1103 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1102 = (1'h0);
  reg [(3'h5):(1'h0)] reg1100 = (1'h0);
  reg [(4'hd):(1'h0)] reg1099 = (1'h0);
  reg [(4'hb):(1'h0)] reg1097 = (1'h0);
  reg [(5'h13):(1'h0)] reg1096 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1095 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1094 = (1'h0);
  reg [(5'h13):(1'h0)] reg1093 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1088 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1087 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1085 = (1'h0);
  reg [(4'he):(1'h0)] reg1084 = (1'h0);
  reg [(5'h10):(1'h0)] reg1083 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1077 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1076 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1075 = (1'h0);
  reg [(4'hd):(1'h0)] reg1074 = (1'h0);
  reg [(4'hb):(1'h0)] reg1065 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1072 = (1'h0);
  reg [(5'h15):(1'h0)] reg1069 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1067 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1063 = (1'h0);
  reg [(5'h16):(1'h0)] reg1062 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1057 = (1'h0);
  reg [(5'h14):(1'h0)] reg1056 = (1'h0);
  reg [(4'hc):(1'h0)] reg1054 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1053 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1050 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1049 = (1'h0);
  reg [(5'h16):(1'h0)] reg1048 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1047 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1041 = (1'h0);
  reg [(4'hf):(1'h0)] reg1039 = (1'h0);
  reg [(3'h6):(1'h0)] reg1037 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1036 = (1'h0);
  reg [(4'h8):(1'h0)] reg1035 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1029 = (1'h0);
  reg [(4'hb):(1'h0)] reg1032 = (1'h0);
  reg [(3'h6):(1'h0)] reg1027 = (1'h0);
  reg [(2'h3):(1'h0)] reg1025 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1023 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1022 = (1'h0);
  reg [(2'h3):(1'h0)] reg1021 = (1'h0);
  reg [(5'h19):(1'h0)] reg1019 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1018 = (1'h0);
  reg [(5'h13):(1'h0)] reg1016 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1008 = (1'h0);
  reg [(5'h17):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1007 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1005 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1001 = (1'h0);
  reg [(2'h3):(1'h0)] reg996 = (1'h0);
  reg [(5'h12):(1'h0)] reg995 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg992 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg990 = (1'h0);
  reg [(5'h19):(1'h0)] reg989 = (1'h0);
  reg [(5'h14):(1'h0)] reg983 = (1'h0);
  reg [(5'h17):(1'h0)] reg982 = (1'h0);
  reg [(4'hb):(1'h0)] reg979 = (1'h0);
  reg [(3'h6):(1'h0)] reg978 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg974 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg972 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg971 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg966 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg964 = (1'h0);
  reg [(4'hf):(1'h0)] reg963 = (1'h0);
  reg [(5'h12):(1'h0)] reg962 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg960 = (1'h0);
  reg [(5'h1d):(1'h0)] reg958 = (1'h0);
  reg [(4'hb):(1'h0)] reg957 = (1'h0);
  reg [(3'h4):(1'h0)] reg954 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg952 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg949 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg944 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg942 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg940 = (1'h0);
  reg [(5'h1a):(1'h0)] reg935 = (1'h0);
  reg [(4'hc):(1'h0)] reg934 = (1'h0);
  reg [(4'ha):(1'h0)] reg932 = (1'h0);
  reg [(5'h1a):(1'h0)] reg930 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg929 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg928 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg925 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg923 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg921 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg920 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg919 = (1'h0);
  reg [(5'h1a):(1'h0)] reg915 = (1'h0);
  reg signed [(4'he):(1'h0)] reg914 = (1'h0);
  reg [(3'h6):(1'h0)] reg912 = (1'h0);
  reg [(4'hc):(1'h0)] reg911 = (1'h0);
  reg [(5'h15):(1'h0)] reg908 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg899 = (1'h0);
  reg [(4'ha):(1'h0)] reg898 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg897 = (1'h0);
  reg [(4'hf):(1'h0)] reg893 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg892 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg886 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg884 = (1'h0);
  reg [(5'h14):(1'h0)] reg883 = (1'h0);
  reg [(4'hd):(1'h0)] reg882 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg880 = (1'h0);
  reg [(5'h15):(1'h0)] reg879 = (1'h0);
  reg [(5'h13):(1'h0)] reg878 = (1'h0);
  reg signed [(4'he):(1'h0)] reg871 = (1'h0);
  reg [(5'h17):(1'h0)] reg875 = (1'h0);
  reg [(5'h1d):(1'h0)] reg872 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg866 = (1'h0);
  reg [(5'h15):(1'h0)] reg861 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg858 = (1'h0);
  reg [(4'hf):(1'h0)] reg857 = (1'h0);
  reg [(5'h12):(1'h0)] reg853 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg849 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg845 = (1'h0);
  reg [(4'hd):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg834 = (1'h0);
  reg signed [(4'he):(1'h0)] reg832 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg831 = (1'h0);
  reg [(3'h4):(1'h0)] reg827 = (1'h0);
  reg [(5'h18):(1'h0)] reg824 = (1'h0);
  reg [(5'h13):(1'h0)] reg822 = (1'h0);
  reg [(3'h7):(1'h0)] reg820 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg816 = (1'h0);
  reg [(4'hf):(1'h0)] reg814 = (1'h0);
  reg [(4'h9):(1'h0)] reg813 = (1'h0);
  reg [(5'h1e):(1'h0)] reg809 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg808 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg806 = (1'h0);
  reg [(3'h6):(1'h0)] reg805 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg804 = (1'h0);
  reg [(5'h1d):(1'h0)] reg797 = (1'h0);
  reg [(3'h7):(1'h0)] reg796 = (1'h0);
  reg [(2'h2):(1'h0)] reg791 = (1'h0);
  reg [(3'h6):(1'h0)] reg789 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg788 = (1'h0);
  reg [(3'h7):(1'h0)] reg787 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg783 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg782 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg780 = (1'h0);
  reg [(3'h5):(1'h0)] reg777 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg776 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg771 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg768 = (1'h0);
  reg [(2'h2):(1'h0)] reg766 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg760 = (1'h0);
  reg [(3'h4):(1'h0)] reg755 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg753 = (1'h0);
  reg [(3'h5):(1'h0)] reg750 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg748 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg747 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg746 = (1'h0);
  reg [(5'h11):(1'h0)] reg743 = (1'h0);
  reg [(5'h18):(1'h0)] reg742 = (1'h0);
  reg [(3'h7):(1'h0)] reg740 = (1'h0);
  reg [(5'h13):(1'h0)] reg735 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg734 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg732 = (1'h0);
  reg [(5'h1a):(1'h0)] reg730 = (1'h0);
  reg [(5'h1d):(1'h0)] reg728 = (1'h0);
  reg [(4'hf):(1'h0)] reg727 = (1'h0);
  reg [(5'h19):(1'h0)] reg726 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg723 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg721 = (1'h0);
  reg [(3'h7):(1'h0)] reg719 = (1'h0);
  reg [(5'h1e):(1'h0)] reg717 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg714 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg712 = (1'h0);
  reg [(5'h17):(1'h0)] reg709 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg707 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg706 = (1'h0);
  reg [(5'h1d):(1'h0)] reg703 = (1'h0);
  reg [(5'h13):(1'h0)] reg702 = (1'h0);
  reg [(3'h4):(1'h0)] reg700 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg699 = (1'h0);
  reg [(5'h1b):(1'h0)] reg698 = (1'h0);
  reg [(4'hb):(1'h0)] reg695 = (1'h0);
  reg [(2'h2):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg691 = (1'h0);
  reg [(2'h3):(1'h0)] reg690 = (1'h0);
  reg [(4'ha):(1'h0)] reg688 = (1'h0);
  reg [(5'h13):(1'h0)] reg684 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg682 = (1'h0);
  reg [(5'h1d):(1'h0)] reg676 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg675 = (1'h0);
  reg [(5'h1c):(1'h0)] reg672 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg667 = (1'h0);
  reg [(4'he):(1'h0)] reg666 = (1'h0);
  reg [(5'h15):(1'h0)] reg664 = (1'h0);
  reg [(4'hc):(1'h0)] reg662 = (1'h0);
  reg [(5'h17):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg655 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg654 = (1'h0);
  reg [(5'h1a):(1'h0)] reg651 = (1'h0);
  reg [(5'h10):(1'h0)] reg650 = (1'h0);
  reg [(4'ha):(1'h0)] reg649 = (1'h0);
  reg signed [(4'he):(1'h0)] reg646 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg640 = (1'h0);
  reg [(2'h2):(1'h0)] reg639 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg635 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg628 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg625 = (1'h0);
  reg [(4'hd):(1'h0)] reg620 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg616 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg615 = (1'h0);
  reg [(4'hd):(1'h0)] reg613 = (1'h0);
  reg [(3'h5):(1'h0)] reg611 = (1'h0);
  reg [(3'h6):(1'h0)] reg607 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg606 = (1'h0);
  reg [(4'he):(1'h0)] reg605 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg604 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg603 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg599 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg598 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg596 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg592 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg589 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg586 = (1'h0);
  reg [(4'he):(1'h0)] reg585 = (1'h0);
  reg [(5'h14):(1'h0)] reg579 = (1'h0);
  reg [(3'h6):(1'h0)] reg575 = (1'h0);
  reg [(5'h12):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg572 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg571 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg569 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg566 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg561 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg558 = (1'h0);
  reg [(4'he):(1'h0)] reg552 = (1'h0);
  reg [(5'h13):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg549 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg546 = (1'h0);
  reg [(5'h13):(1'h0)] reg543 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg542 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg539 = (1'h0);
  reg [(5'h19):(1'h0)] reg537 = (1'h0);
  reg [(5'h15):(1'h0)] reg530 = (1'h0);
  reg signed [(4'he):(1'h0)] reg529 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg528 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg525 = (1'h0);
  reg [(5'h11):(1'h0)] reg522 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg520 = (1'h0);
  reg [(5'h1d):(1'h0)] reg519 = (1'h0);
  reg [(5'h19):(1'h0)] reg516 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg515 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg514 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg512 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg511 = (1'h0);
  reg [(5'h15):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg506 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg503 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg500 = (1'h0);
  reg [(4'hf):(1'h0)] reg498 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg497 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg495 = (1'h0);
  reg [(5'h16):(1'h0)] reg493 = (1'h0);
  reg [(2'h3):(1'h0)] reg490 = (1'h0);
  reg [(5'h13):(1'h0)] reg489 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg486 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg485 = (1'h0);
  reg signed [(4'he):(1'h0)] reg484 = (1'h0);
  reg [(4'h8):(1'h0)] reg482 = (1'h0);
  reg [(5'h1f):(1'h0)] reg469 = (1'h0);
  reg [(5'h14):(1'h0)] reg467 = (1'h0);
  reg [(4'hc):(1'h0)] reg466 = (1'h0);
  reg [(5'h1b):(1'h0)] reg463 = (1'h0);
  reg [(5'h17):(1'h0)] reg460 = (1'h0);
  reg [(4'he):(1'h0)] reg458 = (1'h0);
  reg [(5'h12):(1'h0)] reg457 = (1'h0);
  reg [(3'h6):(1'h0)] reg456 = (1'h0);
  reg [(5'h12):(1'h0)] reg455 = (1'h0);
  reg [(4'h8):(1'h0)] reg454 = (1'h0);
  reg [(4'hc):(1'h0)] reg452 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg450 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg447 = (1'h0);
  reg [(5'h1a):(1'h0)] reg443 = (1'h0);
  reg [(4'ha):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg439 = (1'h0);
  reg [(3'h4):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg434 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg433 = (1'h0);
  reg [(5'h15):(1'h0)] reg1264 = (1'h0);
  reg [(5'h14):(1'h0)] reg1263 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1262 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1259 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1258 = (1'h0);
  reg [(4'hc):(1'h0)] reg1257 = (1'h0);
  reg [(5'h11):(1'h0)] reg1256 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1250 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1249 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1248 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1245 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1244 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1242 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1241 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1240 = (1'h0);
  reg [(3'h5):(1'h0)] reg1237 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1236 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1234 = (1'h0);
  reg [(4'ha):(1'h0)] reg1233 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1232 = (1'h0);
  reg [(4'hc):(1'h0)] reg1227 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1226 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1223 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1220 = (1'h0);
  reg [(5'h18):(1'h0)] reg1219 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1217 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1216 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1212 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1209 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1208 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1206 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1205 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1203 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1202 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1201 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1199 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1198 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1197 = (1'h0);
  reg [(5'h15):(1'h0)] reg1196 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1195 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1193 = (1'h0);
  reg [(5'h16):(1'h0)] reg1192 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1189 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1188 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar1179 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1185 = (1'h0);
  reg [(3'h5):(1'h0)] reg1184 = (1'h0);
  reg [(5'h13):(1'h0)] reg1183 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1182 = (1'h0);
  reg [(4'h9):(1'h0)] reg1174 = (1'h0);
  reg [(4'h9):(1'h0)] reg1173 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar1170 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1170 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1168 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1166 = (1'h0);
  reg [(4'h9):(1'h0)] reg1165 = (1'h0);
  reg [(5'h19):(1'h0)] reg1163 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1162 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1161 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1158 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1157 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1156 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1153 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1152 = (1'h0);
  reg [(5'h19):(1'h0)] reg1149 = (1'h0);
  reg [(5'h11):(1'h0)] reg1145 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1143 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1141 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1140 = (1'h0);
  reg [(4'hd):(1'h0)] reg1139 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1130 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1136 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1135 = (1'h0);
  reg [(5'h15):(1'h0)] reg1133 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1132 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1131 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1130 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1128 = (1'h0);
  reg [(4'hf):(1'h0)] reg1127 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1125 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1124 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1122 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1121 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1118 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1116 = (1'h0);
  reg [(5'h14):(1'h0)] reg1115 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1112 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1111 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1110 = (1'h0);
  reg [(5'h15):(1'h0)] reg1109 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1107 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1105 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1104 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1101 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1098 = (1'h0);
  reg [(3'h7):(1'h0)] reg1092 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1091 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1090 = (1'h0);
  reg [(4'he):(1'h0)] reg1086 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1082 = (1'h0);
  reg [(5'h16):(1'h0)] reg1081 = (1'h0);
  reg [(4'hb):(1'h0)] reg1080 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1079 = (1'h0);
  reg [(5'h16):(1'h0)] reg1078 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1073 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1061 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1060 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1058 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1057 = (1'h0);
  reg [(4'h8):(1'h0)] reg1071 = (1'h0);
  reg [(5'h12):(1'h0)] reg1070 = (1'h0);
  reg [(2'h3):(1'h0)] reg1068 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1066 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1065 = (1'h0);
  reg [(5'h13):(1'h0)] reg1064 = (1'h0);
  reg [(4'he):(1'h0)] forvar1061 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1060 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1059 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1058 = (1'h0);
  reg [(5'h12):(1'h0)] reg1055 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1052 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1051 = (1'h0);
  reg [(5'h14):(1'h0)] reg1046 = (1'h0);
  reg [(4'hc):(1'h0)] reg1045 = (1'h0);
  reg [(5'h15):(1'h0)] reg1044 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1043 = (1'h0);
  reg [(5'h18):(1'h0)] reg1042 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1040 = (1'h0);
  reg [(4'hd):(1'h0)] reg1038 = (1'h0);
  reg [(5'h17):(1'h0)] reg1034 = (1'h0);
  reg [(5'h10):(1'h0)] reg1033 = (1'h0);
  reg [(5'h18):(1'h0)] reg1031 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1030 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1029 = (1'h0);
  reg [(4'hd):(1'h0)] reg1028 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1026 = (1'h0);
  reg [(3'h5):(1'h0)] reg1024 = (1'h0);
  reg [(4'hf):(1'h0)] reg1020 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1017 = (1'h0);
  reg [(4'h8):(1'h0)] reg1015 = (1'h0);
  reg [(4'h8):(1'h0)] reg1014 = (1'h0);
  reg [(3'h5):(1'h0)] reg1013 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1011 = (1'h0);
  reg [(4'h9):(1'h0)] reg1010 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1009 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1008 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1006 = (1'h0);
  reg [(4'hd):(1'h0)] reg1004 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1003 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1002 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1000 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg999 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg998 = (1'h0);
  reg [(4'hd):(1'h0)] forvar989 = (1'h0);
  reg [(5'h1a):(1'h0)] reg997 = (1'h0);
  reg [(3'h7):(1'h0)] reg994 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg993 = (1'h0);
  reg signed [(4'he):(1'h0)] reg991 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg988 = (1'h0);
  reg [(3'h6):(1'h0)] forvar987 = (1'h0);
  reg [(2'h2):(1'h0)] reg986 = (1'h0);
  reg [(4'h8):(1'h0)] forvar985 = (1'h0);
  reg [(5'h1e):(1'h0)] reg984 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg981 = (1'h0);
  reg [(5'h1a):(1'h0)] reg980 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg977 = (1'h0);
  reg [(5'h15):(1'h0)] reg976 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg975 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg973 = (1'h0);
  reg [(4'hc):(1'h0)] reg970 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg969 = (1'h0);
  reg [(2'h3):(1'h0)] reg968 = (1'h0);
  reg [(5'h17):(1'h0)] forvar967 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg965 = (1'h0);
  reg [(4'h8):(1'h0)] reg961 = (1'h0);
  reg [(5'h18):(1'h0)] reg959 = (1'h0);
  reg [(4'hf):(1'h0)] forvar956 = (1'h0);
  reg [(3'h7):(1'h0)] reg955 = (1'h0);
  reg [(4'ha):(1'h0)] reg953 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg951 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg950 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar948 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar947 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg946 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg945 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg943 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg941 = (1'h0);
  reg [(4'h9):(1'h0)] reg939 = (1'h0);
  reg [(5'h12):(1'h0)] reg938 = (1'h0);
  reg [(5'h1e):(1'h0)] reg937 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg936 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar933 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg931 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar925 = (1'h0);
  reg [(5'h16):(1'h0)] reg922 = (1'h0);
  reg [(4'hc):(1'h0)] reg927 = (1'h0);
  reg [(5'h11):(1'h0)] reg926 = (1'h0);
  reg [(5'h11):(1'h0)] reg924 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar922 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg918 = (1'h0);
  reg [(5'h12):(1'h0)] forvar911 = (1'h0);
  reg [(5'h1d):(1'h0)] reg917 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg916 = (1'h0);
  reg [(4'h8):(1'h0)] reg913 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg910 = (1'h0);
  reg [(4'hb):(1'h0)] reg909 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg900 = (1'h0);
  reg [(5'h1b):(1'h0)] reg907 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg906 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg905 = (1'h0);
  reg [(4'hd):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg902 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg901 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar900 = (1'h0);
  reg [(4'hf):(1'h0)] reg896 = (1'h0);
  reg [(4'hf):(1'h0)] reg895 = (1'h0);
  reg [(5'h11):(1'h0)] reg894 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg891 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg890 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg889 = (1'h0);
  reg signed [(4'he):(1'h0)] reg888 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar887 = (1'h0);
  reg [(5'h1d):(1'h0)] reg885 = (1'h0);
  reg [(2'h2):(1'h0)] forvar881 = (1'h0);
  reg [(4'hb):(1'h0)] forvar872 = (1'h0);
  reg [(4'hd):(1'h0)] reg877 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg876 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg874 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg873 = (1'h0);
  reg [(5'h12):(1'h0)] forvar871 = (1'h0);
  reg [(5'h19):(1'h0)] reg870 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg869 = (1'h0);
  reg [(5'h1f):(1'h0)] reg867 = (1'h0);
  reg [(4'he):(1'h0)] reg865 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg864 = (1'h0);
  reg [(5'h1c):(1'h0)] reg863 = (1'h0);
  reg [(5'h12):(1'h0)] reg862 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg860 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg859 = (1'h0);
  reg [(4'h9):(1'h0)] reg856 = (1'h0);
  reg [(5'h14):(1'h0)] reg855 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg854 = (1'h0);
  reg [(5'h1e):(1'h0)] reg852 = (1'h0);
  reg [(3'h4):(1'h0)] reg851 = (1'h0);
  reg [(4'he):(1'h0)] reg850 = (1'h0);
  reg [(5'h16):(1'h0)] reg848 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar847 = (1'h0);
  reg [(4'ha):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg837 = (1'h0);
  reg [(3'h7):(1'h0)] forvar836 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg844 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg843 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg842 = (1'h0);
  reg [(5'h19):(1'h0)] reg841 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar840 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg839 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg838 = (1'h0);
  reg [(5'h18):(1'h0)] forvar837 = (1'h0);
  reg [(4'h8):(1'h0)] reg836 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg835 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg833 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar830 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg829 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg828 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg826 = (1'h0);
  reg [(4'hd):(1'h0)] reg825 = (1'h0);
  reg [(4'hc):(1'h0)] forvar823 = (1'h0);
  reg [(2'h3):(1'h0)] reg821 = (1'h0);
  reg [(2'h2):(1'h0)] reg818 = (1'h0);
  reg [(4'h8):(1'h0)] reg817 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg815 = (1'h0);
  reg [(5'h1c):(1'h0)] reg812 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg811 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar810 = (1'h0);
  reg [(5'h1e):(1'h0)] reg807 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg803 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar802 = (1'h0);
  reg [(3'h7):(1'h0)] reg801 = (1'h0);
  reg [(5'h16):(1'h0)] reg800 = (1'h0);
  reg [(5'h1b):(1'h0)] reg799 = (1'h0);
  reg [(4'he):(1'h0)] forvar798 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg795 = (1'h0);
  reg [(5'h11):(1'h0)] forvar794 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg793 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar792 = (1'h0);
  reg [(5'h13):(1'h0)] reg790 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar786 = (1'h0);
  reg [(5'h18):(1'h0)] reg785 = (1'h0);
  reg [(5'h12):(1'h0)] reg784 = (1'h0);
  reg [(5'h19):(1'h0)] forvar781 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar779 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg778 = (1'h0);
  reg [(4'h9):(1'h0)] reg775 = (1'h0);
  reg [(4'h9):(1'h0)] reg774 = (1'h0);
  reg [(4'hf):(1'h0)] reg773 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar772 = (1'h0);
  reg [(5'h16):(1'h0)] reg770 = (1'h0);
  reg [(5'h1d):(1'h0)] reg769 = (1'h0);
  reg [(3'h7):(1'h0)] reg767 = (1'h0);
  reg [(3'h6):(1'h0)] reg765 = (1'h0);
  reg [(5'h19):(1'h0)] forvar764 = (1'h0);
  reg [(5'h14):(1'h0)] reg763 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg762 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg761 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg758 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar757 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar756 = (1'h0);
  reg [(5'h14):(1'h0)] reg754 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg752 = (1'h0);
  reg [(5'h18):(1'h0)] reg751 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg749 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg744 = (1'h0);
  reg [(4'hd):(1'h0)] reg729 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg745 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar744 = (1'h0);
  reg [(5'h15):(1'h0)] reg741 = (1'h0);
  reg [(3'h4):(1'h0)] reg739 = (1'h0);
  reg [(5'h16):(1'h0)] reg738 = (1'h0);
  reg [(4'hc):(1'h0)] reg737 = (1'h0);
  reg [(3'h7):(1'h0)] reg736 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg733 = (1'h0);
  reg [(4'hf):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar729 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg725 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar722 = (1'h0);
  reg [(5'h1d):(1'h0)] reg720 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar718 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar713 = (1'h0);
  reg [(5'h18):(1'h0)] reg711 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar710 = (1'h0);
  reg [(3'h4):(1'h0)] reg708 = (1'h0);
  reg [(5'h1d):(1'h0)] reg705 = (1'h0);
  reg [(5'h17):(1'h0)] reg704 = (1'h0);
  reg [(5'h16):(1'h0)] forvar701 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg697 = (1'h0);
  reg [(5'h13):(1'h0)] reg696 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg694 = (1'h0);
  reg [(5'h15):(1'h0)] reg692 = (1'h0);
  reg [(4'h9):(1'h0)] reg689 = (1'h0);
  reg [(5'h17):(1'h0)] reg687 = (1'h0);
  reg [(2'h2):(1'h0)] reg686 = (1'h0);
  reg [(5'h15):(1'h0)] reg685 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg680 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar679 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg683 = (1'h0);
  reg [(5'h1f):(1'h0)] reg681 = (1'h0);
  reg [(5'h14):(1'h0)] forvar680 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg679 = (1'h0);
  reg [(4'hb):(1'h0)] reg677 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar674 = (1'h0);
  reg [(5'h14):(1'h0)] reg673 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar671 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg669 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg663 = (1'h0);
  reg [(5'h11):(1'h0)] reg660 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar659 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar658 = (1'h0);
  reg [(4'ha):(1'h0)] reg657 = (1'h0);
  reg signed [(4'he):(1'h0)] reg656 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar653 = (1'h0);
  reg [(4'h8):(1'h0)] reg652 = (1'h0);
  reg [(3'h4):(1'h0)] reg648 = (1'h0);
  reg [(2'h3):(1'h0)] reg647 = (1'h0);
  reg [(3'h6):(1'h0)] reg644 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg643 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg642 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg641 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg638 = (1'h0);
  reg [(5'h13):(1'h0)] reg637 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg636 = (1'h0);
  reg [(4'hd):(1'h0)] reg634 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar633 = (1'h0);
  reg [(3'h4):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar631 = (1'h0);
  reg [(3'h6):(1'h0)] reg630 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg629 = (1'h0);
  reg [(3'h5):(1'h0)] reg627 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg626 = (1'h0);
  reg [(5'h1e):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg622 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar621 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar619 = (1'h0);
  reg [(5'h13):(1'h0)] reg618 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg617 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg614 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg612 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg610 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg609 = (1'h0);
  reg [(5'h1c):(1'h0)] reg608 = (1'h0);
  reg [(5'h16):(1'h0)] reg602 = (1'h0);
  reg [(5'h19):(1'h0)] forvar601 = (1'h0);
  reg [(5'h17):(1'h0)] reg600 = (1'h0);
  reg [(5'h12):(1'h0)] reg597 = (1'h0);
  reg [(4'h9):(1'h0)] forvar595 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg593 = (1'h0);
  reg [(3'h7):(1'h0)] forvar591 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg590 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg588 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg587 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar584 = (1'h0);
  reg [(5'h1f):(1'h0)] reg583 = (1'h0);
  reg [(4'hd):(1'h0)] reg582 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg581 = (1'h0);
  reg [(5'h1e):(1'h0)] reg580 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg578 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar577 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar576 = (1'h0);
  reg [(5'h10):(1'h0)] reg574 = (1'h0);
  reg [(5'h16):(1'h0)] reg570 = (1'h0);
  reg [(5'h1c):(1'h0)] reg568 = (1'h0);
  reg [(4'h8):(1'h0)] reg567 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar565 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg563 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg560 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg559 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar557 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg556 = (1'h0);
  reg [(4'hb):(1'h0)] forvar555 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar554 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg553 = (1'h0);
  reg [(5'h13):(1'h0)] reg550 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar548 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar547 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg545 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar541 = (1'h0);
  reg [(5'h1a):(1'h0)] reg540 = (1'h0);
  reg [(5'h1a):(1'h0)] reg538 = (1'h0);
  reg [(4'hb):(1'h0)] reg536 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg535 = (1'h0);
  reg [(5'h11):(1'h0)] reg534 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg533 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg531 = (1'h0);
  reg [(5'h1b):(1'h0)] reg521 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar502 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg527 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg524 = (1'h0);
  reg [(5'h19):(1'h0)] reg523 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar521 = (1'h0);
  reg [(3'h6):(1'h0)] reg518 = (1'h0);
  reg [(4'hc):(1'h0)] reg517 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg513 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg509 = (1'h0);
  reg [(5'h12):(1'h0)] reg508 = (1'h0);
  reg [(5'h10):(1'h0)] reg507 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg505 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg502 = (1'h0);
  reg [(5'h12):(1'h0)] reg501 = (1'h0);
  reg [(5'h11):(1'h0)] reg499 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg496 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar487 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg494 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg491 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg488 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg487 = (1'h0);
  reg [(5'h1a):(1'h0)] reg483 = (1'h0);
  reg [(5'h1a):(1'h0)] reg481 = (1'h0);
  reg [(5'h1b):(1'h0)] reg480 = (1'h0);
  reg [(3'h7):(1'h0)] reg479 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg477 = (1'h0);
  reg [(5'h14):(1'h0)] reg476 = (1'h0);
  reg [(5'h10):(1'h0)] reg475 = (1'h0);
  reg [(3'h6):(1'h0)] forvar474 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar473 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg472 = (1'h0);
  reg [(5'h1c):(1'h0)] reg471 = (1'h0);
  reg [(4'h9):(1'h0)] reg470 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg468 = (1'h0);
  reg [(5'h1a):(1'h0)] reg465 = (1'h0);
  reg [(5'h1e):(1'h0)] reg464 = (1'h0);
  reg [(5'h17):(1'h0)] reg462 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg461 = (1'h0);
  reg [(5'h13):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar451 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg449 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg446 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg445 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar444 = (1'h0);
  reg [(5'h1a):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg440 = (1'h0);
  reg [(3'h6):(1'h0)] forvar437 = (1'h0);
  reg [(5'h15):(1'h0)] reg436 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg435 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg432 = (1'h0);
  assign y = {wire1265,
                 wire1215,
                 wire1089,
                 wire678,
                 wire670,
                 wire594,
                 wire564,
                 wire431,
                 reg1261,
                 reg1260,
                 reg1255,
                 reg1254,
                 reg1253,
                 reg1252,
                 reg1251,
                 reg1247,
                 reg1246,
                 reg1243,
                 reg1239,
                 reg1238,
                 reg1235,
                 reg1231,
                 reg1230,
                 reg1229,
                 reg1228,
                 reg1225,
                 reg1224,
                 reg1222,
                 reg1221,
                 reg1218,
                 reg1214,
                 reg1213,
                 reg1211,
                 reg1210,
                 reg1207,
                 reg1204,
                 reg1200,
                 reg1194,
                 reg1191,
                 reg1190,
                 reg1187,
                 reg1186,
                 reg1181,
                 reg1180,
                 reg1179,
                 reg1178,
                 reg1177,
                 reg1176,
                 reg1175,
                 reg1172,
                 reg1171,
                 reg1169,
                 reg1167,
                 reg1164,
                 reg1160,
                 reg1159,
                 reg1155,
                 reg1154,
                 reg1151,
                 reg1150,
                 reg1148,
                 reg1147,
                 reg1146,
                 reg1144,
                 reg1142,
                 reg1131,
                 reg1138,
                 reg1137,
                 reg1134,
                 reg1129,
                 reg1126,
                 reg1123,
                 reg1120,
                 reg1119,
                 reg1117,
                 reg1114,
                 reg1113,
                 reg1108,
                 reg1106,
                 reg1103,
                 reg1102,
                 reg1100,
                 reg1099,
                 reg1097,
                 reg1096,
                 reg1095,
                 reg1094,
                 reg1093,
                 reg1088,
                 reg1087,
                 reg1085,
                 reg1084,
                 reg1083,
                 reg1077,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1065,
                 reg1072,
                 reg1069,
                 reg1067,
                 reg1063,
                 reg1062,
                 reg1057,
                 reg1056,
                 reg1054,
                 reg1053,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1047,
                 reg1041,
                 reg1039,
                 reg1037,
                 reg1036,
                 reg1035,
                 reg1029,
                 reg1032,
                 reg1027,
                 reg1025,
                 reg1023,
                 reg1022,
                 reg1021,
                 reg1019,
                 reg1018,
                 reg1016,
                 reg1008,
                 reg1012,
                 reg1007,
                 reg1005,
                 reg1001,
                 reg996,
                 reg995,
                 reg992,
                 reg990,
                 reg989,
                 reg983,
                 reg982,
                 reg979,
                 reg978,
                 reg974,
                 reg972,
                 reg971,
                 reg966,
                 reg964,
                 reg963,
                 reg962,
                 reg960,
                 reg958,
                 reg957,
                 reg954,
                 reg952,
                 reg949,
                 reg944,
                 reg942,
                 reg940,
                 reg935,
                 reg934,
                 reg932,
                 reg930,
                 reg929,
                 reg928,
                 reg925,
                 reg923,
                 reg921,
                 reg920,
                 reg919,
                 reg915,
                 reg914,
                 reg912,
                 reg911,
                 reg908,
                 reg903,
                 reg899,
                 reg898,
                 reg897,
                 reg893,
                 reg892,
                 reg886,
                 reg884,
                 reg883,
                 reg882,
                 reg880,
                 reg879,
                 reg878,
                 reg871,
                 reg875,
                 reg872,
                 reg868,
                 reg866,
                 reg861,
                 reg858,
                 reg857,
                 reg853,
                 reg849,
                 reg845,
                 reg840,
                 reg834,
                 reg832,
                 reg831,
                 reg827,
                 reg824,
                 reg822,
                 reg820,
                 reg819,
                 reg816,
                 reg814,
                 reg813,
                 reg809,
                 reg808,
                 reg806,
                 reg805,
                 reg804,
                 reg797,
                 reg796,
                 reg791,
                 reg789,
                 reg788,
                 reg787,
                 reg783,
                 reg782,
                 reg780,
                 reg777,
                 reg776,
                 reg771,
                 reg768,
                 reg766,
                 reg760,
                 reg755,
                 reg753,
                 reg750,
                 reg748,
                 reg747,
                 reg746,
                 reg743,
                 reg742,
                 reg740,
                 reg735,
                 reg734,
                 reg732,
                 reg730,
                 reg728,
                 reg727,
                 reg726,
                 reg723,
                 reg721,
                 reg719,
                 reg717,
                 reg714,
                 reg712,
                 reg709,
                 reg707,
                 reg706,
                 reg703,
                 reg702,
                 reg700,
                 reg699,
                 reg698,
                 reg695,
                 reg693,
                 reg691,
                 reg690,
                 reg688,
                 reg684,
                 reg682,
                 reg676,
                 reg675,
                 reg672,
                 reg667,
                 reg666,
                 reg664,
                 reg662,
                 reg661,
                 reg655,
                 reg654,
                 reg651,
                 reg650,
                 reg649,
                 reg646,
                 reg645,
                 reg640,
                 reg639,
                 reg635,
                 reg628,
                 reg625,
                 reg620,
                 reg616,
                 reg615,
                 reg613,
                 reg611,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg599,
                 reg598,
                 reg596,
                 reg592,
                 reg589,
                 reg586,
                 reg585,
                 reg579,
                 reg575,
                 reg573,
                 reg572,
                 reg571,
                 reg569,
                 reg566,
                 reg562,
                 reg561,
                 reg558,
                 reg552,
                 reg551,
                 reg549,
                 reg546,
                 reg543,
                 reg542,
                 reg539,
                 reg537,
                 reg530,
                 reg529,
                 reg528,
                 reg525,
                 reg522,
                 reg520,
                 reg519,
                 reg516,
                 reg515,
                 reg514,
                 reg512,
                 reg511,
                 reg510,
                 reg506,
                 reg503,
                 reg500,
                 reg498,
                 reg497,
                 reg495,
                 reg493,
                 reg490,
                 reg489,
                 reg486,
                 reg485,
                 reg484,
                 reg482,
                 reg469,
                 reg467,
                 reg466,
                 reg463,
                 reg460,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg452,
                 reg450,
                 reg447,
                 reg443,
                 reg442,
                 reg439,
                 reg438,
                 reg437,
                 reg434,
                 reg433,
                 reg1264,
                 reg1263,
                 reg1262,
                 reg1259,
                 reg1258,
                 reg1257,
                 reg1256,
                 reg1250,
                 reg1249,
                 reg1248,
                 reg1245,
                 reg1244,
                 reg1242,
                 reg1241,
                 forvar1240,
                 reg1237,
                 reg1236,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1227,
                 reg1226,
                 reg1223,
                 reg1220,
                 reg1219,
                 forvar1217,
                 forvar1216,
                 reg1212,
                 reg1209,
                 reg1208,
                 forvar1206,
                 reg1205,
                 reg1203,
                 reg1202,
                 forvar1201,
                 forvar1199,
                 reg1198,
                 forvar1197,
                 reg1196,
                 reg1195,
                 reg1193,
                 reg1192,
                 forvar1189,
                 reg1188,
                 forvar1179,
                 reg1185,
                 reg1184,
                 reg1183,
                 reg1182,
                 reg1174,
                 reg1173,
                 forvar1170,
                 reg1170,
                 reg1168,
                 reg1166,
                 reg1165,
                 reg1163,
                 reg1162,
                 forvar1161,
                 reg1158,
                 reg1157,
                 reg1156,
                 reg1153,
                 forvar1152,
                 reg1149,
                 reg1145,
                 reg1143,
                 reg1141,
                 reg1140,
                 reg1139,
                 forvar1130,
                 reg1136,
                 reg1135,
                 reg1133,
                 reg1132,
                 forvar1131,
                 reg1130,
                 reg1128,
                 reg1127,
                 reg1125,
                 reg1124,
                 reg1122,
                 reg1121,
                 reg1118,
                 reg1116,
                 reg1115,
                 reg1112,
                 reg1111,
                 reg1110,
                 reg1109,
                 reg1107,
                 reg1105,
                 forvar1104,
                 reg1101,
                 reg1098,
                 reg1092,
                 forvar1091,
                 forvar1090,
                 reg1086,
                 reg1082,
                 reg1081,
                 reg1080,
                 forvar1079,
                 reg1078,
                 reg1073,
                 reg1061,
                 forvar1060,
                 reg1058,
                 forvar1057,
                 reg1071,
                 reg1070,
                 reg1068,
                 reg1066,
                 forvar1065,
                 reg1064,
                 forvar1061,
                 reg1060,
                 reg1059,
                 forvar1058,
                 reg1055,
                 reg1052,
                 reg1051,
                 reg1046,
                 reg1045,
                 reg1044,
                 reg1043,
                 reg1042,
                 reg1040,
                 reg1038,
                 reg1034,
                 reg1033,
                 reg1031,
                 reg1030,
                 forvar1029,
                 reg1028,
                 forvar1026,
                 reg1024,
                 reg1020,
                 forvar1017,
                 reg1015,
                 reg1014,
                 reg1013,
                 reg1011,
                 reg1010,
                 reg1009,
                 forvar1008,
                 forvar1006,
                 reg1004,
                 reg1003,
                 reg1002,
                 reg1000,
                 reg999,
                 reg998,
                 forvar989,
                 reg997,
                 reg994,
                 reg993,
                 reg991,
                 reg988,
                 forvar987,
                 reg986,
                 forvar985,
                 reg984,
                 reg981,
                 reg980,
                 reg977,
                 reg976,
                 reg975,
                 reg973,
                 reg970,
                 reg969,
                 reg968,
                 forvar967,
                 reg965,
                 reg961,
                 reg959,
                 forvar956,
                 reg955,
                 reg953,
                 reg951,
                 reg950,
                 forvar948,
                 forvar947,
                 reg946,
                 reg945,
                 reg943,
                 reg941,
                 reg939,
                 reg938,
                 reg937,
                 reg936,
                 forvar933,
                 reg931,
                 forvar925,
                 reg922,
                 reg927,
                 reg926,
                 reg924,
                 forvar922,
                 reg918,
                 forvar911,
                 reg917,
                 reg916,
                 reg913,
                 reg910,
                 reg909,
                 reg900,
                 reg907,
                 reg906,
                 reg905,
                 reg904,
                 reg902,
                 reg901,
                 forvar900,
                 reg896,
                 reg895,
                 reg894,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 forvar887,
                 reg885,
                 forvar881,
                 forvar872,
                 reg877,
                 reg876,
                 reg874,
                 reg873,
                 forvar871,
                 reg870,
                 reg869,
                 reg867,
                 reg865,
                 reg864,
                 reg863,
                 reg862,
                 reg860,
                 reg859,
                 reg856,
                 reg855,
                 reg854,
                 reg852,
                 reg851,
                 reg850,
                 reg848,
                 forvar847,
                 reg846,
                 reg837,
                 forvar836,
                 reg844,
                 reg843,
                 reg842,
                 reg841,
                 forvar840,
                 reg839,
                 reg838,
                 forvar837,
                 reg836,
                 reg835,
                 reg833,
                 forvar830,
                 reg829,
                 reg828,
                 reg826,
                 reg825,
                 forvar823,
                 reg821,
                 reg818,
                 reg817,
                 reg815,
                 reg812,
                 reg811,
                 forvar810,
                 reg807,
                 reg803,
                 forvar802,
                 reg801,
                 reg800,
                 reg799,
                 forvar798,
                 reg795,
                 forvar794,
                 reg793,
                 forvar792,
                 reg790,
                 forvar786,
                 reg785,
                 reg784,
                 forvar781,
                 forvar779,
                 reg778,
                 reg775,
                 reg774,
                 reg773,
                 forvar772,
                 reg770,
                 reg769,
                 reg767,
                 reg765,
                 forvar764,
                 reg763,
                 reg762,
                 reg761,
                 reg759,
                 reg758,
                 forvar757,
                 forvar756,
                 reg754,
                 reg752,
                 reg751,
                 reg749,
                 reg744,
                 reg729,
                 reg745,
                 forvar744,
                 reg741,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg733,
                 reg731,
                 forvar729,
                 reg725,
                 reg724,
                 forvar722,
                 reg720,
                 forvar718,
                 reg716,
                 reg715,
                 forvar713,
                 reg711,
                 forvar710,
                 reg708,
                 reg705,
                 reg704,
                 forvar701,
                 reg697,
                 reg696,
                 reg694,
                 reg692,
                 reg689,
                 reg687,
                 reg686,
                 reg685,
                 reg680,
                 forvar679,
                 reg683,
                 reg681,
                 forvar680,
                 reg679,
                 reg677,
                 forvar674,
                 reg673,
                 forvar671,
                 reg669,
                 reg668,
                 reg665,
                 reg663,
                 reg660,
                 forvar659,
                 forvar658,
                 reg657,
                 reg656,
                 forvar653,
                 reg652,
                 reg648,
                 reg647,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg638,
                 reg637,
                 reg636,
                 reg634,
                 forvar633,
                 reg632,
                 forvar631,
                 reg630,
                 reg629,
                 reg627,
                 reg626,
                 reg624,
                 reg623,
                 reg622,
                 forvar621,
                 forvar619,
                 reg618,
                 reg617,
                 reg614,
                 reg612,
                 reg610,
                 reg609,
                 reg608,
                 reg602,
                 forvar601,
                 reg600,
                 reg597,
                 forvar595,
                 reg593,
                 forvar591,
                 reg590,
                 reg588,
                 reg587,
                 forvar584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 reg578,
                 forvar577,
                 forvar576,
                 reg574,
                 reg570,
                 reg568,
                 reg567,
                 forvar565,
                 reg563,
                 reg560,
                 reg559,
                 forvar557,
                 reg556,
                 forvar555,
                 forvar554,
                 reg553,
                 reg550,
                 forvar548,
                 forvar547,
                 reg545,
                 reg544,
                 forvar541,
                 reg540,
                 reg538,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg521,
                 forvar502,
                 reg527,
                 reg526,
                 reg524,
                 reg523,
                 forvar521,
                 reg518,
                 reg517,
                 reg513,
                 reg509,
                 reg508,
                 reg507,
                 reg505,
                 reg504,
                 reg502,
                 reg501,
                 reg499,
                 reg496,
                 forvar487,
                 reg494,
                 reg492,
                 reg491,
                 reg488,
                 reg487,
                 reg483,
                 reg481,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 forvar474,
                 forvar473,
                 reg472,
                 reg471,
                 reg470,
                 reg468,
                 reg465,
                 reg464,
                 reg462,
                 reg461,
                 reg459,
                 reg453,
                 forvar451,
                 reg449,
                 reg448,
                 reg446,
                 reg445,
                 forvar444,
                 reg441,
                 reg440,
                 forvar437,
                 reg436,
                 reg435,
                 reg432,
                 (1'h0)};
  assign wire431 = $unsigned(wire430);
  always
    @(posedge clk) begin
      reg432 = ((8'ha6) ?
          wire427[(1'h1):(1'h1)] : (^~((&wire428[(3'h4):(1'h0)]) ?
              $unsigned(wire427) : (~wire429))));
    end
  always
    @(posedge clk) begin
      if (((wire425 == {$signed((~^wire431)),
          ($signed(wire426) <<< (wire429 ? wire426 : (8'hbe))),
          ($signed(wire426) & (wire425 ?
              wire427 : wire428))}) - ($signed(wire430) ?
          ({$unsigned((7'h46)),
              (wire427 & (8'ha2)),
              {wire430}} << wire425[(1'h0):(1'h0)]) : $signed($unsigned({wire428,
              wire429})))))
        begin
          reg433 <= wire427;
          if ((&reg433))
            begin
              reg434 <= ($unsigned((^~wire430[(2'h2):(1'h0)])) ?
                  $unsigned(wire428) : wire429[(3'h5):(3'h4)]);
            end
          else
            begin
              reg435 = (7'h4d);
              reg436 = wire427[(2'h3):(2'h2)];
              reg437 <= (~reg435[(5'h19):(4'he)]);
              reg438 <= wire430[(5'h12):(4'hc)];
              reg439 <= (~wire431);
            end
        end
      else
        begin
          reg435 = reg435;
          reg436 = (~&$signed($signed((|(^~(8'hab))))));
          for (forvar437 = (1'h0); (forvar437 < (3'h6)); forvar437 = (forvar437 + (1'h1)))
            begin
              reg438 <= (((((7'h40) << wire425[(1'h1):(1'h0)]) ?
                          ((~&(7'h45)) ?
                              $unsigned(forvar437) : reg434) : (((8'hbb) ?
                              wire426 : (8'ha5)) <<< $signed(reg438))) ?
                      {$unsigned((wire428 ? reg437 : reg437)),
                          ({reg438} != $unsigned(forvar437))} : forvar437) ?
                  reg438[(1'h0):(1'h0)] : wire431[(2'h2):(1'h1)]);
              reg439 <= reg438;
              reg440 = ((~^wire428) != (~|{{(wire426 ? wire426 : reg436)}}));
              reg441 = $unsigned(forvar437[(3'h4):(2'h3)]);
              reg442 <= ({$unsigned($unsigned((!reg436))),
                  {reg438[(2'h2):(1'h0)],
                      reg434[(5'h14):(5'h11)]}} != {$unsigned(reg439),
                  ($unsigned(wire425) ^~ ((wire431 * (8'hb6)) ?
                      $signed(reg441) : {reg433, reg438, (7'h47)}))});
            end
          reg443 <= $unsigned(($unsigned((reg442 - (reg442 ~^ wire431))) ?
              (($signed(wire428) ? (reg438 ? reg433 : wire429) : reg435) ?
                  {wire425,
                      wire430[(5'h14):(4'he)]} : {reg437[(3'h5):(2'h2)]}) : reg434));
          for (forvar444 = (1'h0); (forvar444 < (1'h1)); forvar444 = (forvar444 + (1'h1)))
            begin
              reg445 = (&reg437[(3'h6):(3'h5)]);
              reg446 = (wire427 >> (reg437[(1'h1):(1'h1)] >> (~|wire430)));
              reg447 <= reg435;
              reg448 = $signed(reg433);
              reg449 = $signed(((|$signed(reg438)) ?
                  {{reg437, forvar437, $unsigned(forvar437)},
                      reg434} : (7'h58)));
              reg450 <= wire431[(5'h18):(3'h4)];
            end
          for (forvar451 = (1'h0); (forvar451 < (3'h6)); forvar451 = (forvar451 + (1'h1)))
            begin
              reg452 <= $unsigned((^{$unsigned(reg449), $signed((~|reg450))}));
              reg453 = ($signed(((^~wire429) ? (7'h47) : (~|(|(7'h4a))))) ?
                  {(&(-reg439))} : {$unsigned($signed($unsigned(reg452)))});
              reg454 <= (($unsigned((^$signed(reg447))) ?
                  $signed(wire426[(5'h10):(2'h3)]) : ((reg443[(4'hd):(4'h8)] ?
                      reg435 : ((8'hbf) ?
                          wire431 : reg434)) || reg449[(3'h7):(3'h7)])) * $signed(reg438[(3'h4):(3'h4)]));
              reg455 <= reg448[(3'h7):(1'h0)];
              reg456 <= (!$signed(reg452[(3'h7):(2'h3)]));
              reg457 <= {(~&{{$unsigned((7'h4d)), reg436, ((7'h48) ^~ reg446)},
                      {(reg448 ? reg454 : reg446), {forvar437}, (+wire429)}}),
                  {reg446,
                      {({reg442} ?
                              $unsigned(reg455) : (reg454 ? reg456 : reg456)),
                          $unsigned($signed(reg445)),
                          $signed((|wire425))},
                      $unsigned((|(reg441 ? wire430 : wire429)))},
                  {(reg447 ?
                          {(forvar437 ? (7'h4b) : forvar451),
                              reg447[(2'h3):(1'h0)]} : reg449[(3'h4):(1'h0)]),
                      $unsigned($signed({reg442, reg452, wire425}))}};
            end
          reg458 <= $signed($unsigned($unsigned(wire425[(1'h1):(1'h1)])));
        end
    end
  always
    @(posedge clk) begin
      reg459 = {($unsigned($signed((8'haa))) ~^ wire426[(4'he):(4'ha)]),
          wire425[(1'h1):(1'h0)],
          ($signed($unsigned($unsigned((8'ha6)))) >>> {$unsigned($signed(wire431)),
              (^~(wire427 ~^ wire425))})};
      reg460 <= reg458;
      if ($signed(wire429))
        begin
          reg461 = (reg459[(4'h9):(3'h6)] ?
              $unsigned(($unsigned((|wire426)) ?
                  (~&$signed(reg452)) : ((~|wire430) ^~ $signed(wire430)))) : reg454[(2'h3):(2'h2)]);
          reg462 = (+(8'hbf));
          reg463 <= $signed($unsigned((~|(reg454[(4'h8):(4'h8)] ?
              (reg438 ? (8'ha4) : reg439) : reg455[(3'h6):(2'h2)]))));
          reg464 = ($unsigned($signed($signed($signed(reg452)))) ?
              reg439[(2'h3):(1'h1)] : ($unsigned($unsigned({reg443})) < (~($signed(reg462) ?
                  (wire428 == (8'hbf)) : reg438[(1'h0):(1'h0)]))));
          reg465 = $signed($signed((reg452 ~^ reg461[(5'h15):(3'h5)])));
          reg466 <= ($signed((wire427[(1'h0):(1'h0)] ?
                  ($signed(reg450) ^~ $signed(reg452)) : $signed((wire428 ?
                      reg457 : (8'haa))))) ?
              reg450[(3'h4):(1'h0)] : ((reg463 ?
                  reg452 : reg437[(3'h6):(3'h4)]) && ($signed($signed(wire426)) ?
                  (+((8'ha6) ? reg465 : reg463)) : wire427[(1'h0):(1'h0)])));
          reg467 <= wire426[(1'h0):(1'h0)];
        end
      else
        begin
          if ($signed(reg460))
            begin
              reg461 = reg462;
              reg462 = $unsigned(({(reg467 & {(7'h57),
                      reg458,
                      reg433})} < {(reg437 ? reg455 : $unsigned((8'ha1))),
                  wire427,
                  ({(7'h41), (7'h52)} ?
                      $signed(reg433) : (reg454 >= reg439))}));
              reg464 = wire428;
              reg465 = (!((&(reg465[(3'h6):(1'h1)] << (8'hbb))) ?
                  (($signed(wire431) ? {reg458} : (reg434 ? reg460 : reg463)) ?
                      reg437[(3'h6):(3'h5)] : reg462[(5'h15):(3'h5)]) : $unsigned(wire427[(1'h0):(1'h0)])));
              reg468 = {reg455};
            end
          else
            begin
              reg463 <= (^reg438);
              reg464 = reg450[(3'h7):(3'h4)];
              reg466 <= (wire426[(1'h1):(1'h0)] ?
                  (~$unsigned((~(~|reg464)))) : {(((wire425 ?
                                  (8'ha4) : reg434) ?
                              (reg454 ? wire429 : reg455) : $unsigned(reg434)) ?
                          {reg439[(4'hf):(3'h5)]} : (~^$signed(reg466)))});
            end
        end
      reg469 <= (-(wire427 ?
          (reg456 ?
              $unsigned({reg439,
                  wire426}) : reg437[(3'h6):(1'h1)]) : reg455[(4'hb):(3'h7)]));
      reg470 = (~|((~^reg437[(3'h4):(3'h4)]) ?
          reg438[(2'h3):(2'h2)] : $signed($unsigned($signed((8'haf))))));
      reg471 = $unsigned(reg468);
      reg472 = $unsigned(reg467);
    end
  always
    @(posedge clk) begin
      for (forvar473 = (1'h0); (forvar473 < (1'h0)); forvar473 = (forvar473 + (1'h1)))
        begin
          for (forvar474 = (1'h0); (forvar474 < (3'h6)); forvar474 = (forvar474 + (1'h1)))
            begin
              reg475 = ($signed((+($unsigned(wire428) ?
                  ((7'h4c) >> (8'hbb)) : {forvar474,
                      wire429}))) <<< reg454[(2'h3):(2'h3)]);
              reg476 = $signed($unsigned($unsigned(($unsigned(wire427) ?
                  (forvar473 <<< reg457) : (reg475 ? wire428 : reg434)))));
              reg477 = $signed({reg439});
            end
          if (reg457)
            begin
              reg478 = (-($unsigned((^(wire431 > (8'ha7)))) & (($unsigned((7'h53)) ?
                      $signed(reg434) : (wire431 - reg467)) ?
                  (|$unsigned(reg469)) : (&(reg452 ? wire426 : reg456)))));
              reg479 = $signed((~&reg457));
              reg480 = wire431[(4'hf):(2'h2)];
              reg481 = $signed($signed($unsigned((!$unsigned(reg457)))));
            end
          else
            begin
              reg478 = (~&reg455[(1'h1):(1'h0)]);
              reg482 <= reg476[(3'h7):(3'h6)];
              reg483 = reg463;
              reg484 <= reg437;
              reg485 <= $signed(reg454);
            end
          reg486 <= {$unsigned($signed((!$unsigned(reg478))))};
        end
      if ($signed(forvar473[(2'h2):(1'h1)]))
        begin
          reg487 = reg456[(3'h6):(2'h3)];
          if ((7'h52))
            begin
              reg488 = ($signed(wire427) + reg450[(3'h7):(1'h1)]);
              reg489 <= ({$unsigned($signed((~|reg442))),
                      ($signed($signed(reg483)) & (~|reg480[(1'h1):(1'h0)])),
                      wire431} ?
                  (reg438[(2'h2):(1'h1)] ?
                      wire425 : ($signed(reg481) | ($signed((7'h52)) ?
                          (reg478 << reg466) : (~reg488)))) : $signed((reg437 || reg467)));
              reg490 <= reg460;
              reg491 = $unsigned((^($unsigned((^reg476)) >= reg460)));
              reg492 = reg486;
            end
          else
            begin
              reg488 = $unsigned({{forvar473[(1'h0):(1'h0)]}});
              reg491 = wire431;
              reg493 <= (-wire430);
              reg494 = $unsigned($signed(reg433));
              reg495 <= reg482[(3'h4):(2'h2)];
            end
        end
      else
        begin
          for (forvar487 = (1'h0); (forvar487 < (3'h6)); forvar487 = (forvar487 + (1'h1)))
            begin
              reg488 = reg460[(4'he):(4'he)];
              reg491 = (-(+wire425[(2'h2):(2'h2)]));
              reg493 <= (~reg482[(3'h6):(2'h3)]);
              reg494 = ((7'h53) < forvar487);
              reg496 = (+reg492[(3'h5):(1'h1)]);
              reg497 <= $unsigned((+reg463));
            end
          if ($unsigned((^(reg480[(5'h12):(4'ha)] ?
              reg457[(2'h3):(1'h1)] : $signed($signed(reg482))))))
            begin
              reg498 <= (^~reg495);
              reg499 = ((forvar487 ?
                      $signed({(reg483 ?
                              forvar474 : reg442)}) : $unsigned(reg447)) ?
                  forvar487[(5'h14):(2'h2)] : reg447);
              reg500 <= reg495[(4'h8):(3'h5)];
            end
          else
            begin
              reg499 = (forvar473[(2'h2):(1'h1)] ?
                  reg438[(3'h4):(1'h0)] : $signed({$signed($signed((7'h56))),
                      (wire431[(5'h14):(4'h9)] ?
                          $unsigned(reg476) : $unsigned(reg457))}));
              reg501 = reg457;
            end
        end
      if (($unsigned(reg442[(3'h7):(3'h5)]) ? reg454[(3'h7):(3'h7)] : reg476))
        begin
          if ((&reg483[(5'h1a):(5'h13)]))
            begin
              reg502 = $signed($signed((^(~&reg452))));
              reg503 <= reg442;
              reg504 = $unsigned(reg475[(4'h8):(3'h5)]);
              reg505 = ((|reg501[(5'h11):(4'he)]) >> (+$signed(reg500)));
            end
          else
            begin
              reg502 = ((reg479[(1'h1):(1'h0)] ?
                  reg475 : $signed((^~reg490[(1'h0):(1'h0)]))) * reg490[(2'h3):(2'h3)]);
            end
          reg506 <= (~(~|{$unsigned($unsigned(reg478)),
              reg447,
              reg494[(1'h1):(1'h1)]}));
          if (((|($signed((reg479 || reg475)) || (~|reg494[(4'he):(4'hd)]))) ?
              $unsigned((~^($unsigned(wire431) * (+reg482)))) : {wire428,
                  (&$unsigned((8'ha2)))}))
            begin
              reg507 = $unsigned(reg497[(1'h1):(1'h1)]);
              reg508 = reg454[(1'h1):(1'h1)];
              reg509 = reg486;
              reg510 <= ((reg492[(1'h1):(1'h1)] < (|($unsigned((7'h45)) << (reg490 ?
                  reg456 : wire426)))) + {(($signed(reg488) ?
                          (~reg478) : $unsigned(reg455)) ?
                      $signed(reg484[(4'hb):(4'ha)]) : (reg489[(5'h12):(3'h4)] || reg509[(2'h2):(1'h0)])),
                  (7'h58)});
              reg511 <= $signed((~&reg455[(4'he):(4'h9)]));
              reg512 <= (-wire431);
            end
          else
            begin
              reg507 = reg447;
              reg510 <= reg491[(1'h1):(1'h0)];
              reg511 <= reg499[(3'h7):(1'h1)];
              reg513 = $unsigned(reg511[(1'h0):(1'h0)]);
              reg514 <= reg447;
              reg515 <= {$signed((8'haa)),
                  (~|$unsigned(reg506)),
                  ((((wire430 == reg497) ?
                      {(8'ha2),
                          reg507} : (reg442 << (7'h54))) && {(reg454 | (7'h48)),
                      $unsigned(reg458)}) >>> (~^$signed((reg442 >= reg497))))};
            end
          if (reg495)
            begin
              reg516 <= {(+reg482),
                  ((~^$signed(reg514[(1'h0):(1'h0)])) ?
                      ((reg499 ? $signed(reg463) : reg513[(4'h9):(2'h3)]) ?
                          (^reg479[(3'h5):(2'h3)]) : reg455[(4'ha):(4'ha)]) : reg490),
                  {(reg447[(3'h4):(2'h2)] == ((~&reg499) ? reg503 : reg486)),
                      reg481[(2'h3):(1'h0)]}};
              reg517 = ($unsigned((~&$unsigned(reg496))) ?
                  $signed(((7'h45) ?
                      (~(reg484 ?
                          reg483 : reg454)) : (~^reg439[(2'h2):(1'h0)]))) : $signed($unsigned(reg505[(1'h1):(1'h1)])));
              reg518 = reg483[(2'h3):(1'h0)];
              reg519 <= (reg433[(4'hf):(3'h7)] ^ $signed((reg493 ?
                  reg508 : reg442)));
            end
          else
            begin
              reg516 <= ((^reg517[(2'h2):(2'h2)]) && (^~reg494[(3'h7):(1'h0)]));
              reg519 <= reg495;
              reg520 <= (+($signed((-$signed(reg487))) ^~ (reg498 ~^ $signed(reg496[(1'h0):(1'h0)]))));
            end
          for (forvar521 = (1'h0); (forvar521 < (1'h0)); forvar521 = (forvar521 + (1'h1)))
            begin
              reg522 <= (|((~|((~|forvar521) ?
                      $signed(reg487) : $unsigned(reg501))) ?
                  $unsigned(reg486) : reg495[(4'hc):(4'hc)]));
            end
          if (reg508)
            begin
              reg523 = reg475[(2'h2):(1'h1)];
              reg524 = reg501[(4'h9):(2'h2)];
              reg525 <= reg496[(3'h4):(2'h2)];
              reg526 = $signed((+(~^(reg502 ~^ (^~reg519)))));
              reg527 = (^~reg511);
            end
          else
            begin
              reg523 = $unsigned((reg452[(3'h6):(3'h6)] & {(wire425 ?
                      {reg495, reg438, wire430} : wire430),
                  reg485[(3'h6):(3'h6)]}));
              reg524 = $unsigned(reg518);
              reg526 = {reg487,
                  (|{{$unsigned(reg522), (8'hab)},
                      (reg478[(2'h3):(1'h0)] >= (8'hb3)),
                      $signed($signed(reg491))}),
                  reg497};
              reg527 = $signed((^(($unsigned((8'hbf)) ?
                  reg438 : reg507) > ($unsigned(reg514) ?
                  reg508 : reg466[(4'ha):(4'h9)]))));
              reg528 <= (+reg509[(4'h9):(4'h8)]);
              reg529 <= (reg476 ^~ reg503);
              reg530 <= (((reg454 ?
                          $signed(reg520[(1'h1):(1'h0)]) : $unsigned((~&reg520))) ?
                      $signed((~^reg458[(3'h5):(3'h4)])) : ((+(reg509 ?
                          reg527 : reg503)) & (8'ha6))) ?
                  (8'ha6) : (|$signed(reg500)));
            end
        end
      else
        begin
          for (forvar502 = (1'h0); (forvar502 < (2'h2)); forvar502 = (forvar502 + (1'h1)))
            begin
              reg503 <= (reg442[(3'h7):(1'h1)] ?
                  {$signed($unsigned(reg515)), reg484[(1'h0):(1'h0)]} : reg501);
              reg504 = $unsigned(wire425);
              reg506 <= $unsigned({(-$signed((^reg476)))});
              reg510 <= $signed(reg456);
              reg511 <= $signed(($signed((reg443 ?
                      $signed((8'ha4)) : (+reg515))) ?
                  reg490 : $signed({{reg457, wire425, reg480},
                      (reg475 ? (8'hb6) : reg515),
                      reg460[(5'h10):(4'hb)]})));
            end
          if (reg492)
            begin
              reg512 <= $signed({((forvar487[(3'h7):(3'h5)] ?
                          {reg509} : reg520) ?
                      {$signed((7'h51)),
                          (^~forvar521),
                          reg525[(3'h5):(1'h1)]} : reg512)});
              reg514 <= $signed($signed($signed((reg511[(2'h2):(1'h1)] ?
                  $signed(reg515) : (~^reg488)))));
              reg517 = {(($signed(reg519[(4'h9):(2'h3)]) ?
                      (forvar487[(5'h1c):(5'h1b)] >>> reg501) : (8'hbd)) + $signed($signed($unsigned(reg460)))),
                  $signed(reg523[(1'h1):(1'h0)])};
              reg519 <= ((reg476[(3'h5):(2'h2)] ?
                      reg466[(2'h3):(2'h3)] : {wire430}) ?
                  (($signed(reg502[(5'h16):(3'h7)]) ?
                      reg457 : (reg514[(1'h0):(1'h0)] ?
                          (~^reg467) : (reg452 << reg514))) >> (~^forvar521)) : reg497);
              reg520 <= $unsigned(reg517[(4'hc):(3'h7)]);
              reg521 = ((($signed($signed(forvar473)) * reg438) ?
                      ({$signed(reg494), $unsigned(wire425)} ?
                          reg483 : ($signed(reg493) ?
                              (reg483 <<< (7'h53)) : $unsigned(reg458))) : $signed($signed((~^reg506)))) ?
                  (~(!$unsigned((reg489 | reg457)))) : (reg460 >> {reg499[(5'h10):(2'h2)],
                      $unsigned(reg509[(1'h0):(1'h0)]),
                      ((reg477 ? (8'hac) : reg443) ? (~&reg499) : wire428)}));
              reg523 = (&(reg511 ?
                  $signed(((reg456 * wire431) * (reg528 ?
                      reg511 : reg463))) : $unsigned({(~^(8'hb0)),
                      {reg439, wire426, reg530}})));
            end
          else
            begin
              reg513 = reg515;
              reg517 = reg495[(4'ha):(2'h3)];
              reg519 <= (|((~&(reg527[(4'ha):(2'h3)] < (reg520 * wire429))) + (reg469[(4'h8):(3'h5)] | $signed((reg530 > reg518)))));
              reg520 <= (8'hb3);
              reg521 = ({({reg450[(3'h7):(1'h0)]} ?
                      ($signed((7'h51)) && $signed(reg483)) : (7'h42))} + {{(~|$unsigned((7'h50))),
                      $signed((reg450 ? reg484 : reg442)),
                      (~&reg493)},
                  reg485[(4'h9):(4'h8)],
                  (~^(((8'hb5) ? reg516 : wire428) ?
                      reg460 : $unsigned(reg469)))});
            end
          if ($signed(((^{$unsigned(reg496), (8'hb2)}) * {$signed((-reg512)),
              $signed((reg516 ? reg457 : reg499)),
              {$unsigned(reg479), $unsigned(wire428), (&wire431)}})))
            begin
              reg524 = $unsigned((~&(($signed(wire429) ?
                  reg526[(2'h3):(2'h3)] : reg502[(5'h13):(4'hf)]) > (wire427[(2'h2):(1'h1)] ?
                  (forvar521 || (7'h4d)) : (reg450 ? reg484 : forvar474)))));
              reg526 = reg439;
              reg528 <= (~&reg495);
            end
          else
            begin
              reg525 <= reg438[(1'h0):(1'h0)];
              reg526 = (~(~&$signed(forvar473[(1'h1):(1'h1)])));
              reg528 <= reg519;
              reg529 <= ({reg434} ?
                  {reg486,
                      {{(~reg434), ((8'hb7) ? reg496 : reg486)},
                          (&reg488),
                          $unsigned((wire427 <<< forvar521))},
                      reg498} : (~&(reg515[(3'h5):(2'h2)] >>> reg466)));
              reg530 <= ({reg438[(2'h3):(1'h1)],
                  $signed(reg443),
                  forvar502[(4'ha):(3'h5)]} - $signed($unsigned({reg478[(5'h18):(5'h13)]})));
              reg531 = ((reg524[(5'h18):(3'h7)] - reg503[(1'h0):(1'h0)]) ?
                  $unsigned(reg518[(3'h5):(1'h1)]) : ($signed(reg490[(2'h2):(1'h0)]) >> reg505[(4'h9):(4'h9)]));
            end
          if ((~&$unsigned((reg483[(5'h18):(5'h14)] <= (~^(reg487 >= wire431))))))
            begin
              reg532 = reg488;
              reg533 = {(reg516 != reg513[(2'h2):(1'h1)]),
                  reg492[(4'hc):(3'h6)]};
              reg534 = (&$signed($unsigned($unsigned((reg478 << reg529)))));
              reg535 = (7'h40);
              reg536 = reg525[(4'ha):(3'h6)];
              reg537 <= ((-reg485) ^~ (reg491 < reg439));
              reg538 = (8'hb6);
            end
          else
            begin
              reg532 = $unsigned(reg527[(5'h1e):(4'hb)]);
              reg537 <= $signed((|$unsigned($signed((reg488 != (8'hbb))))));
              reg538 = $unsigned(($signed(reg488) & reg447));
              reg539 <= $signed(reg523[(5'h12):(4'h8)]);
              reg540 = reg531[(3'h5):(2'h2)];
            end
          for (forvar541 = (1'h0); (forvar541 < (2'h3)); forvar541 = (forvar541 + (1'h1)))
            begin
              reg542 <= (~^{$signed((^~(8'hab))),
                  (+$unsigned(((7'h51) == reg501)))});
              reg543 <= (reg499 ?
                  ({((&forvar487) > (reg447 ? forvar473 : reg529))} ?
                      reg433 : ($signed((reg515 ^ reg532)) ?
                          {reg500, reg521} : (^$unsigned(reg434)))) : reg519);
              reg544 = forvar502[(2'h3):(1'h1)];
              reg545 = ($signed(reg443[(5'h1a):(5'h14)]) ?
                  (($unsigned((reg486 ?
                      wire429 : reg499)) >>> $unsigned($signed(reg525))) * reg502[(4'hc):(4'hb)]) : $unsigned($signed($signed((reg543 ?
                      reg501 : reg522)))));
              reg546 <= reg495[(3'h7):(3'h5)];
            end
        end
      for (forvar547 = (1'h0); (forvar547 < (1'h1)); forvar547 = (forvar547 + (1'h1)))
        begin
          for (forvar548 = (1'h0); (forvar548 < (3'h4)); forvar548 = (forvar548 + (1'h1)))
            begin
              reg549 <= (^~reg493[(4'hf):(3'h7)]);
              reg550 = (8'ha6);
              reg551 <= $signed({(^($unsigned((7'h4a)) ^~ (reg434 == reg536))),
                  reg469});
              reg552 <= $unsigned({reg489});
              reg553 = reg511[(2'h2):(1'h1)];
            end
        end
      for (forvar554 = (1'h0); (forvar554 < (1'h1)); forvar554 = (forvar554 + (1'h1)))
        begin
          for (forvar555 = (1'h0); (forvar555 < (3'h4)); forvar555 = (forvar555 + (1'h1)))
            begin
              reg556 = (reg502 ?
                  $unsigned(($unsigned($signed(reg535)) <<< (reg528 ~^ (reg501 >>> reg504)))) : (^~reg484));
            end
          for (forvar557 = (1'h0); (forvar557 < (3'h5)); forvar557 = (forvar557 + (1'h1)))
            begin
              reg558 <= reg532;
              reg559 = reg482[(1'h1):(1'h1)];
              reg560 = $signed((({{(8'hbf),
                      reg506}} + $unsigned({reg509})) ^ (((reg543 >>> reg545) == reg552[(3'h6):(1'h0)]) != ($signed(reg510) && reg553))));
              reg561 <= $signed($signed((8'haf)));
              reg562 <= $unsigned($signed(($signed(reg514) ?
                  $unsigned(((8'ha6) <<< (7'h4e))) : $signed((reg556 ~^ reg447)))));
            end
          reg563 = reg452[(3'h4):(2'h2)];
        end
    end
  assign wire564 = reg549;
  always
    @(posedge clk) begin
      for (forvar565 = (1'h0); (forvar565 < (1'h1)); forvar565 = (forvar565 + (1'h1)))
        begin
          if (((reg525[(2'h3):(1'h0)] ?
                  ($signed({wire430}) ?
                      $signed({reg512,
                          reg561}) : reg443[(4'h8):(3'h5)]) : wire425[(2'h2):(1'h1)]) ?
              $unsigned($signed(((reg514 && reg500) | $signed(reg515)))) : ((forvar565[(2'h2):(1'h0)] ?
                      (reg458 && (reg539 || reg452)) : ($unsigned(reg438) ?
                          $unsigned(reg562) : $signed((8'ha6)))) ?
                  $unsigned((wire427 ?
                      $signed((8'haf)) : reg484[(1'h0):(1'h0)])) : reg434[(4'h8):(2'h3)])))
            begin
              reg566 <= reg437[(2'h2):(1'h0)];
              reg567 = (!(&(^$signed(reg537[(5'h16):(3'h6)]))));
              reg568 = (!{(~^reg457),
                  ($unsigned($signed((8'hb7))) ?
                      (^~(reg447 >>> reg510)) : (~^(reg452 ?
                          reg438 : reg561)))});
              reg569 <= reg529;
              reg570 = $signed(($signed(($unsigned((7'h57)) ?
                      (-reg500) : (^~reg516))) ?
                  (reg437[(1'h1):(1'h0)] ?
                      $signed($unsigned(reg455)) : ((&reg525) ?
                          (forvar565 && reg469) : reg452)) : ((!reg493) ?
                      $signed((^reg569)) : (|(-reg516)))));
            end
          else
            begin
              reg567 = ({$unsigned($unsigned(reg542[(1'h0):(1'h0)]))} > {(~|wire425[(1'h1):(1'h1)]),
                  (7'h4a),
                  reg546});
              reg568 = reg497;
              reg569 <= $unsigned(reg519[(5'h14):(3'h5)]);
              reg571 <= $unsigned(wire425[(1'h1):(1'h0)]);
              reg572 <= (~&forvar565);
            end
          reg573 <= $signed($signed(reg469[(5'h13):(1'h0)]));
          reg574 = ((($unsigned((reg495 || wire427)) ?
                      (8'ha3) : (reg512 || (!reg443))) ?
                  $unsigned((~^$unsigned(reg458))) : reg512) ?
              $signed({reg463[(5'h13):(4'ha)]}) : reg571);
          reg575 <= $unsigned(($signed($unsigned(reg542[(1'h1):(1'h0)])) ?
              reg442[(3'h7):(2'h3)] : (wire564 == ($unsigned(reg549) <= $signed((7'h43))))));
        end
      for (forvar576 = (1'h0); (forvar576 < (3'h6)); forvar576 = (forvar576 + (1'h1)))
        begin
          for (forvar577 = (1'h0); (forvar577 < (1'h0)); forvar577 = (forvar577 + (1'h1)))
            begin
              reg578 = (reg512 ? $signed(wire564[(1'h1):(1'h1)]) : reg493);
              reg579 <= ($signed($signed(((8'hb6) ^ (wire429 && (8'hbd))))) & (&$signed((reg561[(3'h7):(3'h5)] || wire426[(5'h13):(3'h7)]))));
              reg580 = reg516[(3'h5):(1'h1)];
              reg581 = ((~^{{(8'hb6)}}) ? (|(~&(~reg458))) : (&reg579));
              reg582 = ($signed({{{wire425, reg574}},
                      $unsigned((7'h40)),
                      {(wire428 + reg497)}}) ?
                  (^~(reg458 + $unsigned($signed(reg466)))) : reg514);
              reg583 = $signed($unsigned(reg456));
            end
          for (forvar584 = (1'h0); (forvar584 < (2'h3)); forvar584 = (forvar584 + (1'h1)))
            begin
              reg585 <= reg571;
            end
          if (((($signed(reg529) ?
                  (~reg568) : $unsigned((reg438 ? wire431 : reg434))) ?
              ((~|(reg525 ?
                  (7'h40) : reg443)) >= $signed((|reg485))) : {reg514[(2'h2):(1'h0)],
                  ((reg460 & reg539) ? wire425 : forvar584[(4'h8):(1'h0)]),
                  (~^(reg447 ? reg519 : reg522))}) != reg570[(1'h1):(1'h1)]))
            begin
              reg586 <= reg510[(4'hf):(2'h3)];
              reg587 = $signed(((|wire431) * ($signed((forvar565 ?
                      reg529 : reg447)) ?
                  reg510 : $signed((~^reg515)))));
              reg588 = reg572;
              reg589 <= $unsigned((reg497[(3'h4):(1'h1)] ?
                  reg574 : $signed($unsigned((reg467 | reg578)))));
              reg590 = (reg514[(2'h3):(1'h0)] > wire430[(4'hd):(4'hd)]);
            end
          else
            begin
              reg587 = ($signed((!$signed((|reg552)))) != ($unsigned(reg539) ?
                  $signed(((reg562 ?
                      reg519 : reg519) * (^~reg575))) : reg566[(4'hc):(3'h7)]));
              reg588 = $signed((~^$unsigned((|reg572))));
            end
          for (forvar591 = (1'h0); (forvar591 < (3'h6)); forvar591 = (forvar591 + (1'h1)))
            begin
              reg592 <= reg586;
              reg593 = $unsigned((|reg485[(1'h0):(1'h0)]));
            end
        end
    end
  assign wire594 = ($signed(($unsigned((reg460 != (7'h56))) == $signed(reg546[(3'h4):(2'h2)]))) ?
                       (~^$unsigned((~|((7'h58) - (8'hbe))))) : $signed((&((~^reg498) <= reg551[(5'h10):(2'h2)]))));
  always
    @(posedge clk) begin
      for (forvar595 = (1'h0); (forvar595 < (3'h4)); forvar595 = (forvar595 + (1'h1)))
        begin
          if ($signed(wire426[(5'h18):(3'h6)]))
            begin
              reg596 <= reg520[(2'h3):(1'h0)];
              reg597 = ((reg433 ?
                  wire429[(3'h5):(2'h2)] : (^(-$unsigned(reg511)))) ~^ ((7'h53) & (^~$unsigned(wire564[(1'h0):(1'h0)]))));
              reg598 <= $signed(reg493[(5'h15):(5'h15)]);
              reg599 <= $signed({$unsigned(reg572[(4'he):(4'h9)]),
                  reg443,
                  reg519[(4'h8):(4'h8)]});
            end
          else
            begin
              reg596 <= reg452[(3'h5):(3'h4)];
              reg598 <= (~^{$unsigned((~reg485[(2'h3):(2'h3)])),
                  (((8'hb8) ?
                      $signed(reg439) : reg458[(2'h2):(1'h0)]) <<< (reg437 | (reg466 << wire594)))});
            end
          reg600 = wire564;
          for (forvar601 = (1'h0); (forvar601 < (3'h4)); forvar601 = (forvar601 + (1'h1)))
            begin
              reg602 = (8'ha8);
              reg603 <= (($signed((7'h46)) ?
                  reg486[(1'h0):(1'h0)] : (~^reg485[(4'h8):(3'h5)])) != (~|($signed(((8'ha8) ?
                      reg439 : reg572)) ?
                  reg520[(1'h0):(1'h0)] : $signed($unsigned(reg515)))));
              reg604 <= {$unsigned({($signed(reg572) ?
                          $signed(reg543) : (~|reg525))}),
                  $signed(reg458[(1'h0):(1'h0)])};
            end
          if ({$signed(wire430),
              $unsigned(({(reg528 ? reg603 : reg561), reg433} ?
                  ($signed(reg530) ?
                      (reg571 ?
                          reg525 : reg558) : $unsigned(reg437)) : ((wire429 ?
                      reg519 : reg442) << $unsigned((8'ha3))))),
              reg520[(2'h3):(1'h1)]})
            begin
              reg605 <= ($unsigned(reg586[(5'h17):(4'he)]) == (&(~&$signed((8'ha4)))));
              reg606 <= (~|{(!((reg467 <= reg519) ? (~(7'h55)) : (8'hb0))),
                  reg510[(1'h1):(1'h0)]});
              reg607 <= ($unsigned((~|((reg603 ~^ reg549) ?
                      (wire426 && reg586) : reg443))) ?
                  (reg450 << wire564) : (reg599[(4'h8):(3'h6)] <= (~&($unsigned(reg522) ?
                      (7'h56) : reg463[(4'ha):(4'h8)]))));
              reg608 = ((^reg549[(4'ha):(1'h1)]) ^ {reg539,
                  $signed(reg450),
                  $unsigned(reg457[(1'h1):(1'h1)])});
              reg609 = (!(7'h43));
            end
          else
            begin
              reg608 = (reg566 >>> {$unsigned($unsigned((8'hbc))),
                  (^reg506[(1'h0):(1'h0)]),
                  reg485});
              reg609 = (reg608 ?
                  (($signed($unsigned(reg466)) << (8'ha6)) ^ ((~|reg579[(3'h6):(3'h4)]) ?
                      reg510 : reg561)) : (&(reg455 ~^ $signed(reg571))));
              reg610 = (~^$signed(((~&reg596[(4'he):(3'h4)]) ?
                  (~&(&reg514)) : ((~&reg561) & (&reg543)))));
              reg611 <= (reg552[(3'h5):(1'h0)] >= reg573[(4'h9):(3'h6)]);
              reg612 = reg467;
            end
          reg613 <= (-$unsigned(($signed($signed(reg515)) & {wire430,
              (reg600 + reg510)})));
          if (reg539[(4'h9):(3'h6)])
            begin
              reg614 = $signed(($unsigned($unsigned((reg606 + reg589))) <<< ($unsigned(reg597[(3'h5):(2'h3)]) ?
                  $signed($unsigned(reg539)) : $signed((|reg589)))));
            end
          else
            begin
              reg615 <= $signed(reg575[(2'h3):(2'h2)]);
              reg616 <= (&wire564[(4'h9):(3'h4)]);
              reg617 = reg433[(4'ha):(1'h0)];
              reg618 = reg615[(3'h4):(3'h4)];
            end
        end
      for (forvar619 = (1'h0); (forvar619 < (2'h3)); forvar619 = (forvar619 + (1'h1)))
        begin
          reg620 <= ((~^($signed((reg455 >> (8'haf))) ? reg466 : (^~(8'ha3)))) ?
              reg537[(4'hb):(1'h0)] : ((((~&reg602) << (7'h58)) || ((reg562 ?
                      reg439 : reg529) >>> reg542)) ?
                  wire431 : ((~&reg598[(3'h6):(3'h6)]) ?
                      ((reg566 && reg592) - (^reg614)) : {(wire429 <<< reg585),
                          (reg609 >= reg500),
                          {(8'ha3), reg608}})));
          for (forvar621 = (1'h0); (forvar621 < (2'h2)); forvar621 = (forvar621 + (1'h1)))
            begin
              reg622 = reg455[(4'ha):(2'h2)];
              reg623 = (($unsigned($signed($signed(reg516))) || (+reg439)) ?
                  reg613[(4'h9):(3'h4)] : ($unsigned($signed(reg618)) ?
                      reg546[(1'h1):(1'h0)] : $signed(reg454[(3'h7):(3'h7)])));
              reg624 = reg623;
              reg625 <= {$unsigned({reg503[(1'h0):(1'h0)],
                      ($unsigned(reg454) ?
                          $signed((8'ha5)) : reg469[(4'hb):(1'h1)])}),
                  $signed(reg486[(3'h5):(1'h1)]),
                  reg522[(3'h5):(1'h0)]};
              reg626 = (~|($unsigned({$unsigned(reg525), (~&wire564)}) ?
                  reg460 : $signed(reg443)));
              reg627 = $unsigned(reg542);
              reg628 <= ($unsigned({reg611[(1'h0):(1'h0)],
                      $unsigned($unsigned((7'h41)))}) ?
                  ($signed({{reg456, reg457, reg500}, $unsigned(reg566)}) ?
                      $unsigned($signed((8'ha2))) : $unsigned(({reg490,
                              reg599} ?
                          $signed(reg569) : (reg486 >> reg575)))) : (8'hb3));
            end
        end
      reg629 = {((wire430 ?
                  ($signed((7'h4b)) ^~ {reg579,
                      (8'hb3),
                      reg519}) : $signed({reg447})) ?
              (!(^((8'haf) || reg608))) : reg627[(3'h5):(1'h1)]),
          reg458[(2'h2):(2'h2)],
          (((7'h56) < reg546) << (&(~|((8'hbe) ? (8'hb7) : reg546))))};
      reg630 = $unsigned((reg537[(1'h0):(1'h0)] ?
          (8'ha8) : $signed(((reg612 >= reg485) - (8'hae)))));
      for (forvar631 = (1'h0); (forvar631 < (3'h5)); forvar631 = (forvar631 + (1'h1)))
        begin
          reg632 = reg528;
          for (forvar633 = (1'h0); (forvar633 < (3'h5)); forvar633 = (forvar633 + (1'h1)))
            begin
              reg634 = ($signed(reg608[(5'h10):(4'ha)]) || {((~reg489) ?
                      $signed($signed((7'h4e))) : ($signed(reg626) > $signed((7'h40)))),
                  reg614[(1'h0):(1'h0)]});
              reg635 <= (8'ha4);
              reg636 = $signed({reg624,
                  (~^(reg585 * {reg454, reg469, (7'h55)})),
                  $signed(reg469[(1'h1):(1'h1)])});
              reg637 = ($signed(reg610) <<< $unsigned(reg589));
              reg638 = reg572[(1'h1):(1'h0)];
              reg639 <= reg516;
            end
          reg640 <= (($unsigned((~(reg628 ?
              reg549 : reg438))) ~^ ((^reg628) ^ (-$signed(reg519)))) != (!$signed($unsigned((-reg469)))));
          if (wire426)
            begin
              reg641 = ({(-(reg530 ?
                          ((8'hae) * reg600) : ((8'ha4) ? reg495 : forvar601))),
                      ((+$unsigned(reg575)) <<< ((reg624 ^~ reg443) + (~&reg623))),
                      (~reg539[(3'h5):(2'h3)])} ?
                  $unsigned(reg609[(5'h18):(5'h12)]) : $unsigned(reg438[(3'h4):(3'h4)]));
              reg642 = (~&$signed(reg463[(4'he):(3'h5)]));
              reg643 = (~|$unsigned(((reg525 ^~ reg617) ^ {{reg573}, reg514})));
              reg644 = ($signed((reg497 ?
                      (~|(8'had)) : $signed((reg516 >= reg537)))) ?
                  wire426[(5'h12):(5'h10)] : forvar633[(1'h0):(1'h0)]);
            end
          else
            begin
              reg645 <= (reg615 ?
                  {(reg618[(5'h11):(2'h3)] >= ((reg620 >= reg606) ?
                          $unsigned((8'haa)) : (reg489 ? reg438 : reg450))),
                      reg549[(3'h4):(2'h2)]} : ($unsigned($signed(reg603[(3'h4):(3'h4)])) ?
                      forvar595 : (reg438 != ({reg498, (8'h9c)} ?
                          {reg605, reg525} : reg569))));
              reg646 <= {((&((reg512 ?
                          reg598 : reg520) <<< ((8'ha6) ^~ reg608))) ?
                      ((reg607 ?
                          (reg629 >> reg484) : reg645[(3'h7):(2'h2)]) <= ($unsigned(reg514) && forvar619[(2'h2):(1'h0)])) : ($signed((-reg620)) ~^ ($unsigned(reg592) < $unsigned(reg514)))),
                  {reg609[(5'h1d):(4'ha)],
                      ($unsigned(reg575) ^ (~^$signed(reg549))),
                      $signed(((|(7'h52)) ?
                          $unsigned(reg608) : reg493[(4'h8):(4'h8)]))},
                  $signed(($unsigned((wire428 >> reg460)) == $unsigned(reg599)))};
              reg647 = reg558[(1'h0):(1'h0)];
              reg648 = ((^~reg605[(3'h4):(2'h2)]) ^ $signed(reg572));
              reg649 <= $signed(reg489[(2'h2):(2'h2)]);
              reg650 <= reg562;
              reg651 <= (~{reg614});
            end
          reg652 = ({(|(((8'hb4) ? reg558 : reg607) ?
                      $signed((8'hb3)) : (reg454 ? reg467 : reg506))),
                  ($unsigned((wire430 - reg495)) ?
                      reg515 : $signed((reg510 ^~ reg640)))} ?
              reg609[(5'h19):(5'h12)] : $signed(reg589));
        end
    end
  always
    @(posedge clk) begin
      for (forvar653 = (1'h0); (forvar653 < (3'h4)); forvar653 = (forvar653 + (1'h1)))
        begin
          reg654 <= (!$unsigned($signed(($unsigned(reg551) <<< reg645[(3'h5):(2'h2)]))));
        end
      reg655 <= {reg649};
      reg656 = (reg438[(1'h1):(1'h0)] ?
          (-$signed(reg620)) : reg586[(5'h19):(3'h6)]);
      reg657 = reg519[(4'hd):(3'h7)];
      for (forvar658 = (1'h0); (forvar658 < (2'h3)); forvar658 = (forvar658 + (1'h1)))
        begin
          for (forvar659 = (1'h0); (forvar659 < (2'h3)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 = reg456[(1'h0):(1'h0)];
              reg661 <= $unsigned(reg605);
              reg662 <= reg645[(3'h7):(3'h7)];
              reg663 = reg443[(3'h4):(1'h0)];
            end
          reg664 <= ($unsigned($unsigned({forvar659,
                  $unsigned(reg607),
                  (7'h56)})) ?
              reg522 : (-($unsigned((reg552 != (8'ha6))) ?
                  reg514[(1'h0):(1'h0)] : $unsigned({reg511,
                      (8'hba),
                      reg657}))));
          reg665 = wire428;
          if (reg586)
            begin
              reg666 <= ((+reg463) + $signed(($unsigned($unsigned(reg605)) ~^ $unsigned((forvar658 ?
                  wire425 : forvar659)))));
              reg667 <= reg463[(5'h1a):(3'h7)];
              reg668 = ($unsigned((($unsigned(reg620) ?
                      (reg615 >= reg450) : wire431[(5'h15):(4'hc)]) ?
                  reg651[(1'h1):(1'h0)] : reg579[(1'h0):(1'h0)])) ~^ $unsigned({(8'hb1),
                  ($unsigned(reg645) * $unsigned(reg585)),
                  $unsigned((reg654 != wire428))}));
            end
          else
            begin
              reg666 <= $signed((reg489 >> $unsigned((reg611 ?
                  reg558[(1'h1):(1'h1)] : ((8'ha4) ? reg558 : reg437)))));
              reg667 <= (~^$signed((7'h41)));
            end
          reg669 = $signed($signed($signed($unsigned(forvar659))));
        end
    end
  assign wire670 = ((|reg503[(2'h3):(2'h3)]) ?
                       ($unsigned({reg506,
                           (wire430 ? reg500 : reg571),
                           $unsigned(reg469)}) <<< $signed((((8'h9c) && reg500) == $unsigned(reg434)))) : (reg616 ?
                           (^((reg558 || wire426) << wire594[(3'h7):(3'h5)])) : reg620));
  always
    @(posedge clk) begin
      for (forvar671 = (1'h0); (forvar671 < (2'h2)); forvar671 = (forvar671 + (1'h1)))
        begin
          reg672 <= ($signed((((reg506 ? reg611 : reg654) ?
                  reg598[(3'h7):(3'h5)] : (~^(7'h53))) && reg651[(5'h19):(5'h14)])) ?
              (^reg586) : (|$signed(($signed(reg500) ?
                  wire430 : reg552[(4'ha):(2'h2)]))));
          reg673 = reg667[(3'h5):(1'h1)];
          for (forvar674 = (1'h0); (forvar674 < (3'h6)); forvar674 = (forvar674 + (1'h1)))
            begin
              reg675 <= reg439[(4'hd):(3'h5)];
              reg676 <= ((-(7'h4a)) ? reg606 : (!{$signed($signed(reg467))}));
              reg677 = {reg603, (~reg575[(3'h6):(3'h5)])};
            end
        end
    end
  assign wire678 = (reg514 <= reg562[(3'h6):(3'h4)]);
  always
    @(posedge clk) begin
      if (((^{(!$unsigned(reg539)),
              $signed($unsigned(reg490)),
              ((^reg516) ? $signed((8'hbe)) : {reg585})}) ?
          (+(((reg607 ? reg579 : reg645) ?
                  reg640[(4'hc):(4'hb)] : (reg530 << (8'haa))) ?
              $signed($signed(reg433)) : (&reg439[(5'h11):(4'hc)]))) : (~&(8'hb4))))
        begin
          reg679 = {(reg605 ?
                  $unsigned((!(reg463 ?
                      (8'hb1) : (8'h9f)))) : $signed(($signed(reg640) <<< (+reg485)))),
              ((^reg438) ^~ {$unsigned(reg460[(2'h2):(2'h2)])})};
          for (forvar680 = (1'h0); (forvar680 < (3'h5)); forvar680 = (forvar680 + (1'h1)))
            begin
              reg681 = $signed($signed(((8'hb1) || (+(^~wire426)))));
              reg682 <= (($signed(reg433) > (({reg519, reg558} ?
                  $signed(reg664) : (reg586 != reg500)) >= (~^(reg493 < (7'h4b))))) >> $unsigned((~($unsigned(reg552) >= {reg498,
                  reg466,
                  reg635}))));
              reg683 = (&reg490[(1'h1):(1'h1)]);
            end
        end
      else
        begin
          for (forvar679 = (1'h0); (forvar679 < (2'h2)); forvar679 = (forvar679 + (1'h1)))
            begin
              reg680 = $unsigned((7'h50));
              reg682 <= (^reg645[(3'h4):(1'h0)]);
              reg683 = (|(!(reg460[(4'ha):(4'h8)] ?
                  reg679[(4'hc):(3'h7)] : ((reg485 || forvar680) > reg640[(4'hb):(3'h6)]))));
              reg684 <= reg651;
              reg685 = (~&$unsigned((!reg672)));
              reg686 = (7'h4b);
            end
          reg687 = (((reg649[(1'h0):(1'h0)] ?
                  ($signed((7'h49)) << {reg666, (7'h55), wire564}) : (8'hba)) ?
              {{(-reg467), reg611},
                  (~&(~|reg683))} : $signed(reg529)) >>> ((~&$signed((reg625 <<< reg613))) ~^ ($unsigned(wire670[(2'h2):(2'h2)]) ?
              ($signed(reg437) == (~&reg605)) : $signed(reg611))));
          reg688 <= (^~reg442[(3'h4):(3'h4)]);
          reg689 = reg654;
          reg690 <= (reg511 * $signed(reg433));
          if ((((($signed(reg598) ? (reg466 <<< (8'had)) : reg607) ?
                  $unsigned($unsigned(reg503)) : (+reg542[(1'h1):(1'h0)])) ?
              (~&{((8'ha1) ? reg506 : wire426),
                  $signed(reg450)}) : $unsigned((reg596[(5'h14):(4'hc)] > $signed(reg543)))) | (((-$signed((8'haf))) <= (8'hb7)) >= $unsigned(reg500))))
            begin
              reg691 <= reg528;
              reg692 = $unsigned(reg552[(4'he):(4'he)]);
              reg693 <= reg529;
              reg694 = reg466[(3'h6):(3'h6)];
            end
          else
            begin
              reg691 <= (~|(8'ha7));
              reg692 = reg522[(3'h7):(3'h6)];
              reg694 = reg572;
              reg695 <= reg442[(1'h0):(1'h0)];
              reg696 = reg645;
              reg697 = $signed(reg498[(4'he):(2'h3)]);
              reg698 <= wire425;
            end
        end
      reg699 <= $unsigned((((~^reg495[(4'h8):(4'h8)]) ?
          reg467[(4'hd):(3'h5)] : {(reg439 ? (8'hb5) : reg519),
              (reg454 ? reg434 : reg506),
              reg662[(4'h9):(3'h5)]}) && ($unsigned($signed(reg498)) & (((8'ha8) ^~ reg490) ~^ (reg585 ?
          reg562 : reg551)))));
      reg700 <= (8'hb6);
      for (forvar701 = (1'h0); (forvar701 < (3'h6)); forvar701 = (forvar701 + (1'h1)))
        begin
          if ($unsigned(reg528))
            begin
              reg702 <= reg640[(1'h0):(1'h0)];
              reg703 <= $signed(($unsigned(($unsigned(reg655) ?
                  $signed(reg539) : (~|reg454))) <= $unsigned(reg525)));
              reg704 = reg585[(4'hc):(4'hb)];
              reg705 = {(reg696[(2'h3):(1'h0)] ? forvar680 : reg539),
                  $signed($unsigned($signed(reg516))),
                  (-(reg466 + (((8'haa) > reg680) * reg699[(3'h5):(1'h1)])))};
              reg706 <= reg498;
              reg707 <= $unsigned((($unsigned(reg650) < ((~|reg522) & reg699)) << ((~^$signed(reg615)) ?
                  (((8'hbc) || reg433) * reg511[(1'h1):(1'h1)]) : (+reg685[(2'h2):(1'h1)]))));
              reg708 = $signed(((reg484[(2'h2):(1'h0)] | {(reg528 ?
                      reg662 : (8'ha3)),
                  {reg696}}) ^~ reg598[(4'h8):(2'h3)]));
            end
          else
            begin
              reg702 <= $unsigned(($signed((reg516 >> (8'hbf))) << $unsigned(($unsigned(reg703) != (^~wire594)))));
              reg704 = reg645;
              reg705 = reg585;
              reg706 <= $unsigned(reg569[(4'h8):(4'h8)]);
              reg707 <= (^reg549[(4'hd):(3'h5)]);
              reg709 <= (+(reg592 || $signed(reg691)));
            end
          for (forvar710 = (1'h0); (forvar710 < (2'h2)); forvar710 = (forvar710 + (1'h1)))
            begin
              reg711 = $unsigned((~|({(wire431 ?
                      reg606 : reg442)} != ((~|(8'hb9)) ?
                  (wire678 & reg537) : {reg447}))));
            end
          reg712 <= ($signed(reg596[(1'h1):(1'h1)]) ?
              {{$unsigned((forvar710 ? reg685 : reg434))},
                  $signed({(!reg585),
                      $unsigned(reg650),
                      (reg575 ? reg529 : reg546)}),
                  reg551} : (+($signed((reg693 >> reg606)) ?
                  (|reg687) : ($unsigned(reg433) ~^ $signed(reg458)))));
          for (forvar713 = (1'h0); (forvar713 < (2'h2)); forvar713 = (forvar713 + (1'h1)))
            begin
              reg714 <= $unsigned(((($unsigned(reg454) ?
                          ((7'h47) != reg569) : $signed(reg646)) ?
                      (reg611[(1'h0):(1'h0)] ^~ $unsigned(reg514)) : ($signed(reg605) ?
                          reg662[(1'h0):(1'h0)] : $unsigned((7'h50)))) ?
                  (-reg438) : (reg709[(2'h2):(1'h1)] >> $unsigned(reg460[(3'h4):(2'h3)]))));
              reg715 = reg542;
              reg716 = ((($unsigned((~|reg672)) ?
                  (~^reg530[(5'h10):(1'h1)]) : (reg455[(4'he):(4'hc)] ?
                      $unsigned(reg579) : $signed(reg682))) ^~ (((reg635 < reg490) ?
                  (reg599 > reg543) : (&reg558)) >>> (+(reg437 ^ wire594)))) ^~ reg645);
              reg717 <= {{(reg552[(3'h5):(3'h5)] ?
                          reg709[(5'h12):(4'hd)] : {reg606[(3'h4):(1'h0)],
                              reg433[(3'h4):(1'h1)]}),
                      (~|(^reg604)),
                      ($unsigned($signed(reg530)) ?
                          reg467[(3'h4):(2'h3)] : reg684)}};
            end
          for (forvar718 = (1'h0); (forvar718 < (2'h3)); forvar718 = (forvar718 + (1'h1)))
            begin
              reg719 <= reg692[(1'h1):(1'h0)];
              reg720 = (~^$unsigned((^~reg503[(2'h3):(2'h2)])));
              reg721 <= ($signed(reg698[(5'h13):(4'he)]) >> ($signed($unsigned($signed(reg664))) <<< $unsigned(reg680)));
            end
          for (forvar722 = (1'h0); (forvar722 < (2'h2)); forvar722 = (forvar722 + (1'h1)))
            begin
              reg723 <= (reg586 <= $unsigned($unsigned((7'h4a))));
              reg724 = ({$signed(($unsigned(forvar701) ?
                      (reg569 >>> (8'h9d)) : (!reg672))),
                  $signed($unsigned((reg662 | (7'h50)))),
                  $unsigned(reg438)} | (~$signed(reg685)));
              reg725 = $unsigned((+(~&reg696[(2'h2):(1'h1)])));
              reg726 <= ((((8'hb6) ?
                      $unsigned(reg512) : wire564[(1'h1):(1'h0)]) > reg515[(1'h1):(1'h0)]) ?
                  {((^$signed(reg598)) ? reg721 : reg706[(1'h0):(1'h0)]),
                      (!({reg516, (8'hbb), (8'hb5)} ?
                          $signed(reg676) : (reg696 & reg485)))} : $signed(reg712[(4'ha):(2'h2)]));
              reg727 <= $signed(({reg605,
                      ($signed(reg562) ? {(8'hbe), (7'h49)} : (~|wire425))} ?
                  (~^(^~(reg684 ^ reg706))) : reg681));
            end
        end
      reg728 <= (($signed($unsigned((7'h47))) >> $unsigned($signed($signed(reg661)))) == $unsigned($signed(($signed(reg457) || (reg662 ?
          reg620 : reg571)))));
      if ((((forvar679 ? $signed(reg607[(2'h3):(2'h3)]) : (~(~^wire426))) ?
              $signed(reg625[(1'h0):(1'h0)]) : reg694) ?
          (|((reg604[(4'h8):(3'h6)] ? (7'h4a) : {reg646, reg680}) ?
              (-(reg522 ?
                  reg705 : reg460)) : reg549)) : $unsigned($unsigned({(forvar701 ?
                  reg573 : wire430)}))))
        begin
          for (forvar729 = (1'h0); (forvar729 < (3'h6)); forvar729 = (forvar729 + (1'h1)))
            begin
              reg730 <= reg666[(4'he):(4'h8)];
              reg731 = (($signed(reg572[(3'h4):(2'h2)]) <<< reg434) <= ({$signed(reg486),
                  (reg434[(1'h0):(1'h0)] ? (|reg528) : {wire425})} && reg442));
              reg732 <= $unsigned($signed(reg466));
              reg733 = ((($unsigned(reg613[(4'h8):(2'h2)]) ?
                      $unsigned(reg457[(4'hc):(2'h3)]) : $unsigned((^~(8'hbb)))) & $signed($signed(reg539[(3'h6):(3'h5)]))) ?
                  ((reg439 <= $signed((~|reg715))) ?
                      ($signed((reg546 < reg539)) ?
                          $signed((reg454 ?
                              reg667 : reg463)) : ((reg691 ~^ forvar710) ?
                              (reg709 || reg456) : $unsigned((7'h57)))) : (!reg514[(1'h1):(1'h1)])) : reg679[(5'h15):(4'hb)]);
              reg734 <= $signed(reg506);
              reg735 <= reg728;
            end
          if (((+$unsigned((~&$signed(reg562)))) >>> {{reg586}}))
            begin
              reg736 = (!(!reg434[(4'hf):(4'hf)]));
              reg737 = ((7'h51) ?
                  $unsigned($unsigned($unsigned({reg522}))) : $signed(reg649[(2'h3):(1'h1)]));
              reg738 = forvar718[(1'h0):(1'h0)];
              reg739 = (($signed(({reg569} * (reg456 ?
                  reg585 : reg706))) == (~$signed({reg719}))) ^~ (-$unsigned(((reg522 >> reg467) + $signed(reg542)))));
            end
          else
            begin
              reg740 <= ({reg539,
                      $unsigned({$unsigned(reg683)}),
                      $unsigned(reg724)} ?
                  wire426 : ((reg719 & reg490[(1'h0):(1'h0)]) ?
                      $signed(wire427[(1'h1):(1'h0)]) : ($unsigned($signed(reg661)) ~^ forvar729)));
              reg741 = reg708[(3'h4):(1'h1)];
              reg742 <= $signed(reg628[(2'h2):(1'h0)]);
              reg743 <= ($signed({$signed($signed(reg485))}) * reg717);
            end
          for (forvar744 = (1'h0); (forvar744 < (3'h5)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 = $signed({((reg733 ?
                      (reg500 ?
                          reg667 : reg681) : (~|reg463)) ~^ (^~$signed(reg683))),
                  $signed(($unsigned((8'hab)) ?
                      reg566 : reg437[(3'h4):(3'h4)]))});
            end
          reg746 <= (+(~^reg739[(1'h0):(1'h0)]));
          reg747 <= {(+(^~(((7'h45) << reg539) ?
                  $signed(forvar744) : {reg640, wire678}))),
              (reg551[(3'h6):(3'h6)] ?
                  (+((-reg458) ^ (reg469 - reg709))) : $signed((~|$signed(reg447))))};
          reg748 <= reg549;
        end
      else
        begin
          reg729 = $unsigned(reg457);
          reg730 <= (reg690[(2'h3):(1'h0)] >>> reg438);
          reg731 = {reg635};
          if ((~^(reg520[(1'h0):(1'h0)] ?
              (~reg728) : (($unsigned(reg712) ?
                  (8'h9e) : reg442[(4'ha):(3'h5)]) >= $unsigned((reg675 < reg697))))))
            begin
              reg732 <= $signed($signed(reg628[(5'h12):(4'ha)]));
              reg733 = (reg747 ?
                  (+$signed($signed($unsigned(reg489)))) : reg732[(4'he):(4'he)]);
            end
          else
            begin
              reg732 <= (reg506[(4'hf):(4'he)] != ($unsigned(reg662[(2'h3):(1'h1)]) || ((reg484[(4'h8):(3'h5)] ^ (reg651 ?
                  (8'ha1) : (7'h57))) >>> $unsigned(reg500[(1'h0):(1'h0)]))));
              reg733 = ((8'hbf) < $unsigned(reg579));
              reg736 = $signed($unsigned(reg579));
              reg740 <= reg698;
            end
          if (reg702[(3'h5):(1'h1)])
            begin
              reg741 = $unsigned(reg699[(2'h3):(1'h0)]);
              reg742 <= (((reg720[(5'h15):(5'h15)] ?
                      $signed($unsigned(reg645)) : ((~^(7'h4a)) ?
                          (7'h48) : (~^reg727))) ?
                  reg711 : reg696) ^~ reg490[(2'h3):(2'h2)]);
              reg744 = reg666;
              reg745 = (!(8'hb5));
              reg749 = $signed(($signed(($unsigned(reg598) > (reg666 ^~ reg469))) ^ (~&((reg728 && wire429) ?
                  reg737 : $signed(reg615)))));
              reg750 <= (reg613[(3'h6):(2'h2)] ?
                  $unsigned(($unsigned((reg708 <= reg447)) ^~ $unsigned(reg720))) : $signed($signed((~|$signed(reg705)))));
            end
          else
            begin
              reg741 = reg708[(2'h3):(2'h2)];
              reg742 <= $signed((~{reg717[(4'h8):(1'h0)],
                  (^(reg562 > (7'h47)))}));
              reg744 = reg528;
            end
          reg751 = $signed($signed(reg687[(5'h14):(4'hf)]));
          reg752 = $unsigned(wire564[(2'h3):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      reg753 <= (|reg730);
      reg754 = {$signed({({reg512, reg709, reg700} ?
                  (reg485 ^~ (7'h40)) : (reg676 | reg599)),
              ((reg490 ? reg645 : reg546) ? (~^reg703) : reg707)}),
          (|((^reg721[(1'h0):(1'h0)]) ?
              (^~(!reg458)) : $signed(((8'h9e) ~^ (8'h9d)))))};
      reg755 <= ((wire426 ?
              (!((reg549 ? reg747 : reg529) ?
                  (reg628 >> reg497) : (reg695 ?
                      reg695 : reg489))) : ((|reg740) ? reg549 : (7'h41))) ?
          ($signed(reg740[(2'h2):(2'h2)]) + $signed($unsigned(reg655[(1'h1):(1'h0)]))) : $unsigned($unsigned((^~(reg558 <<< reg572)))));
      for (forvar756 = (1'h0); (forvar756 < (1'h1)); forvar756 = (forvar756 + (1'h1)))
        begin
          for (forvar757 = (1'h0); (forvar757 < (2'h3)); forvar757 = (forvar757 + (1'h1)))
            begin
              reg758 = $signed(reg458);
              reg759 = $unsigned((8'ha2));
              reg760 <= {($signed(reg498[(3'h7):(2'h2)]) != (((reg520 ^ reg528) | ((7'h50) | reg562)) ?
                      (&$signed(reg433)) : {$unsigned((8'hbe)), (~|reg664)}))};
              reg761 = reg434;
              reg762 = $signed($unsigned((~|(^~{reg699, reg514}))));
              reg763 = reg605[(4'h8):(3'h5)];
            end
          for (forvar764 = (1'h0); (forvar764 < (3'h6)); forvar764 = (forvar764 + (1'h1)))
            begin
              reg765 = $unsigned(reg546);
              reg766 <= $unsigned(($signed($signed($signed(wire428))) ?
                  reg572[(4'he):(4'hb)] : reg539[(4'hc):(3'h4)]));
              reg767 = $signed((|reg761));
              reg768 <= ($unsigned(reg613) ~^ $signed({$signed((!reg717)),
                  $signed(((7'h4a) ? reg586 : reg549)),
                  ((~^reg506) ? $unsigned(reg561) : reg450)}));
              reg769 = reg562;
              reg770 = $signed((~&(~reg543)));
              reg771 <= (reg616[(1'h1):(1'h1)] ?
                  (reg522 >>> ({$signed(forvar757),
                          (reg443 ? reg743 : reg542),
                          $unsigned(reg537)} ?
                      $unsigned($signed(reg605)) : ($signed(reg439) > (~^reg730)))) : (reg635 ^~ reg693));
            end
          for (forvar772 = (1'h0); (forvar772 < (1'h0)); forvar772 = (forvar772 + (1'h1)))
            begin
              reg773 = (((reg493[(5'h14):(4'ha)] ?
                  ((reg469 ? reg511 : reg645) ?
                      (reg522 ?
                          reg712 : wire670) : reg746) : forvar756) >>> reg719[(2'h2):(1'h0)]) >> reg551[(4'ha):(1'h0)]);
              reg774 = (~{(7'h58)});
              reg775 = {(reg447[(3'h4):(1'h1)] ^ $unsigned(($signed(reg707) ?
                      (reg607 ? reg743 : reg520) : wire425[(1'h0):(1'h0)])))};
            end
          reg776 <= {(({(reg734 >= (8'hba))} || (((7'h4a) < reg458) ?
                  (7'h46) : (reg458 ? reg682 : reg506))) >> reg562)};
          reg777 <= reg573[(4'ha):(2'h3)];
        end
      reg778 = $signed($unsigned(reg703[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      for (forvar779 = (1'h0); (forvar779 < (3'h6)); forvar779 = (forvar779 + (1'h1)))
        begin
          reg780 <= $signed((~^(reg646 ? $signed((-reg460)) : (~(~^reg651)))));
          for (forvar781 = (1'h0); (forvar781 < (3'h5)); forvar781 = (forvar781 + (1'h1)))
            begin
              reg782 <= reg702;
              reg783 <= reg655[(5'h12):(3'h6)];
              reg784 = (^($unsigned((7'h4c)) ?
                  $signed(reg606) : (~^((reg742 - forvar779) ~^ reg746[(2'h2):(2'h2)]))));
              reg785 = (7'h55);
            end
          for (forvar786 = (1'h0); (forvar786 < (2'h2)); forvar786 = (forvar786 + (1'h1)))
            begin
              reg787 <= (!$signed(((~&reg482[(3'h5):(1'h1)]) ?
                  ((~|reg703) ?
                      $unsigned((7'h53)) : (reg512 | reg691)) : (wire430 ?
                      reg702 : $signed(reg484)))));
              reg788 <= ($unsigned((-$unsigned((&(7'h49))))) * $signed($signed($unsigned($unsigned(reg603)))));
              reg789 <= $signed($signed({((^~(8'hb4)) <<< reg511[(2'h2):(1'h0)]),
                  reg606}));
              reg790 = $signed(($signed((&reg688[(2'h2):(2'h2)])) ?
                  $signed((^(reg437 ?
                      reg539 : reg717))) : (~|reg649[(4'ha):(3'h6)])));
              reg791 <= $signed((~reg484));
            end
        end
      for (forvar792 = (1'h0); (forvar792 < (3'h4)); forvar792 = (forvar792 + (1'h1)))
        begin
          reg793 = (|reg628);
          for (forvar794 = (1'h0); (forvar794 < (1'h0)); forvar794 = (forvar794 + (1'h1)))
            begin
              reg795 = $signed((~^(~^$signed((^~reg605)))));
              reg796 <= (7'h53);
            end
          reg797 <= (reg748 ?
              $unsigned((($unsigned((7'h53)) ?
                  (reg511 || reg784) : (reg467 ?
                      reg537 : (7'h52))) >>> ((~reg699) || (reg748 ?
                  reg529 : reg695)))) : $signed($unsigned($unsigned((|reg706)))));
          for (forvar798 = (1'h0); (forvar798 < (1'h1)); forvar798 = (forvar798 + (1'h1)))
            begin
              reg799 = (^(({{wire425}, $signed(reg511)} ?
                      reg575 : (((7'h53) & reg589) >>> reg529)) ?
                  (&reg575[(3'h4):(1'h0)]) : (~^(((8'ha3) ? reg457 : reg734) ?
                      (~|reg433) : ((7'h41) <<< (8'hb4))))));
            end
        end
      reg800 = ({reg529[(4'he):(1'h0)],
              ((reg780[(5'h17):(2'h2)] ^ reg528) ?
                  reg455 : reg490[(1'h0):(1'h0)]),
              ((+(+reg795)) ?
                  {forvar786[(4'hd):(4'hd)],
                      $unsigned((8'ha8))} : (!(reg543 > reg466)))} ?
          reg519 : (&($unsigned(reg664) ? {$unsigned(reg651)} : reg575)));
      reg801 = (forvar798 + reg447[(1'h1):(1'h1)]);
      for (forvar802 = (1'h0); (forvar802 < (3'h5)); forvar802 = (forvar802 + (1'h1)))
        begin
          if (wire594[(2'h3):(2'h2)])
            begin
              reg803 = $signed((((reg782[(2'h2):(1'h1)] - (reg456 ^ reg782)) ?
                      $unsigned($unsigned(reg707)) : reg717[(5'h16):(4'he)]) ?
                  (^$signed($signed(reg728))) : reg735));
              reg804 <= (&forvar798);
              reg805 <= {{reg740}, reg640[(5'h12):(5'h12)]};
              reg806 <= $unsigned((~|reg466[(2'h2):(2'h2)]));
            end
          else
            begin
              reg804 <= (~^(reg667 && reg454));
              reg807 = (8'haf);
            end
          reg808 <= (-$signed(reg734));
          reg809 <= $unsigned(reg649[(4'h8):(2'h3)]);
          for (forvar810 = (1'h0); (forvar810 < (2'h2)); forvar810 = (forvar810 + (1'h1)))
            begin
              reg811 = {$signed((~^(~|$unsigned(reg457)))),
                  $signed(($signed((reg486 <= (8'hb6))) * (~(reg613 ?
                      (8'ha5) : (7'h53)))))};
              reg812 = (reg776[(4'h9):(3'h4)] ?
                  (!(+$unsigned((reg537 - reg661)))) : (+$unsigned(forvar798[(4'hc):(4'ha)])));
              reg813 <= $signed(reg777);
            end
          reg814 <= reg732;
          reg815 = {((reg490[(2'h3):(2'h3)] ?
                  reg721[(3'h6):(3'h5)] : (8'ha9)) >>> reg788[(5'h14):(3'h7)]),
              {(($unsigned(reg688) & (reg806 ~^ reg706)) ?
                      reg561[(1'h1):(1'h0)] : ((wire425 < reg592) <<< ((8'ha8) ?
                          reg489 : reg709)))}};
        end
      if ((|($signed(($unsigned(reg709) > (reg613 ? reg795 : reg776))) ?
          $unsigned(($unsigned(reg777) <<< reg796[(1'h1):(1'h1)])) : ($signed({reg766}) & ((&reg438) * reg793)))))
        begin
          reg816 <= reg795[(4'hc):(2'h2)];
          reg817 = (&$unsigned($unsigned(reg571[(1'h0):(1'h0)])));
          reg818 = $signed(reg651[(1'h1):(1'h1)]);
          reg819 <= ((~reg558[(2'h3):(2'h3)]) ?
              {$unsigned(reg625[(4'h8):(3'h5)]),
                  ($signed(((8'haa) >> reg490)) + (reg699[(2'h3):(2'h2)] ?
                      reg817 : $unsigned(reg620))),
                  (8'haa)} : $signed((^($signed((7'h55)) ?
                  $signed(reg503) : {reg732, reg753}))));
          reg820 <= reg585[(4'hb):(4'hb)];
        end
      else
        begin
          reg817 = reg515;
          reg819 <= reg511;
          reg821 = $signed(reg490[(1'h0):(1'h0)]);
          reg822 <= (reg768 & (^{reg467,
              $signed((~&(8'h9e))),
              ($signed(reg603) ? (|reg611) : ((8'ha7) ? reg438 : reg730))}));
          for (forvar823 = (1'h0); (forvar823 < (2'h2)); forvar823 = (forvar823 + (1'h1)))
            begin
              reg824 <= $unsigned(((reg817[(1'h0):(1'h0)] <= (^~(reg820 ?
                  reg537 : reg780))) | (|$unsigned(reg456))));
              reg825 = reg520;
              reg826 = $signed($signed((~|reg506)));
              reg827 <= (-(reg746[(1'h1):(1'h1)] != $signed(reg690[(1'h1):(1'h0)])));
              reg828 = ((!{reg456}) < ((-((forvar792 ? reg655 : reg771) ?
                  $signed(reg667) : reg495[(4'he):(1'h0)])) >= $unsigned({$signed(forvar802),
                  (+reg528),
                  ((7'h57) == reg579)})));
            end
          reg829 = $unsigned({(((reg690 ? reg458 : (8'h9d)) ?
                  wire564[(3'h5):(2'h3)] : reg719[(3'h7):(2'h3)]) <<< reg611)});
          for (forvar830 = (1'h0); (forvar830 < (3'h4)); forvar830 = (forvar830 + (1'h1)))
            begin
              reg831 <= $unsigned(($unsigned(reg719[(3'h7):(3'h6)]) ?
                  (7'h56) : (!($signed(reg438) ?
                      (reg828 ? reg782 : reg466) : (reg516 != reg558)))));
              reg832 <= reg799[(2'h2):(1'h1)];
              reg833 = $unsigned({$unsigned(($signed(reg714) ?
                      $unsigned(reg620) : reg815[(5'h1c):(5'h19)]))});
              reg834 <= $unsigned($signed((&reg755[(2'h3):(2'h3)])));
              reg835 = (reg799[(4'h9):(1'h0)] > $unsigned(reg566));
            end
        end
      if (((reg825 ? reg782[(1'h0):(1'h0)] : $signed({reg829[(4'he):(4'hd)]})) ?
          $unsigned(($signed((8'hb6)) ?
              wire670 : $signed((reg585 ? reg795 : reg730)))) : (8'haa)))
        begin
          reg836 = reg625[(1'h1):(1'h1)];
          for (forvar837 = (1'h0); (forvar837 < (3'h5)); forvar837 = (forvar837 + (1'h1)))
            begin
              reg838 = $unsigned(reg572[(1'h1):(1'h1)]);
            end
          reg839 = $unsigned($unsigned(reg730));
          for (forvar840 = (1'h0); (forvar840 < (1'h0)); forvar840 = (forvar840 + (1'h1)))
            begin
              reg841 = (((reg655 ?
                  $signed($signed((7'h54))) : reg703[(5'h15):(2'h2)]) * {(-reg688),
                  forvar810,
                  reg651[(2'h3):(1'h1)]}) ^ reg746);
              reg842 = $signed((7'h49));
              reg843 = (^~reg684[(5'h12):(2'h3)]);
              reg844 = $signed((((7'h52) && reg566[(2'h3):(1'h0)]) ?
                  $unsigned((((7'h56) >>> reg698) <<< $unsigned(reg714))) : reg691[(3'h6):(1'h1)]));
            end
        end
      else
        begin
          for (forvar836 = (1'h0); (forvar836 < (2'h2)); forvar836 = (forvar836 + (1'h1)))
            begin
              reg837 = ({(~|reg833[(3'h5):(2'h2)])} <<< reg562[(4'ha):(4'h8)]);
              reg840 <= {{$unsigned($signed($unsigned(reg815))),
                      (~&((reg684 ? reg817 : reg691) ?
                          (reg454 ? reg727 : reg826) : $unsigned(reg528)))},
                  reg603};
              reg841 = (reg790[(1'h0):(1'h0)] > reg452);
              reg845 <= {((7'h41) - (~{$signed(reg780),
                      reg789[(1'h1):(1'h1)],
                      $unsigned((8'hb7))})),
                  $signed(reg784),
                  $signed(reg607[(2'h3):(1'h0)])};
            end
          reg846 = ({$signed(reg546[(4'hb):(3'h6)]),
              reg486,
              reg529[(2'h2):(1'h1)]} >= reg655[(4'h9):(1'h1)]);
          for (forvar847 = (1'h0); (forvar847 < (3'h6)); forvar847 = (forvar847 + (1'h1)))
            begin
              reg848 = (~^(((-reg539) ?
                  (-{reg463,
                      reg525,
                      (7'h43)}) : $unsigned((forvar798 - reg552))) | $unsigned(((~|reg572) & {reg469,
                  reg596,
                  reg607}))));
              reg849 <= (reg516 ?
                  $unsigned($unsigned(((!reg562) >>> (^reg433)))) : reg650[(5'h10):(4'h8)]);
              reg850 = ((~|$signed({reg450[(1'h1):(1'h1)],
                  $signed(reg750),
                  $signed((8'ha4))})) & (+{wire431[(5'h17):(4'hb)]}));
              reg851 = (reg777[(3'h5):(3'h5)] > ((8'ha2) ?
                  (^(~&(&reg585))) : $signed($unsigned(reg822[(2'h3):(1'h0)]))));
              reg852 = reg691[(5'h11):(4'hf)];
              reg853 <= reg447[(1'h1):(1'h0)];
            end
          if (($signed(reg664[(4'h8):(2'h3)]) - reg516))
            begin
              reg854 = (({reg695, {{forvar810}}} ?
                  {((forvar786 >= wire670) == reg490[(1'h0):(1'h0)]),
                      ({reg598, forvar836, reg831} ?
                          $signed(reg654) : (reg495 ?
                              forvar840 : reg835))} : reg606) == $signed(($signed($unsigned(reg748)) ?
                  {{reg816, reg542},
                      $signed(reg463)} : reg740[(3'h6):(2'h2)])));
              reg855 = reg845[(1'h1):(1'h1)];
              reg856 = ((reg495[(4'ha):(2'h2)] ?
                      reg562[(3'h4):(2'h2)] : ((forvar792[(5'h14):(3'h4)] - {reg434,
                          (7'h43)}) <<< ((reg727 | reg811) ?
                          reg740[(3'h4):(3'h4)] : reg695[(4'h8):(3'h7)]))) ?
                  (~&{(!reg717),
                      $unsigned((&wire431))}) : ((((reg551 == reg784) ^~ (8'hab)) ?
                          $signed(reg829[(5'h15):(4'h8)]) : ((reg646 ?
                                  reg522 : reg676) ?
                              {(7'h44), (7'h47), reg808} : reg820)) ?
                      ($unsigned(reg486[(1'h0):(1'h0)]) | reg589) : reg832));
            end
          else
            begin
              reg857 <= (&forvar786);
              reg858 <= (wire430 ?
                  (((~^{reg529}) ?
                      $signed($unsigned(reg460)) : {reg734[(5'h12):(5'h10)]}) >>> ($unsigned((reg558 ?
                      (8'ha5) : (7'h47))) <<< (reg836[(3'h6):(3'h4)] ?
                      ((8'hba) << reg723) : reg571))) : (^~reg442));
              reg859 = (~^forvar836);
            end
          if ($signed(((&wire594[(3'h7):(1'h0)]) ~^ forvar802[(2'h3):(2'h2)])))
            begin
              reg860 = reg469;
            end
          else
            begin
              reg860 = ($signed(reg655) ?
                  $signed((^$signed($signed(reg613)))) : reg467[(4'hb):(1'h1)]);
              reg861 <= (^(|reg639));
              reg862 = reg783;
              reg863 = reg552;
              reg864 = (^reg661);
              reg865 = $signed((($unsigned((reg755 ?
                  reg714 : reg695)) && (~&$signed((8'hb5)))) != (~^reg458)));
              reg866 <= (forvar847 ?
                  ($signed(reg635[(5'h13):(3'h4)]) ?
                      ((~&(8'had)) | ({reg460, reg796, reg442} ?
                          reg746[(1'h1):(1'h0)] : {reg865,
                              forvar847})) : $signed($unsigned((reg811 <<< wire429)))) : (reg734 ?
                      reg782[(4'h8):(2'h3)] : (!$unsigned($unsigned(reg821)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg867 = $signed(((($unsigned(reg797) ~^ $unsigned(reg849)) <= reg695) >>> $unsigned(reg734[(3'h4):(2'h2)])));
    end
  always
    @(posedge clk) begin
      reg868 <= {($unsigned(reg816[(3'h4):(1'h0)]) << $signed({$unsigned(wire426),
              {reg579, reg467}})),
          (+(&({(8'hae)} >>> reg753[(2'h3):(1'h0)]))),
          (wire428[(3'h7):(1'h1)] + (reg782 <<< (8'hb5)))};
      if ((($unsigned({$unsigned(reg832),
                  $unsigned(reg654),
                  reg732[(3'h7):(3'h5)]}) ?
              reg796[(1'h0):(1'h0)] : (!((reg858 <<< reg688) <<< (reg734 ~^ reg558)))) ?
          $unsigned(reg522[(2'h3):(2'h3)]) : reg598[(3'h5):(3'h4)]))
        begin
          reg869 = $unsigned((7'h54));
          reg870 = reg691;
          for (forvar871 = (1'h0); (forvar871 < (3'h4)); forvar871 = (forvar871 + (1'h1)))
            begin
              reg872 <= reg869[(5'h17):(3'h7)];
              reg873 = (7'h40);
              reg874 = ($signed(reg599[(4'hb):(1'h0)]) ?
                  {{$signed((7'h54))},
                      reg688[(4'h8):(2'h2)],
                      (~&$unsigned($signed(reg490)))} : $signed(($unsigned(reg503[(1'h1):(1'h0)]) != $signed($signed(reg690)))));
              reg875 <= ($signed((8'ha7)) | (8'h9f));
              reg876 = (!{(reg768 ?
                      $unsigned($signed((8'hac))) : ($signed(reg806) ?
                          {(8'ha2)} : (~|reg691))),
                  reg572});
              reg877 = {reg787,
                  ({(&reg698[(5'h12):(1'h1)])} ^~ (($signed(reg700) ?
                      $unsigned(wire594) : {reg654,
                          reg797,
                          reg866}) ~^ $signed($unsigned(reg439)))),
                  (($signed((&reg726)) == $signed((reg516 ?
                      (8'hbc) : reg442))) || {($unsigned(reg529) <= $unsigned(reg575)),
                      $signed({(8'hbc), reg566, wire429})})};
            end
        end
      else
        begin
          reg869 = $signed((reg748[(4'h9):(3'h5)] ?
              reg740[(2'h3):(1'h0)] : reg598[(3'h5):(3'h4)]));
          reg871 <= $unsigned($signed(({reg625[(4'ha):(3'h5)], (|(8'haf))} ?
              reg599[(2'h3):(1'h0)] : $signed((^~reg780)))));
          for (forvar872 = (1'h0); (forvar872 < (3'h6)); forvar872 = (forvar872 + (1'h1)))
            begin
              reg873 = ($signed((~|wire594)) ?
                  ((($unsigned(reg497) <<< $signed(reg748)) ?
                          reg814 : reg452[(2'h2):(1'h1)]) ?
                      $signed(reg562[(3'h6):(3'h5)]) : ($signed($unsigned(reg452)) ?
                          $signed((reg824 < forvar872)) : ({reg662,
                              reg858,
                              reg605} ^~ (7'h41)))) : ((7'h53) ?
                      ($unsigned((reg712 != reg813)) >>> reg760[(1'h0):(1'h0)]) : (($unsigned(reg661) == wire429) ?
                          $unsigned((8'hb1)) : (reg814[(3'h5):(2'h2)] ?
                              ((7'h51) ? (8'haa) : reg808) : {(8'haa),
                                  reg456,
                                  (7'h49)}))));
              reg875 <= (((^$unsigned({reg442})) * reg484) ?
                  {(~$unsigned((reg682 ? reg706 : reg845))),
                      $signed(($signed(reg740) | (&reg806))),
                      (~reg579)} : reg742[(4'hb):(4'h8)]);
              reg876 = (7'h58);
              reg877 = (reg748 ? reg603[(3'h5):(2'h3)] : reg834);
              reg878 <= $signed((^~$unsigned((&reg571))));
              reg879 <= reg516;
            end
        end
      reg880 <= $signed(reg676[(4'ha):(3'h6)]);
    end
  always
    @(posedge clk) begin
      for (forvar881 = (1'h0); (forvar881 < (2'h2)); forvar881 = (forvar881 + (1'h1)))
        begin
          if ({((reg645 ?
                      (reg484 ?
                          (~&reg603) : (reg661 ?
                              wire564 : (7'h41))) : $unsigned((|(7'h47)))) ?
                  $signed(reg490[(1'h0):(1'h0)]) : (reg707[(2'h3):(2'h2)] ^ reg806)),
              reg433})
            begin
              reg882 <= reg743;
              reg883 <= $signed({reg528, $signed($unsigned((8'hb6)))});
              reg884 <= forvar881[(1'h0):(1'h0)];
            end
          else
            begin
              reg885 = reg510;
              reg886 <= ($unsigned(reg640) | ({reg579[(1'h0):(1'h0)],
                      $unsigned((reg520 | reg639)),
                      (~reg490)} ?
                  reg530 : {{$unsigned(reg791), {reg546, reg740}},
                      ($signed(reg747) ^ reg661[(5'h15):(4'h8)])}));
            end
          for (forvar887 = (1'h0); (forvar887 < (3'h4)); forvar887 = (forvar887 + (1'h1)))
            begin
              reg888 = reg695;
              reg889 = reg805;
            end
          if (reg572)
            begin
              reg890 = $unsigned((~($signed($unsigned(reg655)) + ($unsigned((8'haf)) ?
                  reg611[(2'h3):(1'h1)] : $unsigned(reg503)))));
              reg891 = reg592[(3'h4):(2'h3)];
              reg892 <= ($signed(((7'h4b) ? reg884 : reg635)) < (7'h54));
              reg893 <= ($signed($signed(reg866[(3'h6):(1'h0)])) ?
                  reg458 : $unsigned((reg840 ~^ ((reg662 ? reg654 : reg714) ?
                      (^~(7'h52)) : (reg640 != reg747)))));
              reg894 = reg606[(5'h12):(4'ha)];
              reg895 = reg572;
              reg896 = {(^~$signed((forvar881 != reg662))),
                  $unsigned($unsigned((wire564[(3'h7):(2'h2)] <<< (reg546 & (8'h9c))))),
                  $signed($signed((reg489 ?
                      $unsigned((8'ha8)) : (reg732 ? reg883 : reg598))))};
            end
          else
            begin
              reg890 = (&(reg740 >= ({((7'h45) ? reg675 : (8'hb9)),
                  $signed(reg693),
                  $signed(reg740)} >> $signed(reg484[(4'ha):(2'h2)]))));
              reg892 <= $signed(((+$signed((^reg719))) ?
                  ((|(reg698 ? reg640 : reg495)) ?
                      (-(wire430 ? reg886 : reg709)) : {{(7'h56),
                              reg640,
                              reg787}}) : ((reg728[(5'h18):(5'h16)] >> (8'h9e)) - (((8'hbc) <<< reg522) < $unsigned(reg598)))));
            end
          reg897 <= ({($signed($signed(wire426)) ?
                  reg645[(1'h1):(1'h1)] : (8'ha1))} - {wire426});
        end
      if (reg552[(4'hb):(3'h4)])
        begin
          reg898 <= (^({reg672, reg443[(1'h0):(1'h0)]} ?
              (reg879 ?
                  $unsigned(reg780) : {(~^reg750)}) : $signed($signed(((7'h40) ?
                  reg789 : (8'had))))));
          reg899 <= $unsigned(reg562);
          for (forvar900 = (1'h0); (forvar900 < (2'h3)); forvar900 = (forvar900 + (1'h1)))
            begin
              reg901 = reg700;
              reg902 = $unsigned($unsigned($signed((forvar881[(1'h0):(1'h0)] * reg728))));
              reg903 <= (^(~|reg457[(1'h0):(1'h0)]));
            end
          reg904 = reg888[(4'h8):(1'h0)];
          reg905 = ($signed($signed(reg628)) ?
              ((8'h9d) * $signed(reg777)) : ({((reg816 ?
                      (7'h4b) : reg895) << $unsigned(reg500)),
                  $signed($unsigned(reg897)),
                  {(^~reg611)}} | (^$unsigned(reg723[(3'h4):(2'h2)]))));
          reg906 = reg454;
          reg907 = (7'h4b);
        end
      else
        begin
          if ($signed($signed(reg879[(3'h4):(1'h0)])))
            begin
              reg898 <= $signed((reg707[(1'h1):(1'h1)] | $unsigned((reg664 ?
                  {reg589, reg452} : {reg899}))));
              reg900 = reg650[(2'h3):(1'h0)];
              reg903 <= {reg592,
                  {(+$unsigned(reg437[(2'h3):(1'h1)])),
                      $unsigned({reg748,
                          reg895[(4'ha):(2'h3)],
                          (reg676 >>> reg490)}),
                      reg433}};
              reg904 = (($signed({$signed(reg456),
                      reg651}) ^~ (!((reg813 && (7'h41)) ?
                      (~|reg486) : (reg743 > reg698)))) ?
                  (^reg549[(4'hc):(4'h8)]) : reg896);
            end
          else
            begin
              reg898 <= ((reg635[(5'h12):(3'h5)] * $signed({(reg861 || wire430),
                  ((8'ha8) == reg485)})) <<< reg719);
              reg899 <= reg897[(1'h1):(1'h1)];
              reg900 = reg573;
            end
          reg908 <= {(^~$signed((8'hba))),
              (~&(8'ha9)),
              {(((reg596 ? reg766 : reg516) ~^ reg787) | $signed({reg782,
                      reg813,
                      reg750})),
                  (&$unsigned(wire428[(3'h7):(3'h4)]))}};
        end
      reg909 = (reg808 && $unsigned((~^$signed(reg433[(4'hc):(4'hb)]))));
      if ({reg503[(2'h3):(2'h3)], reg806})
        begin
          reg910 = reg776;
          reg911 <= reg702[(3'h4):(2'h3)];
          if (reg776[(4'h8):(3'h6)])
            begin
              reg912 <= $signed((|(-{(~|reg605), (reg676 >> reg607)})));
              reg913 = reg433[(1'h1):(1'h1)];
              reg914 <= (reg884[(3'h7):(3'h7)] != ((!$signed((~|reg510))) ?
                  reg447[(3'h4):(1'h1)] : (({reg575,
                      (8'hbe),
                      reg776} && (reg858 ? reg489 : reg743)) || reg908)));
            end
          else
            begin
              reg913 = wire427;
              reg914 <= (-$unsigned(((7'h4d) ?
                  reg484[(4'he):(4'hd)] : (reg746 ? reg522 : wire431))));
              reg915 <= $signed(((|$unsigned((reg613 & reg520))) < reg503));
              reg916 = $signed(($unsigned(reg898[(3'h5):(2'h2)]) * $signed(reg702[(4'h8):(1'h0)])));
              reg917 = (reg598[(4'h9):(3'h4)] << $signed($unsigned((8'hb9))));
            end
        end
      else
        begin
          reg910 = (^$unsigned(($unsigned(reg604[(1'h0):(1'h0)]) < reg750[(3'h5):(3'h4)])));
          for (forvar911 = (1'h0); (forvar911 < (3'h5)); forvar911 = (forvar911 + (1'h1)))
            begin
              reg912 <= (($unsigned($signed($signed(reg649))) || (((reg573 ?
                      reg572 : reg542) != reg917) ^ ((reg661 ?
                      reg904 : reg482) < $signed(reg611)))) ?
                  reg546 : (&(~|(7'h53))));
            end
          reg914 <= ($unsigned(reg707) ?
              reg734 : (+{reg460[(4'hb):(3'h4)],
                  (wire427 <<< $unsigned(reg755)),
                  reg882}));
        end
      if ((~|$signed($signed((~|(~reg755))))))
        begin
          reg918 = reg510;
          if ((~&reg886[(2'h2):(1'h0)]))
            begin
              reg919 <= reg809;
            end
          else
            begin
              reg919 <= $unsigned($signed($signed($signed(reg709[(4'hb):(1'h0)]))));
              reg920 <= ($signed($signed(((reg571 ? (7'h43) : wire564) ?
                  $signed(reg528) : (~reg717)))) ^~ (^$signed(($signed(reg569) ~^ reg894[(2'h2):(1'h0)]))));
            end
          reg921 <= wire431[(3'h5):(1'h0)];
          for (forvar922 = (1'h0); (forvar922 < (3'h6)); forvar922 = (forvar922 + (1'h1)))
            begin
              reg923 <= $signed(reg788);
              reg924 = reg827[(2'h3):(1'h0)];
              reg925 <= (~|{reg551[(2'h2):(2'h2)]});
              reg926 = (~&reg755);
              reg927 = {$signed(($unsigned((reg783 ^ reg514)) << (reg735[(4'hb):(1'h0)] | (!reg514)))),
                  (!(^((7'h52) - reg613[(1'h0):(1'h0)]))),
                  $signed(reg746[(3'h4):(2'h3)])};
            end
          reg928 <= reg666[(4'h9):(1'h1)];
          reg929 <= $signed($unsigned($unsigned({$unsigned(reg814),
              $signed(reg893),
              $unsigned(reg639)})));
          reg930 <= (($unsigned(reg561[(5'h13):(1'h0)]) | ((+{(7'h42),
                  reg907,
                  reg484}) - (8'hb1))) ?
              reg573 : $signed($unsigned(reg879[(4'h8):(3'h5)])));
        end
      else
        begin
          reg919 <= $signed($signed({((reg909 != (7'h51)) ?
                  (reg787 ? reg493 : reg495) : $signed(reg914)),
              reg579,
              (&$unsigned(reg883))}));
          if ((reg885 * $unsigned(((~|(reg452 ? reg892 : reg831)) ?
              (reg606 ?
                  reg878[(3'h7):(1'h1)] : (reg743 != reg892)) : $signed((~reg646))))))
            begin
              reg922 = (7'h54);
              reg923 <= ((+$signed($unsigned(reg928))) ?
                  forvar887[(4'hc):(4'h8)] : $signed(reg699[(2'h3):(2'h3)]));
            end
          else
            begin
              reg922 = reg434[(3'h5):(2'h2)];
            end
          reg924 = ({((8'hbe) * (8'hbe)),
                  {$signed($unsigned((7'h53))), reg787}} ?
              $signed(reg493[(3'h5):(3'h4)]) : ((~&$signed((^~forvar911))) ?
                  reg814[(3'h6):(3'h6)] : (reg804[(4'hd):(3'h5)] - $unsigned((reg691 ?
                      wire430 : reg503)))));
          for (forvar925 = (1'h0); (forvar925 < (1'h1)); forvar925 = (forvar925 + (1'h1)))
            begin
              reg926 = reg712;
              reg927 = reg796[(2'h3):(1'h0)];
            end
          reg928 <= {((((reg604 ?
                      reg871 : reg917) != $unsigned(reg599)) >>> (8'hbb)) ?
                  (~&(reg639[(2'h2):(2'h2)] & (~^reg598))) : (reg806[(1'h0):(1'h0)] ?
                      reg639[(1'h1):(1'h1)] : forvar925[(2'h2):(1'h1)])),
              reg543,
              {($unsigned({reg858, reg672}) ?
                      ($unsigned(reg666) ~^ (reg690 & reg605)) : ((reg878 ?
                          reg452 : reg466) && (reg911 ? reg776 : reg592))),
                  {reg730}}};
          reg931 = $signed(reg699[(1'h0):(1'h0)]);
          reg932 <= (^~$signed(reg889));
        end
      for (forvar933 = (1'h0); (forvar933 < (2'h3)); forvar933 = (forvar933 + (1'h1)))
        begin
          if ($unsigned(reg808[(4'ha):(1'h1)]))
            begin
              reg934 <= $unsigned((($signed(reg805) ?
                  (!wire670[(1'h0):(1'h0)]) : $unsigned((reg598 + reg447))) <<< $unsigned($signed({reg605,
                  reg905,
                  (7'h46)}))));
              reg935 <= (~|($unsigned(reg905) >>> $signed($signed((-reg776)))));
              reg936 = (^~reg537[(4'hd):(4'hd)]);
              reg937 = reg552;
              reg938 = (+(~&$signed((|reg519[(4'hd):(3'h6)]))));
              reg939 = ({reg539} <= reg805[(2'h3):(1'h0)]);
            end
          else
            begin
              reg934 <= (reg888 ? reg460[(5'h12):(5'h12)] : reg907);
              reg936 = $signed($signed({(reg809[(5'h1e):(5'h14)] != $signed(reg732)),
                  $signed((|reg497))}));
              reg940 <= ((reg937 ?
                      reg640[(5'h1c):(3'h5)] : (~($unsigned((7'h53)) ?
                          $signed(reg495) : $signed((8'hbe))))) ?
                  (((8'hae) < $unsigned((reg904 & (7'h55)))) <= $signed(({reg649,
                          reg905,
                          reg675} ?
                      $signed(reg586) : (reg768 ? reg493 : reg529)))) : reg709);
              reg941 = reg804;
            end
          reg942 <= reg926[(3'h4):(2'h3)];
          reg943 = (~reg437);
          reg944 <= reg768;
        end
      reg945 = (reg539[(1'h0):(1'h0)] ?
          (~^reg813) : $signed(reg721[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg946 = $signed(reg929[(5'h19):(4'hc)]);
      for (forvar947 = (1'h0); (forvar947 < (1'h1)); forvar947 = (forvar947 + (1'h1)))
        begin
          for (forvar948 = (1'h0); (forvar948 < (2'h2)); forvar948 = (forvar948 + (1'h1)))
            begin
              reg949 <= $unsigned(wire425);
              reg950 = (~&reg771[(4'h8):(3'h7)]);
              reg951 = (reg940[(5'h14):(3'h6)] >= $signed({((reg878 ?
                          reg452 : reg434) ?
                      (+reg585) : (reg510 >> reg911)),
                  {$unsigned(reg522)},
                  $signed(reg520[(2'h2):(1'h0)])}));
              reg952 <= reg797;
              reg953 = $signed(wire427);
              reg954 <= (~&reg651[(3'h5):(1'h1)]);
            end
          reg955 = (reg777[(1'h1):(1'h0)] < reg940);
          for (forvar956 = (1'h0); (forvar956 < (1'h1)); forvar956 = (forvar956 + (1'h1)))
            begin
              reg957 <= $unsigned(reg651);
              reg958 <= reg592;
              reg959 = (|reg592);
              reg960 <= $signed(reg695);
              reg961 = reg434;
              reg962 <= ((reg666[(2'h2):(2'h2)] ?
                      $signed({$signed(reg514), reg820}) : (^(8'hb3))) ?
                  ((({reg959, reg706, reg709} ?
                      (!reg649) : (reg908 ?
                          reg558 : reg562)) <= {(^~reg892)}) < (&reg616[(1'h1):(1'h0)])) : $unsigned($signed(reg897[(5'h17):(4'ha)])));
            end
          reg963 <= (reg892 ?
              reg814 : {$signed(($unsigned(reg935) ?
                      (reg789 || reg960) : (~^reg450))),
                  $unsigned(reg598[(2'h2):(2'h2)]),
                  reg727[(4'h8):(3'h6)]});
        end
      reg964 <= $signed({(8'h9d),
          ((~|reg562) ?
              $unsigned($unsigned(reg788)) : $signed(reg457[(4'hc):(4'hc)]))});
    end
  always
    @(posedge clk) begin
      reg965 = $signed($signed(($unsigned($signed((8'had))) << $signed(reg814[(4'hb):(2'h3)]))));
      reg966 <= reg586[(5'h15):(5'h12)];
      for (forvar967 = (1'h0); (forvar967 < (3'h4)); forvar967 = (forvar967 + (1'h1)))
        begin
          reg968 = reg664;
          reg969 = (^((~^({reg727, reg824, reg575} ?
                  wire427[(1'h0):(1'h0)] : (~|wire429))) ?
              ($unsigned((reg730 ?
                  reg721 : reg562)) << (^{reg615})) : (~|(^~$signed(reg942)))));
          if (((~|$unsigned($unsigned(reg664))) ?
              ((((reg460 ? reg928 : reg675) >>> (reg666 ?
                      reg776 : reg768)) ^~ $signed((reg698 >> reg439))) ?
                  reg620[(4'hb):(4'hb)] : {(((8'hb6) ~^ reg857) ?
                          (reg498 ? reg558 : reg604) : (~&(7'h4a))),
                      reg447,
                      reg911[(2'h2):(1'h1)]}) : reg525[(3'h7):(1'h1)]))
            begin
              reg970 = $unsigned((reg944 ^~ reg482[(3'h5):(1'h0)]));
            end
          else
            begin
              reg971 <= ($signed(($unsigned({reg898, reg942}) ?
                  $unsigned(reg882) : $unsigned($unsigned(reg712)))) != {reg893[(1'h0):(1'h0)],
                  $signed(((&(8'hba)) ?
                      ((7'h48) ? reg845 : reg490) : (&wire670))),
                  reg592[(3'h5):(3'h5)]});
              reg972 <= reg650;
              reg973 = (((&(&reg923)) ?
                  reg934 : (~&((8'ha7) ?
                      (reg573 | reg579) : (reg667 && reg552)))) << ((reg645[(2'h3):(1'h1)] ?
                      ($signed(reg880) <= {reg930, reg969, reg615}) : (reg703 ?
                          (^reg964) : ((8'ha9) ? reg819 : reg897))) ?
                  reg748[(2'h2):(1'h1)] : $unsigned(($signed((8'ha3)) ?
                      reg603[(4'ha):(4'ha)] : $signed(wire429)))));
              reg974 <= ({(((reg820 ^ reg868) ?
                              {reg726, (8'ha2)} : (~|reg721)) ?
                          (~(reg503 ?
                              reg768 : reg520)) : reg861[(5'h10):(4'hc)]),
                      {(-((8'hbd) ? reg969 : reg858)),
                          $signed((|wire678)),
                          $signed((reg857 ? reg537 : reg952))}} ?
                  {reg512, reg972} : (($signed(reg489[(2'h3):(2'h2)]) ?
                          reg969[(3'h7):(3'h6)] : reg672) ?
                      (~^reg690) : reg586));
              reg975 = ({(($signed((7'h46)) ?
                              $unsigned(reg789) : reg450[(2'h2):(2'h2)]) ?
                          reg746 : $unsigned((8'ha0))),
                      reg482,
                      $unsigned((reg853 ?
                          $signed(reg469) : (reg886 ? (8'haf) : reg651)))} ?
                  reg607[(3'h4):(1'h1)] : reg734);
              reg976 = reg439[(3'h4):(2'h2)];
            end
          if (($signed($signed(reg899)) ?
              reg571[(2'h2):(2'h2)] : {(reg516[(4'he):(1'h0)] ?
                      $signed((reg934 <= reg753)) : $signed((^(8'ha9)))),
                  (-(^(reg882 ? reg976 : reg589)))}))
            begin
              reg977 = reg975;
              reg978 <= (7'h57);
              reg979 <= reg872[(5'h1a):(4'hc)];
              reg980 = $signed($signed(reg952));
              reg981 = reg569;
            end
          else
            begin
              reg977 = (($signed($signed((^reg871))) | $unsigned(reg675[(4'ha):(1'h1)])) <= {reg639,
                  $unsigned($signed($signed(reg455)))});
              reg978 <= $signed(((7'h55) * (((wire427 || reg857) >> $unsigned((8'hab))) * ($unsigned(reg966) >= (reg957 ?
                  reg820 : reg954)))));
              reg980 = ((~^reg964) + reg438);
              reg982 <= wire678;
              reg983 <= (~|{$signed((reg693 ? {reg783} : $signed(reg561))),
                  {((reg519 ? (7'h4d) : reg727) ?
                          reg871[(4'ha):(4'h9)] : reg605)},
                  $unsigned($signed($unsigned((7'h48))))});
              reg984 = (reg780 > reg727[(4'he):(3'h4)]);
            end
          for (forvar985 = (1'h0); (forvar985 < (2'h3)); forvar985 = (forvar985 + (1'h1)))
            begin
              reg986 = ($unsigned(($signed($unsigned(reg966)) ?
                  reg979[(3'h6):(2'h2)] : $unsigned($signed(reg734)))) + $unsigned(reg437[(2'h3):(2'h3)]));
            end
          for (forvar987 = (1'h0); (forvar987 < (2'h3)); forvar987 = (forvar987 + (1'h1)))
            begin
              reg988 = (reg966[(2'h3):(2'h2)] ^~ {(&((+forvar985) ?
                      reg919[(4'hd):(3'h6)] : (reg454 ? reg791 : reg983)))});
            end
        end
      if ((reg782[(4'h9):(4'h9)] + $unsigned((^~reg882[(1'h0):(1'h0)]))))
        begin
          reg989 <= {{(~|($signed((7'h41)) || reg845))},
              reg573,
              (!reg923[(4'h9):(1'h1)])};
          reg990 <= reg666[(2'h3):(2'h2)];
          if ((!(^~(($unsigned(reg971) ? (wire430 * (8'hb1)) : reg522) ?
              reg455 : ($signed(reg853) ?
                  reg512[(5'h10):(2'h3)] : {(7'h44), reg662, reg514})))))
            begin
              reg991 = ((({reg510, reg734, (8'hb0)} ?
                      $unsigned((reg714 ? reg962 : reg771)) : $signed((reg463 ?
                          reg734 : reg599))) >> (^((reg654 - (8'hbe)) ?
                      reg768[(2'h3):(2'h2)] : (reg447 ^ reg964)))) ?
                  $unsigned((|reg575)) : (^~$unsigned($signed($signed(reg571)))));
              reg992 <= forvar967[(4'hb):(3'h6)];
            end
          else
            begin
              reg991 = $signed(reg746[(3'h4):(2'h2)]);
              reg993 = reg605;
              reg994 = $signed(({reg964[(3'h5):(3'h5)],
                  reg925[(5'h14):(1'h1)]} <<< $signed($signed($signed(reg788)))));
              reg995 <= (-$signed((~&$unsigned($unsigned(reg840)))));
            end
          reg996 <= wire564[(3'h6):(2'h2)];
          reg997 = {reg655[(4'hc):(4'ha)],
              reg573,
              {($signed($signed(reg728)) ?
                      $unsigned($signed(wire678)) : reg734[(2'h2):(1'h0)])}};
        end
      else
        begin
          for (forvar989 = (1'h0); (forvar989 < (3'h4)); forvar989 = (forvar989 + (1'h1)))
            begin
              reg990 <= (7'h4b);
              reg992 <= (reg930[(4'h9):(3'h4)] ?
                  reg919 : (|(^reg969[(4'hc):(3'h6)])));
              reg995 <= (~^{{$unsigned((~|reg598)),
                      reg966[(3'h4):(3'h4)],
                      $unsigned(reg466[(4'ha):(4'ha)])},
                  $unsigned($unsigned({reg861, reg503}))});
              reg997 = reg442[(2'h3):(2'h2)];
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg750)
        begin
          reg998 = $unsigned(reg930[(2'h3):(1'h1)]);
          if ($unsigned(((reg728 ?
                  (reg607[(1'h0):(1'h0)] ?
                      reg771 : ((7'h55) || (8'hb7))) : ($unsigned(reg721) ?
                      (7'h55) : $signed(reg768))) ?
              reg920[(4'hd):(1'h1)] : (8'hbb))))
            begin
              reg999 = reg542;
              reg1000 = reg791;
            end
          else
            begin
              reg1001 <= {((($unsigned(reg682) ?
                      (&reg639) : reg463) <<< reg603) | reg734)};
              reg1002 = reg561[(5'h1b):(4'hc)];
              reg1003 = ((reg486[(5'h11):(4'ha)] >= $unsigned(($unsigned(reg712) ?
                  reg646 : (reg433 & reg942)))) * $unsigned($unsigned(($unsigned(reg522) ?
                  (reg706 ? wire429 : reg503) : $unsigned(reg649)))));
              reg1004 = {(~|reg546[(2'h2):(2'h2)]),
                  ($unsigned((~^(reg972 ? wire670 : (8'hbe)))) ?
                      (reg782[(2'h3):(1'h0)] ?
                          (reg734 <= reg695[(4'ha):(1'h0)]) : (&(+reg996))) : $signed({reg845,
                          ((7'h47) ? reg849 : (7'h4e))}))};
              reg1005 <= reg726;
            end
          for (forvar1006 = (1'h0); (forvar1006 < (2'h2)); forvar1006 = (forvar1006 + (1'h1)))
            begin
              reg1007 <= $signed({reg899});
            end
          for (forvar1008 = (1'h0); (forvar1008 < (1'h1)); forvar1008 = (forvar1008 + (1'h1)))
            begin
              reg1009 = reg816;
              reg1010 = {(~|reg579)};
              reg1011 = {$unsigned(reg437[(2'h3):(1'h1)]),
                  $unsigned($unsigned(($unsigned(reg978) ?
                      $signed(reg845) : $unsigned(reg1002)))),
                  (~&$unsigned($signed(reg992)))};
              reg1012 <= (~&reg982);
            end
        end
      else
        begin
          reg1001 <= ((reg688[(3'h6):(3'h5)] ?
              (8'hb4) : reg861[(5'h11):(2'h2)]) ^~ $signed($unsigned($signed($signed(reg983)))));
          reg1005 <= ((({$unsigned((7'h4b)),
                      (reg746 == reg452)} <= $signed((8'hb5))) ?
                  $signed((^reg620[(4'h9):(1'h1)])) : (~^$unsigned((reg978 ?
                      reg983 : reg611)))) ?
              reg561 : reg989[(5'h18):(4'hf)]);
          for (forvar1006 = (1'h0); (forvar1006 < (1'h1)); forvar1006 = (forvar1006 + (1'h1)))
            begin
              reg1007 <= (((~|(reg463[(5'h11):(5'h10)] + ((8'h9e) ?
                          reg808 : reg1007))) ?
                      {($signed(reg450) ?
                              (7'h56) : reg661[(4'hb):(4'h8)])} : ((~^wire564) >> $unsigned(reg458))) ?
                  $unsigned({$unsigned($signed(reg952))}) : ((!reg514) ?
                      $signed($unsigned($signed(reg443))) : $unsigned((~^$signed(reg709)))));
              reg1008 <= ($unsigned((|((~^reg558) ?
                  (reg858 <<< reg699) : $unsigned(reg551)))) >= ($signed((|reg458[(4'ha):(1'h1)])) | ($unsigned($signed(reg983)) ?
                  $signed($signed(reg808)) : forvar1008[(5'h13):(1'h1)])));
              reg1012 <= wire594[(2'h2):(2'h2)];
              reg1013 = reg998[(5'h10):(3'h5)];
              reg1014 = reg586[(4'hb):(1'h0)];
              reg1015 = $unsigned((+$unsigned($unsigned($unsigned(reg972)))));
            end
          reg1016 <= $unsigned($unsigned(((8'hb0) ?
              reg776 : (((7'h40) < reg861) <<< (reg831 ? reg434 : (7'h41))))));
          for (forvar1017 = (1'h0); (forvar1017 < (1'h0)); forvar1017 = (forvar1017 + (1'h1)))
            begin
              reg1018 <= $signed(reg992[(3'h7):(1'h0)]);
              reg1019 <= reg883;
              reg1020 = $signed(reg998);
              reg1021 <= {(^reg992[(5'h12):(2'h2)]),
                  ((reg616[(1'h1):(1'h1)] != {{reg974, reg519, reg662},
                      (reg655 * reg721),
                      reg662}) && (|(reg551[(3'h6):(1'h1)] <= (reg944 ?
                      reg585 : reg796))))};
              reg1022 <= $unsigned(({{reg875, (reg840 != reg771)},
                      (~|(~|reg439)),
                      reg1019} ?
                  reg735 : $unsigned($signed({reg899}))));
            end
          if ((reg684[(4'h9):(4'h8)] >>> reg735))
            begin
              reg1023 <= reg971[(2'h2):(1'h1)];
            end
          else
            begin
              reg1024 = reg437[(3'h4):(1'h1)];
              reg1025 <= $unsigned((8'h9f));
            end
          for (forvar1026 = (1'h0); (forvar1026 < (1'h0)); forvar1026 = (forvar1026 + (1'h1)))
            begin
              reg1027 <= (reg511[(1'h0):(1'h0)] ?
                  reg911[(1'h1):(1'h0)] : (~&reg966));
            end
        end
      reg1028 = $unsigned(((^(~^(reg511 ?
          reg964 : reg640))) ^ $unsigned(wire670[(1'h0):(1'h0)])));
      if ((|(^reg649[(4'ha):(4'ha)])))
        begin
          for (forvar1029 = (1'h0); (forvar1029 < (3'h4)); forvar1029 = (forvar1029 + (1'h1)))
            begin
              reg1030 = (((8'hb4) >= ($signed(reg1000) ?
                      reg963 : ((^(7'h51)) ?
                          (reg1027 >> reg511) : reg915[(5'h16):(4'hf)]))) ?
                  reg484[(3'h4):(3'h4)] : reg806);
              reg1031 = (reg1014 ?
                  ($signed((~&reg589[(1'h1):(1'h0)])) && reg808[(3'h4):(2'h3)]) : reg463[(4'he):(2'h2)]);
              reg1032 <= ((^~{(~$unsigned((8'hbe))),
                      {$signed(reg897)},
                      $unsigned((reg573 >= reg928))}) ?
                  reg551[(4'h9):(1'h1)] : (reg999 ^~ (~|reg646)));
              reg1033 = wire430;
            end
          reg1034 = $unsigned((($signed((reg599 ?
                  reg515 : reg886)) >= ((wire428 ?
                  reg832 : reg1005) ^~ {(8'haa)})) ?
              reg434[(1'h0):(1'h0)] : $unsigned(reg949)));
        end
      else
        begin
          if ((&($signed((^~$signed(reg958))) << (+((reg992 ?
              reg753 : reg1021) || reg691[(3'h4):(1'h0)])))))
            begin
              reg1029 <= reg747[(5'h10):(4'h9)];
              reg1030 = (~$signed(wire670[(2'h2):(1'h0)]));
              reg1032 <= (reg957 ?
                  (7'h4c) : {(8'hbb),
                      $signed(((reg1009 ?
                          reg832 : reg546) == ((8'hbb) * reg603)))});
              reg1035 <= reg999;
              reg1036 <= $unsigned({(|((7'h46) <<< (reg1000 > reg551)))});
              reg1037 <= ($unsigned((reg805[(1'h1):(1'h0)] * (~&(~&(8'ha2))))) ?
                  ($unsigned(({reg628, reg484} ^~ (~&reg824))) ?
                      {$unsigned((reg592 ?
                              reg1001 : reg516))} : $unsigned((reg598[(3'h5):(2'h3)] <<< $unsigned(reg1015)))) : ($unsigned((reg562 ?
                          reg957 : {reg655, reg824})) ?
                      {$unsigned($unsigned(reg878)),
                          reg1003,
                          reg796} : $signed((8'hbb))));
              reg1038 = $signed(((~&(!$signed((8'hb0)))) != $signed($signed({reg834}))));
            end
          else
            begin
              reg1030 = $unsigned(reg966[(3'h5):(1'h0)]);
              reg1032 <= (&(reg528[(1'h1):(1'h1)] ?
                  ($signed($signed(reg551)) < reg972[(5'h10):(4'hc)]) : reg791[(1'h0):(1'h0)]));
              reg1035 <= reg667;
              reg1036 <= (reg482[(3'h6):(1'h1)] ?
                  reg606[(3'h4):(2'h2)] : ($unsigned($signed($signed(reg966))) || (($unsigned(reg675) * reg726[(5'h10):(5'h10)]) > reg747[(3'h5):(3'h5)])));
              reg1038 = reg925;
            end
          if ((^reg1038[(4'h9):(3'h5)]))
            begin
              reg1039 <= (&(reg1011 ?
                  (^$unsigned(reg497[(1'h1):(1'h0)])) : reg640[(4'h8):(2'h2)]));
              reg1040 = reg651;
              reg1041 <= reg912;
              reg1042 = (($signed({(7'h4e)}) ?
                  reg651 : (reg558 ?
                      ((reg1023 ?
                          reg628 : (7'h4a)) <<< reg693[(2'h2):(2'h2)]) : (~|reg606[(5'h14):(3'h5)]))) > reg1002);
              reg1043 = $unsigned($unsigned({reg727[(3'h4):(2'h2)]}));
              reg1044 = reg490;
              reg1045 = (|((({reg827} ?
                      (reg783 ? (7'h57) : (8'ha1)) : $unsigned(reg514)) ?
                  ((reg934 ?
                      reg528 : reg688) + (reg880 ^ (8'haa))) : $unsigned((reg920 ?
                      (7'h4c) : reg814))) >> $unsigned($unsigned(reg732[(4'hb):(4'h9)]))));
            end
          else
            begin
              reg1040 = $unsigned(reg814);
              reg1042 = reg746;
            end
          reg1046 = $signed($signed({$signed((^reg719)),
              ($unsigned(reg816) <<< reg1044[(4'ha):(2'h2)])}));
          reg1047 <= {$unsigned(({{reg914},
                  $signed(reg789),
                  reg1036} <= reg645))};
          if ({(reg571[(3'h4):(1'h0)] ?
                  reg849[(5'h1a):(3'h4)] : $unsigned(reg1012))})
            begin
              reg1048 <= (~{$signed($signed($signed(reg899))),
                  $signed((reg740[(3'h5):(1'h1)] ^~ (reg960 ?
                      reg789 : reg645)))});
              reg1049 <= (((-(7'h42)) ?
                      (reg592[(4'hb):(4'h8)] != reg999) : {$signed($signed((8'hb0))),
                          (reg1003 ? reg620 : $unsigned(reg514))}) ?
                  reg820 : (((~(reg500 << (8'h9d))) & $unsigned(reg898)) >= $signed(reg635[(5'h16):(5'h14)])));
              reg1050 <= {(((reg878 ?
                      {reg442,
                          forvar1026,
                          reg484} : (reg625 - (8'ha1))) < $signed($unsigned(reg486))) & (reg808[(2'h2):(2'h2)] | reg809[(4'hb):(2'h2)])),
                  reg805,
                  {($signed((reg543 ? reg495 : (7'h57))) ?
                          reg510[(2'h2):(1'h1)] : reg512),
                      reg804}};
              reg1051 = (^(^~(-reg486)));
            end
          else
            begin
              reg1048 <= $unsigned($signed($signed((reg635 ?
                  $unsigned(forvar1006) : $signed(reg974)))));
              reg1051 = $unsigned(reg1014[(2'h2):(2'h2)]);
              reg1052 = (~$signed(((~$unsigned(reg1045)) <<< {(reg709 == reg730)})));
              reg1053 <= reg893[(2'h3):(2'h3)];
              reg1054 <= $unsigned(reg529);
              reg1055 = (~|((+{$signed(reg628),
                  (~|(7'h45)),
                  (reg1001 ~^ reg928)}) <<< $unsigned((~&$unsigned(wire428)))));
            end
        end
      reg1056 <= $signed(((|((reg806 > (7'h4a)) > reg571[(2'h3):(1'h0)])) <= ((+(^reg809)) ?
          reg1020[(4'hc):(1'h1)] : $unsigned($signed(reg1018)))));
      if (($signed(reg868[(4'he):(2'h2)]) << (~^($unsigned({reg661}) <= reg777))))
        begin
          reg1057 <= reg1021;
          for (forvar1058 = (1'h0); (forvar1058 < (3'h4)); forvar1058 = (forvar1058 + (1'h1)))
            begin
              reg1059 = $signed(reg662);
              reg1060 = reg1040;
            end
          for (forvar1061 = (1'h0); (forvar1061 < (2'h2)); forvar1061 = (forvar1061 + (1'h1)))
            begin
              reg1062 <= ($signed(reg503) ?
                  $unsigned(reg971[(1'h1):(1'h1)]) : (~(&(8'h9f))));
              reg1063 <= reg1057;
              reg1064 = reg484[(4'hc):(2'h2)];
            end
          for (forvar1065 = (1'h0); (forvar1065 < (2'h3)); forvar1065 = (forvar1065 + (1'h1)))
            begin
              reg1066 = (|({{(reg676 * reg875), (|(7'h43))},
                      (+reg912[(3'h5):(1'h1)]),
                      reg495[(1'h0):(1'h0)]} ?
                  $signed($signed(reg1033)) : ({(reg1048 ? reg915 : reg1037)} ?
                      $unsigned((reg551 ? reg485 : reg1005)) : reg721)));
              reg1067 <= $unsigned((^~reg748));
              reg1068 = (reg460[(2'h2):(2'h2)] ?
                  $unsigned((reg978 ?
                      ((reg721 > reg824) + reg1012[(5'h13):(1'h1)]) : $signed((^~reg1048)))) : reg979[(4'h8):(1'h0)]);
              reg1069 <= (~$signed($unsigned((7'h42))));
              reg1070 = ($signed(reg783) ?
                  $unsigned(reg490[(1'h0):(1'h0)]) : ((-reg516[(5'h17):(3'h6)]) ?
                      (reg1018 ?
                          $signed((|reg466)) : ((^~reg433) ?
                              (reg579 * reg1051) : (reg1044 ?
                                  reg872 : reg442))) : reg690[(1'h1):(1'h1)]));
              reg1071 = $signed($signed(reg515));
            end
          reg1072 <= reg861[(3'h6):(2'h2)];
        end
      else
        begin
          for (forvar1057 = (1'h0); (forvar1057 < (2'h3)); forvar1057 = (forvar1057 + (1'h1)))
            begin
              reg1058 = {reg1057};
              reg1059 = ($unsigned(reg635) ?
                  {(!(7'h47))} : (((&reg579[(5'h11):(4'h8)]) | ((~reg886) ?
                          $signed(reg831) : (forvar1058 ? reg592 : reg1000))) ?
                      {reg1043[(3'h7):(3'h5)],
                          (-{reg809}),
                          (((8'hae) != reg646) > {reg789,
                              reg693,
                              reg506})} : ($signed((reg516 ~^ reg1042)) ?
                          reg783 : reg849)));
            end
          for (forvar1060 = (1'h0); (forvar1060 < (2'h2)); forvar1060 = (forvar1060 + (1'h1)))
            begin
              reg1061 = $unsigned((reg930[(1'h1):(1'h0)] ?
                  reg528 : $signed({(reg579 ? (8'h9d) : reg978)})));
              reg1064 = reg930[(3'h5):(3'h5)];
              reg1065 <= {{reg797}};
              reg1067 <= reg748;
              reg1069 <= reg458[(3'h6):(3'h6)];
              reg1070 = reg628;
            end
          if ((~&$unsigned((reg914 == ((-reg813) == (reg974 ?
              reg706 : (8'ha2)))))))
            begin
              reg1071 = {reg1003, reg651[(1'h1):(1'h0)], reg734[(3'h6):(3'h5)]};
              reg1072 <= $unsigned($signed((((reg1048 - reg666) ?
                      $unsigned(reg897) : reg1000[(1'h0):(1'h0)]) ?
                  (~|reg819[(3'h7):(3'h6)]) : ($signed(reg572) <= (reg485 && reg497)))));
              reg1073 = reg463;
              reg1074 <= {reg693, reg1052[(4'ha):(2'h3)]};
              reg1075 <= {reg853[(3'h4):(1'h1)]};
              reg1076 <= ($signed({$signed(((8'ha7) <<< reg929))}) ?
                  $unsigned(wire678) : reg820);
              reg1077 <= reg832[(4'hd):(3'h4)];
            end
          else
            begin
              reg1071 = $unsigned(reg1001[(4'ha):(1'h1)]);
              reg1073 = reg949;
              reg1078 = (&{{(&reg932),
                      ((+reg1036) >= (^reg932)),
                      (^~(reg603 ? wire431 : reg1036))},
                  ((reg611 ? $unsigned(reg732) : ((8'ha0) ? reg808 : (7'h51))) ?
                      (-$signed(reg1054)) : (&(+(8'hb3)))),
                  ({(reg857 ? (8'hb2) : reg868),
                          reg717[(3'h4):(3'h4)],
                          $unsigned(reg525)} ?
                      (forvar1008 & $signed(reg537)) : ((reg469 || reg455) ?
                          $signed((8'ha7)) : $unsigned((7'h54))))});
            end
        end
      for (forvar1079 = (1'h0); (forvar1079 < (1'h1)); forvar1079 = (forvar1079 + (1'h1)))
        begin
          if (($signed(({(wire678 << reg1001)} + $signed({reg819}))) ?
              ($signed(reg672) ?
                  $signed(reg691[(4'he):(1'h0)]) : $signed((7'h45))) : reg1075[(2'h2):(2'h2)]))
            begin
              reg1080 = (((^$unsigned((reg1057 ?
                      forvar1017 : (7'h57)))) == (-reg892)) ?
                  (&reg1019[(3'h7):(3'h4)]) : ($signed(((reg562 && reg992) ?
                      reg688[(4'ha):(1'h1)] : (reg884 ?
                          reg463 : reg806))) != {(|{reg486})}));
              reg1081 = reg983[(5'h10):(5'h10)];
              reg1082 = reg1024[(1'h1):(1'h1)];
              reg1083 <= (((~{{reg928}}) ?
                      reg611[(3'h5):(2'h2)] : (reg515 ?
                          {{reg706, (7'h40), reg766},
                              (reg1057 ? reg482 : reg782),
                              reg1050} : reg780[(5'h1b):(4'ha)])) ?
                  (^~{reg666[(1'h1):(1'h1)]}) : $unsigned({$signed(reg750[(1'h0):(1'h0)])}));
              reg1084 <= (~(($unsigned(reg819[(1'h1):(1'h1)]) * ((~reg897) ~^ reg703)) ?
                  reg824 : {(8'hab),
                      ($unsigned(reg613) != $unsigned(forvar1079))}));
              reg1085 <= reg746[(3'h6):(1'h0)];
              reg1086 = $unsigned(($signed({(reg512 ?
                      reg1022 : reg990)}) * ((~(reg1035 ? reg1056 : reg702)) ?
                  $signed($signed(reg834)) : ($signed(reg1007) ?
                      {reg539, reg755} : (~&forvar1029)))));
            end
          else
            begin
              reg1080 = reg662;
            end
          if ($unsigned({$signed({(7'h50), (reg706 ? (7'h56) : reg552)})}))
            begin
              reg1087 <= reg598;
            end
          else
            begin
              reg1087 <= $unsigned(($signed({$signed(reg872),
                  reg787[(3'h4):(2'h3)],
                  (~|reg514)}) >> (~&$signed((~reg954)))));
              reg1088 <= reg460[(3'h4):(2'h3)];
            end
        end
    end
  assign wire1089 = ((^~reg515[(1'h1):(1'h0)]) ?
                        reg511[(1'h1):(1'h0)] : $unsigned(reg940[(2'h3):(2'h3)]));
  always
    @(posedge clk) begin
      for (forvar1090 = (1'h0); (forvar1090 < (3'h6)); forvar1090 = (forvar1090 + (1'h1)))
        begin
          for (forvar1091 = (1'h0); (forvar1091 < (3'h4)); forvar1091 = (forvar1091 + (1'h1)))
            begin
              reg1092 = ((!(((^~(7'h4c)) >> (wire678 || reg753)) ?
                  reg797[(4'ha):(2'h3)] : $unsigned({reg1016,
                      reg469}))) - $signed(reg1076[(3'h5):(3'h4)]));
            end
          if (reg495[(2'h3):(1'h0)])
            begin
              reg1093 <= ({$signed((~|((8'ha1) ? reg921 : reg1085))),
                      (^$signed(wire594[(1'h0):(1'h0)])),
                      $signed($unsigned({reg872, reg522}))} ?
                  $signed(($unsigned(reg732) ?
                      (reg1001 >= $unsigned(reg1037)) : (reg726[(3'h6):(1'h1)] ?
                          (8'hab) : $signed(reg742)))) : reg1057[(2'h2):(1'h1)]);
              reg1094 <= $unsigned($signed((((reg934 * reg1032) ?
                  $unsigned(reg516) : reg1065) >> $signed(((8'ha4) ?
                  reg519 : (7'h42))))));
              reg1095 <= (-(reg561[(5'h18):(2'h2)] ?
                  $signed(((~reg897) > reg530[(3'h7):(3'h7)])) : $unsigned(((&reg880) ?
                      reg512[(3'h4):(1'h1)] : $signed(reg1029)))));
              reg1096 <= reg693;
              reg1097 <= (($signed($unsigned($unsigned(reg589))) == ($signed({(8'h9d)}) ?
                  $unsigned(wire427) : ((7'h52) ?
                      reg616[(1'h1):(1'h0)] : {(7'h58),
                          (8'hbb)}))) <<< {reg1056[(4'hb):(3'h7)],
                  reg719[(1'h0):(1'h0)]});
            end
          else
            begin
              reg1098 = (-(~&$signed((-(^~reg1084)))));
              reg1099 <= ($unsigned((-($signed(reg966) >>> $signed((7'h4f))))) ?
                  $unsigned($unsigned((^~reg1075))) : (&(((reg1016 ?
                          (8'hb7) : reg546) ?
                      $signed((8'hbc)) : (^(8'ha3))) >> ((reg940 >= reg592) ?
                      $signed((8'ha1)) : reg605[(4'h8):(1'h0)]))));
              reg1100 <= reg822[(3'h7):(3'h4)];
              reg1101 = $signed({reg579[(5'h11):(4'hb)]});
              reg1102 <= reg1035;
              reg1103 <= $signed({$signed(reg899),
                  ($unsigned((reg1083 ? reg872 : reg515)) ?
                      $signed((!reg1097)) : ((reg460 | reg723) ?
                          reg703[(5'h12):(1'h1)] : {reg661, reg1077})),
                  (|((~|reg1001) >> {reg592}))});
            end
          for (forvar1104 = (1'h0); (forvar1104 < (2'h3)); forvar1104 = (forvar1104 + (1'h1)))
            begin
              reg1105 = reg966[(3'h6):(1'h0)];
              reg1106 <= reg1085[(5'h13):(5'h10)];
              reg1107 = {reg766, reg746};
              reg1108 <= ($signed((reg598[(2'h2):(1'h0)] - (reg543[(3'h7):(1'h1)] ^ $unsigned(reg766)))) ?
                  (($unsigned({reg868,
                      reg646,
                      reg1022}) - $unsigned(reg469[(5'h16):(5'h11)])) <= $unsigned((|{(7'h54)}))) : (~^$signed((7'h4b))));
              reg1109 = (^$signed((^($signed(reg768) ^ (reg748 >= wire678)))));
              reg1110 = ({($unsigned({wire429}) <<< reg575[(3'h5):(3'h5)])} ^~ {reg690});
            end
          if ($unsigned(($unsigned(({(8'h9e)} ?
              (~|reg438) : (~|reg1065))) >>> reg1097[(3'h4):(1'h0)])))
            begin
              reg1111 = (~^$unsigned($unsigned(wire427)));
              reg1112 = ($signed(reg699) ~^ reg882);
              reg1113 <= ($signed(reg730) ?
                  {reg857,
                      ($signed({reg599, reg1035, reg460}) != ((reg942 ?
                              reg586 : reg1023) ?
                          (|reg1095) : (reg546 ? reg562 : reg503))),
                      reg489[(4'h9):(4'h9)]} : $signed((&$unsigned(reg849[(3'h4):(1'h1)]))));
              reg1114 <= $signed({$unsigned(reg1057), reg516[(4'hc):(2'h2)]});
              reg1115 = (reg915 ?
                  reg586[(5'h1a):(5'h12)] : $signed($unsigned(((7'h50) ?
                      (&reg437) : reg903[(2'h3):(2'h3)]))));
              reg1116 = $signed({$unsigned($unsigned((8'hac)))});
              reg1117 <= reg1032[(3'h5):(2'h3)];
            end
          else
            begin
              reg1113 <= reg1023;
              reg1114 <= {(reg439 - {reg1025[(1'h0):(1'h0)]})};
              reg1115 = reg957[(1'h0):(1'h0)];
              reg1116 = (~|$unsigned($signed(reg878[(1'h1):(1'h1)])));
              reg1118 = $unsigned({(reg816 ?
                      {(reg561 >> (7'h47)),
                          (reg561 || reg760),
                          $signed((7'h56))} : $unsigned((reg530 ?
                          (7'h46) : (8'hb2))))});
              reg1119 <= ($signed((reg484[(4'hb):(3'h7)] + ((reg827 ?
                      reg493 : reg616) - reg549))) ?
                  (reg616 ?
                      reg646 : (|reg746)) : ($signed(reg433) - (reg655[(5'h11):(5'h10)] ^ {(8'ha9),
                      reg912})));
              reg1120 <= $signed((~&reg750[(3'h4):(2'h2)]));
            end
          reg1121 = reg875;
          reg1122 = $signed($unsigned((^$signed(reg806[(3'h4):(2'h3)]))));
          reg1123 <= ($signed($unsigned(($signed(reg996) * $unsigned(reg646)))) | reg787[(1'h1):(1'h1)]);
        end
      reg1124 = ((~^({reg463,
              (reg748 ? reg454 : reg952)} & ($signed(reg897) | reg776))) ?
          reg620[(4'hc):(1'h1)] : $unsigned((^($unsigned((7'h58)) ?
              (reg912 ? (8'hb0) : (8'hb1)) : reg925))));
      reg1125 = $signed(((~&{$unsigned(reg1048)}) ?
          ($unsigned((-reg604)) ?
              wire428[(2'h3):(1'h0)] : $signed($signed(reg511))) : reg1100));
    end
  always
    @(posedge clk) begin
      reg1126 <= (|reg566[(4'h9):(2'h2)]);
      reg1127 = (reg747[(5'h13):(3'h6)] - $unsigned(reg898[(1'h1):(1'h1)]));
      if (((reg1123[(5'h15):(4'hd)] ?
          $unsigned((~(7'h55))) : (-{(^~reg750),
              $unsigned(reg871)})) < (&reg1008)))
        begin
          reg1128 = $unsigned($signed($unsigned({(reg886 ? reg982 : reg728),
              reg861})));
          reg1129 <= (reg579[(4'hb):(4'hb)] ?
              ({$unsigned((+reg596)), (|reg500)} ?
                  (((reg604 + (7'h58)) != $signed(reg520)) ?
                      (((7'h47) ?
                          reg883 : reg1094) << $signed(reg599)) : (reg605 ?
                          $unsigned(reg452) : reg460[(3'h7):(2'h3)])) : (-reg995)) : reg606[(2'h3):(1'h0)]);
          reg1130 = (!{(7'h4f)});
          for (forvar1131 = (1'h0); (forvar1131 < (3'h6)); forvar1131 = (forvar1131 + (1'h1)))
            begin
              reg1132 = (|reg1099);
              reg1133 = (8'hbb);
              reg1134 <= (!$unsigned((|reg912[(2'h2):(2'h2)])));
              reg1135 = $unsigned({$signed((reg455 ?
                      $signed((8'hae)) : (|reg693))),
                  (|(&(~&reg589))),
                  reg834[(4'hf):(2'h2)]});
              reg1136 = reg1056;
              reg1137 <= ($unsigned((~^({reg750,
                  (8'hab)} > reg442[(2'h2):(2'h2)]))) - $unsigned((reg433 << $unsigned((reg912 ?
                  reg457 : reg747)))));
            end
          reg1138 <= $unsigned($signed(reg566));
        end
      else
        begin
          reg1129 <= reg1008;
          for (forvar1130 = (1'h0); (forvar1130 < (3'h4)); forvar1130 = (forvar1130 + (1'h1)))
            begin
              reg1131 <= ((7'h43) <= ($unsigned($signed((8'ha2))) - $signed(reg740)));
              reg1134 <= reg995[(4'he):(3'h6)];
              reg1137 <= reg740;
              reg1139 = reg886;
              reg1140 = (8'h9e);
              reg1141 = (&reg707[(1'h1):(1'h1)]);
            end
          if ((((7'h42) ? reg1041 : (8'hbb)) == reg706[(4'hb):(3'h6)]))
            begin
              reg1142 <= (~|($signed(reg746[(3'h6):(3'h4)]) >> reg728[(5'h18):(4'hf)]));
              reg1143 = ((~($signed(reg1057[(1'h1):(1'h0)]) < reg768[(2'h3):(2'h2)])) > $unsigned($signed((^$unsigned((8'h9e))))));
              reg1144 <= (~|reg455);
              reg1145 = (({($unsigned(reg712) ?
                          (reg753 ?
                              reg872 : (7'h44)) : (wire670 ^ reg971))} ^~ {reg1037[(3'h6):(2'h2)]}) ?
                  $signed(reg529) : ($signed(({reg1077} <<< $signed(reg1117))) >= (reg1032[(4'h9):(1'h0)] * reg875)));
              reg1146 <= reg1049;
              reg1147 <= $signed(reg934);
              reg1148 <= $signed($unsigned(({$signed(reg712),
                  $unsigned(reg787),
                  (reg454 & reg450)} + $unsigned({reg822, reg1037}))));
            end
          else
            begin
              reg1142 <= {$signed($signed(((!(8'ha0)) ?
                      (~^reg575) : (~reg1023)))),
                  (reg983[(5'h12):(4'hd)] ?
                      $unsigned((reg791[(1'h1):(1'h0)] ?
                          reg457[(2'h2):(1'h1)] : {reg611,
                              reg452,
                              reg1134})) : {{$unsigned(reg721),
                              ((8'ha7) ^~ (7'h4d))},
                          ((~&reg516) ? {(7'h42), reg516} : $unsigned((8'hbc))),
                          ($unsigned(reg972) ?
                              (reg458 + (7'h57)) : $unsigned(reg957))}),
                  $signed((~|$signed($signed((8'ha5)))))};
              reg1144 <= {$unsigned($unsigned($signed((reg511 ^~ reg879))))};
              reg1145 = $signed($unsigned({reg1133, reg552}));
              reg1149 = reg958[(4'hb):(4'hb)];
              reg1150 <= ((^$unsigned(($unsigned((8'hbf)) - (-reg1012)))) > $signed({((reg915 >>> reg1008) ?
                      {wire678} : reg797),
                  $signed(reg974[(2'h3):(1'h1)])}));
              reg1151 <= wire431;
            end
          for (forvar1152 = (1'h0); (forvar1152 < (3'h5)); forvar1152 = (forvar1152 + (1'h1)))
            begin
              reg1153 = ({reg1102,
                  $signed($unsigned((reg1140 ? (8'ha1) : reg1113))),
                  {$signed(reg805[(1'h1):(1'h0)]),
                      reg827[(2'h2):(1'h1)]}} > (~&(reg1012 ?
                  (reg490[(2'h3):(1'h0)] ?
                      (reg707 & reg1076) : reg783[(3'h7):(2'h3)]) : $signed((&reg1132)))));
              reg1154 <= ({reg871,
                      ((~|(reg808 > reg486)) >> $unsigned((reg780 << reg921)))} ?
                  ((reg484[(1'h0):(1'h0)] ^ (^~(reg831 ?
                      reg485 : reg740))) < (&$unsigned(reg1041))) : ({(~^(reg1117 << reg958)),
                      reg515[(3'h6):(2'h2)]} >>> wire670));
              reg1155 <= {(~$signed(reg684)),
                  (reg1138 ?
                      reg1132 : $signed(((reg640 >= reg972) ?
                          $unsigned(reg1127) : reg949[(4'hc):(4'hb)])))};
              reg1156 = $signed((&(~^((reg1094 >> reg723) ?
                  reg604 : reg514[(2'h2):(1'h1)]))));
              reg1157 = {$unsigned((~|{(~^reg949)})),
                  $unsigned(((reg791 ? reg607 : reg485[(3'h5):(3'h5)]) ?
                      {(~|(8'hb2))} : $unsigned((~|reg788)))),
                  $signed((^reg768))};
              reg1158 = forvar1131[(4'hb):(1'h0)];
            end
          reg1159 <= reg1149[(4'hc):(4'h9)];
          reg1160 <= $unsigned(reg691);
          for (forvar1161 = (1'h0); (forvar1161 < (1'h1)); forvar1161 = (forvar1161 + (1'h1)))
            begin
              reg1162 = ($unsigned(reg1019) ?
                  ((~|reg1018) >>> $signed(((reg1012 ? (7'h4d) : reg1069) ?
                      (reg893 - reg661) : (^reg882)))) : reg1039[(4'hd):(3'h5)]);
              reg1163 = $unsigned($signed($signed(({reg971} ?
                  $signed(reg605) : reg929))));
              reg1164 <= reg903[(4'hc):(3'h7)];
              reg1165 = ((~&(&$unsigned(reg511[(2'h2):(2'h2)]))) ?
                  reg519[(3'h5):(2'h3)] : $unsigned(reg438[(2'h3):(1'h0)]));
              reg1166 = {$unsigned(reg635[(4'he):(4'h8)]),
                  $signed({{{reg616, reg469}, (reg1057 ? reg607 : reg760)},
                      ($signed(reg1036) > reg599),
                      ($unsigned(reg809) << (~^reg897))}),
                  reg808[(4'ha):(4'h9)]};
              reg1167 <= reg1137[(4'he):(1'h1)];
              reg1168 = ((^~$signed((&(reg834 ? reg771 : reg930)))) ?
                  (7'h50) : (~|((+(reg820 ?
                      reg1088 : reg849)) <= (reg1130 || $signed(reg482)))));
            end
        end
      reg1169 <= {(+(~|reg691)), reg899};
      if ((!reg820[(3'h7):(1'h0)]))
        begin
          reg1170 = {reg661[(2'h2):(1'h0)], reg709};
        end
      else
        begin
          for (forvar1170 = (1'h0); (forvar1170 < (3'h4)); forvar1170 = (forvar1170 + (1'h1)))
            begin
              reg1171 <= (!$signed($signed(((reg1032 ?
                  wire431 : (8'had)) > reg635))));
            end
          reg1172 <= {($signed((8'ha7)) & $unsigned((^~(reg971 ~^ reg783))))};
          reg1173 = $unsigned({$unsigned({(^reg1048), reg1145}), reg872});
          reg1174 = (reg1067[(1'h0):(1'h0)] ?
              $unsigned(reg1148) : reg1094[(1'h0):(1'h0)]);
          reg1175 <= {$unsigned((((^reg666) + (~&reg791)) ?
                  {reg645[(1'h0):(1'h0)]} : (!$unsigned(reg746)))),
              (+{$unsigned((reg824 * reg605))})};
        end
      reg1176 <= {(reg485[(2'h3):(1'h0)] ? reg776[(4'hd):(3'h4)] : reg1022),
          $signed(reg525[(2'h2):(1'h1)]),
          (reg469 ?
              (wire1089[(2'h2):(1'h0)] ^~ $unsigned((reg1120 ?
                  reg605 : reg819))) : (reg460 && (((7'h42) >> reg607) << $signed((7'h44)))))};
      reg1177 <= reg813;
    end
  always
    @(posedge clk) begin
      if (reg1088[(4'hc):(4'ha)])
        begin
          reg1178 <= $unsigned(reg813);
          reg1179 <= (reg942 ?
              $unsigned((~|(-(reg1087 ?
                  reg1019 : reg963)))) : ($signed(reg1154) ?
                  reg730[(4'h9):(1'h0)] : reg768[(2'h3):(2'h2)]));
          if ($unsigned($unsigned($signed((~^(reg935 ? reg1008 : reg1096))))))
            begin
              reg1180 <= ((~reg603) >> $unsigned($signed(reg1057)));
              reg1181 <= (reg957[(3'h4):(1'h1)] ?
                  (~$signed((reg746 <= (8'ha3)))) : ($signed($unsigned((reg442 >> reg596))) >= reg935[(4'hc):(3'h4)]));
              reg1182 = reg1072[(2'h3):(2'h2)];
              reg1183 = (({(~(!reg1113)),
                  (~&reg1160[(1'h0):(1'h0)]),
                  (^reg607[(3'h4):(2'h3)])} ^ reg928[(1'h1):(1'h1)]) << (-reg845));
              reg1184 = ($unsigned(reg735[(5'h10):(3'h4)]) <<< $signed((&(!$signed(reg1126)))));
              reg1185 = ((~&(~$signed(reg982[(4'he):(4'hd)]))) ?
                  reg921 : $signed(reg1094[(2'h2):(1'h1)]));
              reg1186 <= ((reg706 ?
                  $signed(reg1179[(4'hd):(2'h3)]) : (8'ha7)) ^~ ({((reg1032 ?
                          reg962 : reg640) | reg1023[(5'h18):(1'h0)]),
                      $unsigned(reg611[(1'h0):(1'h0)]),
                      reg1039} ?
                  reg732 : {((reg819 != reg466) ~^ $signed(reg791))}));
            end
          else
            begin
              reg1180 <= reg1047[(2'h2):(2'h2)];
              reg1182 = {reg698[(2'h2):(1'h0)],
                  (reg512 != reg493[(2'h2):(2'h2)]),
                  reg1148[(5'h11):(3'h4)]};
              reg1183 = (({{reg1185[(1'h0):(1'h0)],
                      (reg599 ? reg971 : reg995),
                      reg726}} && (reg1001[(2'h3):(2'h3)] <<< reg551)) <<< $unsigned((reg1054 ?
                  (reg469 << $signed(reg871)) : $unsigned((reg1148 != reg707)))));
              reg1184 = reg490;
              reg1186 <= reg543[(5'h13):(4'h9)];
              reg1187 <= $signed(((~^({reg849,
                  reg1012,
                  reg747} >= $signed(reg551))) * reg561));
            end
        end
      else
        begin
          reg1178 <= {(~^reg662[(4'ha):(2'h2)])};
          for (forvar1179 = (1'h0); (forvar1179 < (2'h3)); forvar1179 = (forvar1179 + (1'h1)))
            begin
              reg1182 = (&$signed(($signed($signed(reg466)) ?
                  reg882 : $signed(((8'hb3) > reg707)))));
              reg1183 = $unsigned($unsigned({(8'hba),
                  (reg911[(3'h6):(1'h0)] ? (8'hae) : reg486[(4'h8):(4'h8)])}));
              reg1184 = reg1106;
              reg1185 = reg543;
              reg1188 = ($unsigned((&reg776[(4'h9):(4'h9)])) ?
                  reg458[(3'h6):(1'h0)] : reg1037[(3'h6):(1'h0)]);
            end
          for (forvar1189 = (1'h0); (forvar1189 < (3'h4)); forvar1189 = (forvar1189 + (1'h1)))
            begin
              reg1190 <= (!(($signed((reg1181 < reg954)) << (^$signed((8'ha7)))) ?
                  ((~^reg1048[(4'hc):(3'h7)]) || reg771) : (reg1126 ?
                      reg921 : (~{reg1095, reg1032, reg1056}))));
              reg1191 <= (^~(reg1001[(4'he):(1'h0)] ^~ (+$signed(reg589[(4'h8):(1'h0)]))));
              reg1192 = reg1164[(5'h13):(4'he)];
              reg1193 = $unsigned(reg672[(3'h6):(3'h5)]);
              reg1194 <= reg853[(3'h5):(3'h4)];
            end
          reg1195 = ({$unsigned($unsigned((reg952 ?
                  reg1047 : wire426)))} || reg1155[(3'h6):(3'h5)]);
          reg1196 = $signed(reg1114);
        end
      for (forvar1197 = (1'h0); (forvar1197 < (2'h2)); forvar1197 = (forvar1197 + (1'h1)))
        begin
          reg1198 = (reg514[(2'h2):(2'h2)] ?
              reg437 : (-$unsigned(({reg919,
                  reg827,
                  (7'h53)} >>> $signed(reg990)))));
        end
      for (forvar1199 = (1'h0); (forvar1199 < (3'h4)); forvar1199 = (forvar1199 + (1'h1)))
        begin
          reg1200 <= $unsigned(reg1047[(1'h0):(1'h0)]);
          for (forvar1201 = (1'h0); (forvar1201 < (3'h6)); forvar1201 = (forvar1201 + (1'h1)))
            begin
              reg1202 = {(~^reg1196)};
              reg1203 = (7'h49);
              reg1204 <= (reg1146[(4'h9):(2'h2)] ?
                  reg780 : ($unsigned($signed($signed(reg824))) || ({(reg506 ?
                          reg886 : reg857)} <<< reg1138)));
              reg1205 = $signed({$unsigned((~(reg552 ? (8'ha0) : wire429))),
                  reg528[(1'h1):(1'h0)],
                  reg457[(4'hb):(4'h8)]});
            end
          for (forvar1206 = (1'h0); (forvar1206 < (2'h3)); forvar1206 = (forvar1206 + (1'h1)))
            begin
              reg1207 <= {(7'h47)};
              reg1208 = reg1138[(3'h5):(3'h4)];
            end
          if ($signed({$unsigned(reg1148[(4'hc):(2'h2)]),
              {($signed(reg766) <= (!reg529)),
                  $unsigned(((8'hae) | reg706)),
                  $signed((reg1047 ^ reg514))},
              (7'h44)}))
            begin
              reg1209 = (reg1008[(1'h1):(1'h1)] ?
                  reg1205[(4'he):(2'h2)] : reg760);
              reg1210 <= (($signed(((^reg1151) ?
                      (|reg942) : (reg684 || reg1095))) ^~ ($unsigned(((7'h41) | reg755)) ?
                      {{reg443, reg990}} : $unsigned((reg586 ?
                          reg603 : reg1096)))) ?
                  $signed($unsigned(reg1100[(1'h0):(1'h0)])) : $unsigned(reg1106));
              reg1211 <= {($signed(((reg849 ?
                          reg1202 : (7'h4e)) << reg921[(4'ha):(3'h7)])) ?
                      {$unsigned(((7'h50) ?
                              reg1083 : reg639))} : (&reg542[(1'h0):(1'h0)]))};
              reg1212 = $unsigned(((!reg742) ?
                  reg552 : ($signed(((8'ha7) ~^ reg552)) >> reg497[(1'h0):(1'h0)])));
              reg1213 <= ({(8'ha1)} ?
                  {$unsigned({(reg695 ?
                              (7'h4e) : reg485)})} : ({(wire428[(2'h2):(1'h1)] >> $signed((7'h53))),
                          reg490[(2'h2):(1'h0)],
                          $unsigned($signed(reg1012))} ?
                      (reg964 & $signed((+reg820))) : (!($signed(reg820) ?
                          (reg450 <= wire428) : $signed((8'ha9))))));
              reg1214 <= ((^reg530) <<< $unsigned($signed(reg1120[(3'h6):(2'h3)])));
            end
          else
            begin
              reg1210 <= $unsigned(reg450);
              reg1211 <= (reg586[(4'ha):(2'h2)] >>> (~&(|reg1179)));
            end
        end
    end
  assign wire1215 = $unsigned({$unsigned(((reg503 - (8'ha7)) ?
                            (reg1076 ~^ reg525) : $signed(reg748))),
                        $unsigned(reg734[(5'h1d):(5'h13)])});
  always
    @(posedge clk) begin
      for (forvar1216 = (1'h0); (forvar1216 < (2'h3)); forvar1216 = (forvar1216 + (1'h1)))
        begin
          for (forvar1217 = (1'h0); (forvar1217 < (2'h3)); forvar1217 = (forvar1217 + (1'h1)))
            begin
              reg1218 <= reg893[(4'h8):(3'h6)];
              reg1219 = ($signed($unsigned($unsigned($signed(reg520)))) ?
                  $unsigned($unsigned($unsigned(((8'hbe) > reg530)))) : $signed(reg625));
              reg1220 = reg514;
              reg1221 <= $signed(reg482[(1'h0):(1'h0)]);
              reg1222 <= $signed((|reg866[(4'h9):(4'h9)]));
              reg1223 = ((!reg979) - (^reg603[(1'h0):(1'h0)]));
              reg1224 <= $signed(($signed(((reg511 <<< reg639) > $signed(reg1032))) && $unsigned((^~reg503[(2'h2):(1'h1)]))));
            end
          if (($unsigned(reg866) >>> reg709[(5'h17):(4'hb)]))
            begin
              reg1225 <= (~&$unsigned((($unsigned((8'hb4)) ?
                  $unsigned(reg796) : reg1137[(5'h11):(4'hc)]) - reg698[(5'h10):(3'h7)])));
              reg1226 = $signed(wire594[(4'hc):(4'hb)]);
              reg1227 = (-{$signed($unsigned(reg1087[(3'h5):(2'h2)])),
                  reg611[(3'h5):(1'h1)]});
            end
          else
            begin
              reg1226 = $unsigned($unsigned(reg599));
              reg1228 <= ($signed((wire564[(4'h8):(2'h3)] ?
                  reg650[(4'hd):(4'hb)] : $unsigned((~&(8'hb1))))) >> {(-reg747),
                  (($signed(reg1147) ?
                      reg782 : {wire1089}) - (^$unsigned(reg1117))),
                  {reg728[(4'hc):(3'h4)],
                      (^((7'h43) ^ reg1072)),
                      {((7'h4f) ? (7'h42) : reg1096), $unsigned((8'haa))}}});
            end
          if (reg882[(4'h8):(4'h8)])
            begin
              reg1229 <= {$signed($signed(((!reg551) & reg1036)))};
              reg1230 <= reg552;
              reg1231 <= {(~({{reg447},
                      {wire1089, reg1074, (8'ha3)},
                      (reg911 <<< reg650)} <= $signed($unsigned(reg654)))),
                  ($unsigned((-reg1084)) ?
                      reg575[(2'h3):(2'h3)] : (reg707[(2'h3):(1'h1)] != reg992[(1'h1):(1'h1)]))};
              reg1232 = ((($signed(wire426[(5'h19):(1'h0)]) >>> $signed(reg672)) != (7'h55)) > $unsigned(reg654));
              reg1233 = $unsigned($signed($unsigned((~&wire678[(2'h3):(1'h0)]))));
              reg1234 = (reg1063 * (reg921[(3'h5):(1'h1)] + ($signed((8'ha2)) ?
                  (~&(reg528 < reg1171)) : (reg1056 | (reg463 * reg712)))));
            end
          else
            begin
              reg1229 <= $signed(forvar1216[(5'h11):(2'h2)]);
              reg1232 = ((reg912 ?
                      (($signed(reg1181) ?
                              reg972[(4'hd):(4'h9)] : $unsigned(reg469)) ?
                          ($unsigned(reg546) ?
                              (&(7'h46)) : {reg603,
                                  (8'hb8)}) : reg1175) : reg1207[(3'h5):(2'h3)]) ?
                  $unsigned($unsigned(reg1005)) : wire678[(3'h7):(3'h6)]);
              reg1235 <= reg457[(4'hd):(1'h1)];
              reg1236 = ((~&(reg620 ?
                      $signed((~^reg1041)) : {$unsigned(reg640),
                          (reg814 <= (8'hb5)),
                          {reg755, reg452, reg872}})) ?
                  ((&(-{reg755, reg882})) ^ ($unsigned((reg454 ?
                      (7'h54) : reg510)) + ((8'h9f) || (reg813 ?
                      reg1134 : reg871)))) : (($signed({reg469}) >= $signed(reg1214[(5'h13):(2'h3)])) && ((((7'h56) ?
                          reg930 : reg816) ?
                      {reg1025,
                          reg1229,
                          reg1234} : $unsigned(reg452)) ^ (7'h43))));
            end
          reg1237 = ({reg573[(2'h3):(1'h0)],
                  reg743[(4'hd):(3'h5)],
                  $signed((~^(reg1069 ? reg1142 : reg676)))} ?
              reg1077[(5'h1a):(4'hb)] : reg806[(3'h7):(3'h7)]);
        end
      reg1238 <= reg511;
      reg1239 <= reg717[(4'hc):(3'h7)];
      for (forvar1240 = (1'h0); (forvar1240 < (3'h6)); forvar1240 = (forvar1240 + (1'h1)))
        begin
          if ((({((reg1056 ? reg433 : (8'h9f)) ^~ ((7'h57) ? reg586 : reg979)),
                      (~^$signed((8'h9e)))} ?
                  reg443 : $signed(((reg1095 <<< reg883) <<< {reg813}))) ?
              ($signed(reg766) ?
                  $unsigned(($unsigned(reg605) ^ $signed(reg777))) : reg1001[(1'h1):(1'h0)]) : {(reg1054 != $unsigned(reg1072[(4'hc):(3'h5)])),
                  ($unsigned(reg963) || $signed(reg746)),
                  $signed({(reg650 ? reg957 : reg732),
                      (reg655 - reg1039),
                      $unsigned(reg1167)})}))
            begin
              reg1241 = reg520[(1'h0):(1'h0)];
              reg1242 = $signed($signed(({reg1186} ^~ ((reg1008 ?
                  reg1085 : reg911) <<< $signed(reg957)))));
            end
          else
            begin
              reg1243 <= $signed(reg1049[(4'hb):(4'h9)]);
              reg1244 = {$signed(reg700[(2'h3):(1'h0)])};
              reg1245 = (reg433 >= (reg1056[(4'hb):(4'hb)] >>> $unsigned(((reg804 && reg552) << reg1186[(1'h1):(1'h0)]))));
              reg1246 <= {$signed((($unsigned(reg438) > (reg935 + reg1037)) | $unsigned(reg586[(5'h10):(5'h10)])))};
              reg1247 <= (~|(7'h4e));
              reg1248 = $signed(reg1025[(2'h3):(2'h3)]);
            end
          if (((+(~{(reg814 == reg1227)})) < reg450[(2'h2):(1'h0)]))
            begin
              reg1249 = reg740;
              reg1250 = $signed($signed((-reg562)));
            end
          else
            begin
              reg1251 <= reg1146[(4'ha):(3'h5)];
              reg1252 <= $signed((-((8'ha5) && (reg723[(3'h4):(2'h3)] ?
                  (reg460 ? (7'h55) : reg780) : $unsigned(reg437)))));
              reg1253 <= {reg558[(2'h3):(1'h0)]};
              reg1254 <= ($signed({reg1248,
                  $signed($unsigned(reg920)),
                  ({reg1119} | (~(7'h48)))}) == reg972[(3'h4):(2'h3)]);
              reg1255 <= ($signed($unsigned(((reg562 <= reg604) ?
                      reg572 : {reg700}))) ?
                  reg871[(3'h5):(2'h3)] : reg466);
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg1194)
        begin
          reg1256 = wire425;
          reg1257 = reg1027[(3'h6):(3'h5)];
          if ($unsigned((reg1019 ?
              reg734 : {reg796,
                  $signed((reg1181 <= reg897)),
                  $unsigned((reg915 ? reg995 : wire430))})))
            begin
              reg1258 = $signed(($unsigned(reg1225[(3'h5):(2'h3)]) ?
                  $signed($signed($unsigned((8'hb1)))) : $signed(reg771)));
              reg1259 = reg1178[(4'he):(4'hc)];
            end
          else
            begin
              reg1258 = reg495;
              reg1260 <= {reg1097[(1'h1):(1'h0)],
                  (reg983[(5'h10):(4'h9)] == reg949[(4'he):(4'h8)])};
              reg1261 <= $unsigned((reg467 < reg814));
              reg1262 = {(~^(!(!reg542))),
                  ((^~reg1172) >= reg1260[(1'h0):(1'h0)]),
                  (({$signed((8'hb4))} & (^(reg455 ?
                      reg1062 : (7'h55)))) > $unsigned((+$unsigned(reg928))))};
              reg1263 = {reg438};
              reg1264 = $signed((-$unsigned((!$signed(reg960)))));
            end
        end
      else
        begin
          reg1260 <= ((((^$unsigned((8'hb6))) ?
                  (~{reg944, (8'hbb), reg485}) : {(7'h54),
                      $signed(reg529),
                      reg1005}) ?
              reg1065[(4'hb):(3'h6)] : ({$unsigned(reg490)} ?
                  reg1204[(4'he):(4'ha)] : $signed((^~reg1150)))) >>> reg525[(3'h7):(2'h2)]);
          reg1262 = $unsigned($signed(reg990));
        end
    end
  assign wire1265 = $signed($unsigned(reg1224));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module179
#(parameter param312 = {(~|((((7'h44) >= (8'haa)) >= (!(7'h43))) < (((8'ha6) ^ (8'hb4)) <<< ((8'hbf) + (8'h9e))))), (~|((|((7'h53) ? (8'hb1) : (8'ha2))) + {{(8'ha1), (7'h44)}, ((8'hb0) & (7'h58))}))})
(y, clk, wire185, wire184, wire183, wire182, wire181, wire180);
  output wire [(32'h79f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire185;
  input wire signed [(3'h6):(1'h0)] wire184;
  input wire signed [(5'h1a):(1'h0)] wire183;
  input wire signed [(4'hb):(1'h0)] wire182;
  input wire [(5'h19):(1'h0)] wire181;
  input wire [(4'hd):(1'h0)] wire180;
  wire signed [(5'h1e):(1'h0)] wire311;
  wire [(3'h4):(1'h0)] wire310;
  wire [(4'hc):(1'h0)] wire237;
  wire [(3'h4):(1'h0)] wire236;
  wire signed [(5'h17):(1'h0)] wire188;
  reg signed [(4'h9):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg307 = (1'h0);
  reg [(5'h18):(1'h0)] reg305 = (1'h0);
  reg [(5'h10):(1'h0)] reg304 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg303 = (1'h0);
  reg [(5'h1c):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg298 = (1'h0);
  reg [(4'hd):(1'h0)] reg297 = (1'h0);
  reg [(3'h4):(1'h0)] reg296 = (1'h0);
  reg [(3'h5):(1'h0)] reg295 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg293 = (1'h0);
  reg [(3'h7):(1'h0)] reg290 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg289 = (1'h0);
  reg [(4'h8):(1'h0)] reg287 = (1'h0);
  reg [(5'h1d):(1'h0)] reg285 = (1'h0);
  reg [(4'ha):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg281 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg277 = (1'h0);
  reg [(4'he):(1'h0)] reg276 = (1'h0);
  reg [(5'h11):(1'h0)] reg275 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg270 = (1'h0);
  reg [(5'h18):(1'h0)] reg269 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg265 = (1'h0);
  reg [(4'hc):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg258 = (1'h0);
  reg [(5'h14):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg254 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg249 = (1'h0);
  reg [(4'hc):(1'h0)] reg245 = (1'h0);
  reg [(5'h14):(1'h0)] reg235 = (1'h0);
  reg [(5'h1e):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg233 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg230 = (1'h0);
  reg [(5'h1a):(1'h0)] reg229 = (1'h0);
  reg [(4'h8):(1'h0)] reg227 = (1'h0);
  reg [(4'hc):(1'h0)] reg226 = (1'h0);
  reg [(3'h5):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg220 = (1'h0);
  reg [(3'h7):(1'h0)] reg218 = (1'h0);
  reg [(5'h1b):(1'h0)] reg217 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg216 = (1'h0);
  reg [(4'ha):(1'h0)] reg215 = (1'h0);
  reg [(3'h6):(1'h0)] reg214 = (1'h0);
  reg [(4'hf):(1'h0)] reg213 = (1'h0);
  reg [(5'h15):(1'h0)] reg212 = (1'h0);
  reg [(3'h6):(1'h0)] reg209 = (1'h0);
  reg [(5'h1e):(1'h0)] reg204 = (1'h0);
  reg [(5'h14):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg196 = (1'h0);
  reg [(2'h2):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg187 = (1'h0);
  reg [(2'h3):(1'h0)] reg186 = (1'h0);
  reg [(4'ha):(1'h0)] reg308 = (1'h0);
  reg [(3'h6):(1'h0)] reg306 = (1'h0);
  reg [(4'hc):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg301 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar299 = (1'h0);
  reg [(3'h4):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg292 = (1'h0);
  reg [(5'h19):(1'h0)] reg291 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg288 = (1'h0);
  reg [(3'h4):(1'h0)] reg286 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar284 = (1'h0);
  reg [(5'h1c):(1'h0)] reg283 = (1'h0);
  reg [(3'h5):(1'h0)] reg280 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar279 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg272 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg271 = (1'h0);
  reg [(4'hc):(1'h0)] reg267 = (1'h0);
  reg [(5'h10):(1'h0)] reg263 = (1'h0);
  reg [(3'h5):(1'h0)] forvar262 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg261 = (1'h0);
  reg [(4'hc):(1'h0)] reg260 = (1'h0);
  reg [(5'h10):(1'h0)] reg259 = (1'h0);
  reg [(5'h10):(1'h0)] reg257 = (1'h0);
  reg [(4'hd):(1'h0)] reg255 = (1'h0);
  reg [(5'h16):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg251 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg250 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg248 = (1'h0);
  reg [(5'h12):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg246 = (1'h0);
  reg [(5'h11):(1'h0)] forvar244 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar243 = (1'h0);
  reg [(3'h7):(1'h0)] reg242 = (1'h0);
  reg [(4'hb):(1'h0)] reg241 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg240 = (1'h0);
  reg [(5'h13):(1'h0)] forvar239 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar238 = (1'h0);
  reg [(4'hc):(1'h0)] reg232 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar228 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg225 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar224 = (1'h0);
  reg [(4'hb):(1'h0)] reg223 = (1'h0);
  reg signed [(4'he):(1'h0)] reg221 = (1'h0);
  reg [(5'h15):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg211 = (1'h0);
  reg [(2'h3):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg199 = (1'h0);
  reg [(5'h1f):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg207 = (1'h0);
  reg [(2'h2):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg205 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg201 = (1'h0);
  reg [(4'ha):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar199 = (1'h0);
  reg [(3'h7):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg197 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg195 = (1'h0);
  reg [(4'hc):(1'h0)] forvar194 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar193 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg192 = (1'h0);
  reg [(5'h10):(1'h0)] reg191 = (1'h0);
  reg [(5'h15):(1'h0)] reg190 = (1'h0);
  assign y = {wire311,
                 wire310,
                 wire237,
                 wire236,
                 wire188,
                 reg309,
                 reg307,
                 reg305,
                 reg304,
                 reg303,
                 reg300,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg293,
                 reg290,
                 reg289,
                 reg287,
                 reg285,
                 reg282,
                 reg281,
                 reg277,
                 reg276,
                 reg275,
                 reg273,
                 reg270,
                 reg269,
                 reg268,
                 reg266,
                 reg265,
                 reg264,
                 reg258,
                 reg256,
                 reg254,
                 reg253,
                 reg249,
                 reg245,
                 reg235,
                 reg234,
                 reg233,
                 reg230,
                 reg229,
                 reg227,
                 reg226,
                 reg222,
                 reg220,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg209,
                 reg204,
                 reg203,
                 reg202,
                 reg196,
                 reg189,
                 reg187,
                 reg186,
                 reg308,
                 reg306,
                 reg302,
                 reg301,
                 forvar299,
                 reg294,
                 reg292,
                 reg291,
                 reg288,
                 reg286,
                 forvar284,
                 reg283,
                 reg280,
                 forvar279,
                 reg278,
                 reg274,
                 reg272,
                 reg271,
                 reg267,
                 reg263,
                 forvar262,
                 reg261,
                 reg260,
                 reg259,
                 reg257,
                 reg255,
                 reg252,
                 reg251,
                 reg250,
                 reg248,
                 reg247,
                 reg246,
                 forvar244,
                 forvar243,
                 reg242,
                 reg241,
                 reg240,
                 forvar239,
                 forvar238,
                 reg232,
                 reg231,
                 forvar228,
                 reg225,
                 forvar224,
                 reg223,
                 reg221,
                 reg219,
                 reg211,
                 reg210,
                 reg199,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg201,
                 reg200,
                 forvar199,
                 reg198,
                 reg197,
                 reg195,
                 forvar194,
                 forvar193,
                 reg192,
                 reg191,
                 reg190,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg186 <= ($unsigned($signed(wire181[(3'h4):(3'h4)])) && $signed($unsigned($signed((wire183 ?
          wire183 : wire183)))));
      reg187 <= (-(!{(((8'h9e) << (7'h43)) ?
              $unsigned((8'ha3)) : $unsigned(wire181)),
          (reg186[(1'h1):(1'h0)] ~^ (^wire182))}));
    end
  assign wire188 = $unsigned(reg186);
  always
    @(posedge clk) begin
      reg189 <= (wire184 ^ ((~|reg186[(2'h3):(1'h0)]) <<< wire182[(4'h8):(3'h6)]));
      reg190 = reg186[(1'h1):(1'h0)];
      reg191 = ($signed($signed((!(wire188 ?
          (8'h9c) : wire188)))) >>> ($signed(reg187) ?
          ($unsigned($signed(wire188)) <= (~^(^~(7'h48)))) : ((wire182[(3'h7):(3'h7)] | (wire188 >>> wire182)) - $signed((+(8'ha8))))));
      reg192 = (~((~(~^(!wire183))) < ((^$unsigned(reg189)) ?
          ((wire180 == reg190) << (wire184 < (8'hb3))) : {wire185,
              wire183[(4'hc):(4'hb)]})));
      for (forvar193 = (1'h0); (forvar193 < (1'h1)); forvar193 = (forvar193 + (1'h1)))
        begin
          for (forvar194 = (1'h0); (forvar194 < (1'h1)); forvar194 = (forvar194 + (1'h1)))
            begin
              reg195 = wire184[(1'h0):(1'h0)];
              reg196 <= wire188;
              reg197 = ($unsigned(($unsigned({reg190, reg196}) ?
                      reg190[(5'h13):(3'h7)] : (~|wire180[(3'h6):(1'h1)]))) ?
                  {((reg190[(3'h4):(1'h1)] >> (reg189 ~^ wire184)) ?
                          forvar194 : ({(8'ha5),
                              wire180,
                              forvar194} == reg187[(5'h10):(1'h1)]))} : $unsigned($unsigned($unsigned($signed((8'hb5))))));
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed((&{wire184[(3'h6):(2'h2)]})))
        begin
          reg198 = ((((~&$unsigned(wire185)) && {$unsigned(wire181)}) ?
                  reg187 : wire181[(2'h2):(1'h0)]) ?
              reg187 : (~^$unsigned(({reg189, reg189, reg186} ?
                  (8'ha9) : (~^wire185)))));
          for (forvar199 = (1'h0); (forvar199 < (3'h5)); forvar199 = (forvar199 + (1'h1)))
            begin
              reg200 = $signed(($unsigned((wire182 <= wire180[(4'h8):(3'h4)])) ?
                  $unsigned(($signed(wire185) >> reg198[(2'h3):(2'h3)])) : wire184));
              reg201 = forvar199;
            end
          if ((7'h50))
            begin
              reg202 <= (reg189 << ($unsigned(wire185) ?
                  (((8'hbb) <<< (!(8'hac))) ?
                      ({reg187, (7'h4e), reg189} ?
                          (|reg201) : (reg201 ? reg196 : wire180)) : ({wire183,
                              wire181} ?
                          $signed(wire185) : (wire181 | reg189))) : {($signed(wire182) | (!reg187)),
                      ($unsigned(reg196) * $unsigned(reg198)),
                      (-$unsigned(wire183))}));
              reg203 <= ($signed($signed($signed(((7'h43) ?
                  reg189 : (7'h54))))) != (reg187[(5'h1f):(5'h18)] || {(wire188[(4'hb):(3'h7)] ?
                      wire184[(2'h3):(2'h2)] : (-wire185)),
                  (|(reg202 ? wire185 : wire184))}));
              reg204 <= $unsigned(wire183[(4'hb):(1'h0)]);
              reg205 = (((^$unsigned($unsigned(wire183))) ~^ wire180) ?
                  ($unsigned(wire180) & $unsigned(($signed(wire185) ?
                      $signed(reg203) : {reg204,
                          forvar199,
                          reg186}))) : $signed($signed(({reg198} <<< wire180[(4'hd):(1'h1)]))));
            end
          else
            begin
              reg205 = forvar199;
              reg206 = {$unsigned(reg200),
                  (~&$unsigned($signed($signed(wire184))))};
            end
          reg207 = wire180;
          reg208 = $unsigned(((^~(^(8'hb6))) >= $signed(($unsigned(wire183) && wire188[(5'h11):(4'h8)]))));
          reg209 <= (-reg208[(3'h6):(1'h1)]);
        end
      else
        begin
          reg198 = (((8'ha5) ?
              {$signed((wire184 ? (7'h4b) : wire185))} : {reg202[(4'ha):(1'h1)],
                  $unsigned($signed(reg186))}) ^~ reg187[(2'h2):(1'h0)]);
          if ($unsigned(reg208[(5'h1e):(4'h8)]))
            begin
              reg199 = $unsigned(({reg203[(3'h4):(2'h2)],
                  ((wire188 + reg206) ?
                      (reg209 ? reg201 : (8'ha1)) : $signed(reg204)),
                  wire180[(3'h7):(3'h7)]} ^~ ((8'hb7) ?
                  ($unsigned(reg204) ?
                      wire180[(2'h2):(1'h0)] : $signed((8'ha3))) : $signed((reg206 ?
                      (8'ha4) : reg205)))));
              reg200 = wire184[(3'h5):(2'h3)];
              reg201 = {reg204,
                  (^(^$signed((reg199 | reg206)))),
                  ($signed(reg208) ?
                      (8'h9c) : (($signed(reg187) ?
                          (reg201 | (8'h9f)) : (^~(7'h4d))) ^ $unsigned((reg207 & (8'hb0)))))};
            end
          else
            begin
              reg199 = ((|(($signed((8'hb1)) ?
                  reg202 : $signed((8'hbd))) <= wire184)) || (^~reg208[(5'h10):(4'he)]));
              reg202 <= ($signed((+({wire188, (7'h44), reg203} ?
                      {(7'h4b), wire180, (8'ha4)} : (+reg202)))) ?
                  $unsigned($unsigned(wire188)) : (+{((8'ha3) ?
                          reg196 : reg187),
                      $signed(forvar199[(2'h3):(1'h1)])}));
              reg205 = ((-reg209[(3'h6):(2'h3)]) ?
                  wire185[(3'h5):(2'h3)] : {$unsigned(((wire188 * wire180) ?
                          {reg199, reg204} : reg187[(5'h18):(4'hc)]))});
              reg206 = reg204;
            end
          if (wire180)
            begin
              reg207 = (((reg209 ?
                      ({reg199, reg208} - reg204) : (((7'h54) << reg201) ?
                          {(8'ha2)} : $unsigned(reg202))) | reg207) ?
                  wire188 : (8'hb2));
              reg208 = reg203;
            end
          else
            begin
              reg209 <= ((|$signed(((+reg205) ?
                      $signed((7'h50)) : (reg202 - reg198)))) ?
                  $unsigned((reg205[(1'h1):(1'h0)] ^~ wire184)) : $signed($unsigned(((wire180 != (7'h46)) * (~^reg200)))));
              reg210 = reg199;
              reg211 = ((~|wire185[(3'h4):(3'h4)]) ?
                  $unsigned(reg209) : reg204);
            end
          if (((wire185[(3'h7):(1'h0)] >> {reg210}) ?
              ($signed($signed(wire185)) ?
                  reg205 : {((8'ha0) + reg206)}) : {($signed(((8'hae) ?
                      wire182 : reg186)) >= ((^(7'h4c)) ?
                      $unsigned(reg196) : $signed(reg209)))}))
            begin
              reg212 <= $signed($unsigned(wire180[(4'hd):(3'h6)]));
              reg213 <= (!$signed(wire182));
            end
          else
            begin
              reg212 <= $signed(reg208[(4'h9):(3'h5)]);
              reg213 <= wire188;
              reg214 <= {(wire181[(3'h5):(1'h0)] > ((reg198[(3'h7):(3'h5)] ?
                          {reg209} : (reg186 == reg196)) ?
                      $signed(((8'hb3) == reg186)) : $unsigned((^~(8'hbe)))))};
              reg215 <= reg203[(5'h12):(2'h2)];
              reg216 <= reg186;
              reg217 <= (reg189[(1'h0):(1'h0)] || {$unsigned({(reg209 ?
                          wire184 : (8'ha5))})});
            end
          if (reg198[(1'h0):(1'h0)])
            begin
              reg218 <= {$signed((reg186[(1'h1):(1'h0)] ?
                      $signed($unsigned(reg212)) : ($signed(reg200) < $unsigned((7'h57))))),
                  wire181[(5'h15):(5'h15)]};
              reg219 = ((~^$signed(reg203[(4'hb):(3'h4)])) ~^ (($unsigned((~reg209)) ?
                  $signed((reg204 | reg215)) : $signed($unsigned((8'ha5)))) + ($signed(reg203[(1'h1):(1'h0)]) != (^{reg203}))));
              reg220 <= $unsigned((&$unsigned((^{reg209}))));
              reg221 = $signed({(+$unsigned({reg204, reg203}))});
            end
          else
            begin
              reg218 <= ($unsigned(((reg212[(4'he):(4'h9)] ?
                          {reg204} : $signed((8'hb9))) ?
                      (!(reg212 ? reg186 : reg219)) : (|$unsigned(wire182)))) ?
                  ($signed((reg186[(2'h2):(1'h0)] * (forvar199 ?
                          wire180 : reg210))) ?
                      reg216 : (^((reg208 ?
                          reg218 : reg202) || reg204))) : ((~|wire182) <<< {{(^~(8'hb3))}}));
              reg219 = ($unsigned($unsigned(((reg196 ?
                      reg213 : reg205) * (~|wire182)))) ?
                  reg211[(4'hf):(3'h5)] : (($signed(wire182) + $unsigned(wire183)) > (~|$unsigned($signed(reg201)))));
              reg220 <= $unsigned($signed(((reg189 ?
                      $signed(reg215) : reg209[(1'h0):(1'h0)]) ?
                  reg213[(4'hc):(1'h1)] : (((8'hb0) ?
                      reg198 : (8'hb8)) + (reg205 ? (8'ha1) : wire185)))));
              reg222 <= $unsigned($unsigned(reg217[(3'h4):(3'h4)]));
              reg223 = (&((reg208 >= reg199[(4'he):(4'he)]) ?
                  reg200[(1'h1):(1'h0)] : wire180[(4'hb):(3'h7)]));
            end
        end
      for (forvar224 = (1'h0); (forvar224 < (3'h5)); forvar224 = (forvar224 + (1'h1)))
        begin
          if ((wire181 >= ($signed((reg202 ?
                  $unsigned(reg219) : (reg216 != reg213))) ?
              wire184 : (|({reg203} < (8'hb9))))))
            begin
              reg225 = $unsigned(reg222[(1'h0):(1'h0)]);
              reg226 <= {(8'ha3),
                  $signed(reg222[(3'h4):(1'h1)]),
                  $signed($unsigned(forvar224[(4'hc):(1'h1)]))};
              reg227 <= ((reg203 ?
                  {$signed($unsigned(wire188))} : reg186[(2'h2):(1'h0)]) * wire181[(5'h16):(5'h15)]);
            end
          else
            begin
              reg225 = ((|(($signed(wire183) ^ reg200) * $unsigned(wire181))) ?
                  wire185 : {$unsigned($unsigned(reg210))});
            end
          for (forvar228 = (1'h0); (forvar228 < (3'h6)); forvar228 = (forvar228 + (1'h1)))
            begin
              reg229 <= $signed({$unsigned(reg207[(4'hb):(3'h7)]),
                  wire182,
                  ({(reg227 == reg214)} ?
                      (~^$unsigned(wire184)) : {(reg211 ? reg198 : reg220),
                          reg205,
                          (reg198 ? reg216 : (7'h56))})});
              reg230 <= reg200[(4'h9):(2'h3)];
              reg231 = $unsigned($signed((!(~&(wire183 ? wire183 : (8'ha6))))));
              reg232 = wire185[(2'h2):(1'h1)];
            end
          reg233 <= (wire181[(4'h9):(3'h6)] <<< ($signed($signed(forvar224)) ^ $signed((reg204 ?
              reg213 : {(8'hac), wire188, reg229}))));
          reg234 <= {(reg226[(3'h5):(1'h1)] <= (($signed(forvar224) >= (~^reg196)) >> $signed($unsigned(reg227)))),
              (reg187 ?
                  reg204[(4'hf):(2'h2)] : ($unsigned($signed(wire184)) ?
                      {(reg207 ? (8'hbb) : reg225)} : ((reg205 <<< (7'h47)) ?
                          (wire182 ?
                              reg205 : reg232) : reg217[(3'h6):(3'h4)]))),
              (~&wire184[(2'h2):(2'h2)])};
          reg235 <= reg212[(3'h7):(2'h3)];
        end
    end
  assign wire236 = $unsigned($unsigned($signed(reg213[(2'h2):(1'h0)])));
  assign wire237 = (^~$signed(((wire185[(3'h5):(2'h2)] >>> $unsigned(reg235)) == $signed((reg215 || wire188)))));
  always
    @(posedge clk) begin
      for (forvar238 = (1'h0); (forvar238 < (3'h4)); forvar238 = (forvar238 + (1'h1)))
        begin
          for (forvar239 = (1'h0); (forvar239 < (3'h5)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg240 = ((7'h57) >>> (reg227 | (wire181[(2'h2):(1'h1)] | (!wire181))));
              reg241 = ($unsigned((~^(((7'h45) ? reg215 : (8'h9e)) ?
                  wire180 : reg216))) > reg203[(4'h9):(4'h8)]);
              reg242 = reg234;
            end
        end
      for (forvar243 = (1'h0); (forvar243 < (1'h0)); forvar243 = (forvar243 + (1'h1)))
        begin
          for (forvar244 = (1'h0); (forvar244 < (1'h1)); forvar244 = (forvar244 + (1'h1)))
            begin
              reg245 <= {(reg235[(4'he):(4'hc)] >> $signed((~|(forvar239 <<< wire183)))),
                  $unsigned({reg187}),
                  $signed(forvar239)};
              reg246 = (!reg242);
              reg247 = $signed($unsigned({((7'h46) == {wire237, reg233})}));
              reg248 = (({$unsigned($signed(reg246)),
                          $signed((reg212 - reg230))} ?
                      $signed((~^(!reg227))) : ((reg204 ^ (reg242 ?
                              reg187 : wire188)) ?
                          {$signed(reg202),
                              wire183[(5'h14):(5'h14)],
                              reg247} : ((+reg230) ?
                              reg212 : (wire236 || reg189)))) ?
                  $signed(reg186) : ({{{reg186, reg209, forvar239}},
                      $unsigned($signed(reg235)),
                      (^((8'ha2) ?
                          wire188 : reg214))} >> $signed((&$unsigned(wire188)))));
              reg249 <= ($signed((&(-$unsigned(wire236)))) ?
                  reg196 : reg215[(1'h0):(1'h0)]);
              reg250 = (reg245[(4'ha):(2'h3)] && reg235[(4'hf):(3'h7)]);
            end
          reg251 = $signed($unsigned((reg196 <= $unsigned(((7'h44) || reg220)))));
          if ($unsigned($unsigned(($unsigned($signed(reg247)) < reg246))))
            begin
              reg252 = ((reg189 ~^ ((reg251 == {reg230,
                      forvar238}) ~^ $unsigned($unsigned(reg202)))) ?
                  (reg213[(4'he):(3'h5)] ?
                      ($signed((reg216 ? reg218 : reg233)) ?
                          (^(reg215 ? reg246 : reg229)) : (~^{reg196,
                              reg218})) : $unsigned(((wire236 ?
                              (7'h51) : forvar243) ?
                          (reg241 ?
                              (8'ha2) : reg249) : (7'h45)))) : (($unsigned(reg217[(5'h1b):(4'hc)]) * (reg229[(4'h9):(1'h1)] | $signed(reg251))) ?
                      reg218[(3'h7):(3'h4)] : ({(reg218 <= reg251),
                          $signed(forvar244)} >> ((wire236 | wire236) << reg212[(1'h1):(1'h0)]))));
              reg253 <= reg226;
              reg254 <= (!$signed($signed($unsigned((7'h40)))));
            end
          else
            begin
              reg252 = reg202[(5'h15):(4'hf)];
              reg253 <= (reg218[(3'h7):(3'h6)] ~^ reg235[(4'hf):(1'h1)]);
              reg255 = $unsigned({reg254});
              reg256 <= ($signed(wire183[(1'h1):(1'h1)]) ~^ $signed((&$signed((&(8'h9d))))));
              reg257 = {{{$unsigned(reg217)},
                      (^~$unsigned(reg230[(4'h8):(1'h1)]))},
                  ($unsigned(reg187) ?
                      $signed({$unsigned(reg222),
                          reg218[(3'h5):(2'h3)]}) : $signed((7'h40)))};
            end
          if ((!$unsigned(wire180)))
            begin
              reg258 <= $signed(({{(~^wire237), {reg257}},
                      ((7'h49) ^~ (reg249 * wire237)),
                      (|(~|reg254))} ?
                  reg222[(2'h2):(1'h1)] : reg257));
              reg259 = ($unsigned((^$unsigned(((8'ha1) > reg254)))) ?
                  reg187 : reg227);
              reg260 = $signed(($signed($signed((-reg249))) ?
                  reg256 : ($signed((reg234 ?
                      (7'h4c) : reg196)) < (&$unsigned(reg241)))));
              reg261 = {reg226};
            end
          else
            begin
              reg259 = (&reg203[(4'hb):(3'h6)]);
              reg260 = (~^$signed(reg256[(2'h3):(1'h0)]));
              reg261 = (~&$unsigned(((+(-reg247)) == $signed(((8'hb6) ?
                  reg186 : reg261)))));
            end
          for (forvar262 = (1'h0); (forvar262 < (1'h0)); forvar262 = (forvar262 + (1'h1)))
            begin
              reg263 = ({$signed($signed($unsigned(reg214))),
                  $signed((!wire182))} != (~&$unsigned($signed($signed(wire181)))));
              reg264 <= ({({reg245, (reg256 ? wire182 : reg212)} ?
                          reg257 : (&wire183)),
                      ($signed($signed(reg226)) + {$unsigned(reg229),
                          $unsigned((8'ha7)),
                          reg189})} ?
                  (8'h9f) : $signed((wire184[(3'h4):(1'h1)] > $unsigned({(8'h9e),
                      reg241}))));
              reg265 <= reg217;
              reg266 <= $unsigned(({($unsigned(reg253) ?
                      (reg263 ?
                          reg229 : (8'hab)) : $unsigned(reg213))} && (reg261[(5'h15):(3'h4)] ~^ $signed($signed(reg234)))));
              reg267 = ((8'hb8) ?
                  {$signed(($unsigned(wire183) ?
                          reg264[(3'h5):(2'h2)] : $unsigned(reg229))),
                      $unsigned($unsigned($signed((8'hb6))))} : $unsigned((wire236 ?
                      $signed((^~reg218)) : reg256[(4'hf):(4'hc)])));
              reg268 <= (|((8'hbd) ?
                  ({reg254[(4'ha):(1'h1)], (reg259 ? reg227 : reg261)} ?
                      ((~^forvar262) ?
                          $unsigned(reg209) : ((8'ha4) || reg256)) : reg187) : ((~|$signed(reg187)) <<< $signed(((7'h55) ?
                      reg254 : (7'h51))))));
              reg269 <= (~^reg189);
            end
          if (forvar239[(1'h0):(1'h0)])
            begin
              reg270 <= (7'h54);
            end
          else
            begin
              reg271 = ($unsigned((^~(reg240 <= (!reg266)))) << $signed((((^reg258) || $signed(reg259)) * {$signed(reg212),
                  {reg220}})));
              reg272 = $unsigned($signed({reg234[(5'h12):(1'h1)]}));
              reg273 <= reg250;
              reg274 = (8'ha4);
              reg275 <= $signed(forvar262);
              reg276 <= reg220[(2'h3):(2'h2)];
              reg277 <= reg254[(3'h4):(2'h2)];
            end
        end
      reg278 = wire188[(4'h9):(1'h0)];
      for (forvar279 = (1'h0); (forvar279 < (2'h2)); forvar279 = (forvar279 + (1'h1)))
        begin
          reg280 = reg233;
          if (($signed({reg230[(2'h3):(1'h1)],
                  $signed(reg229[(4'ha):(4'h8)])}) ?
              reg217 : (7'h52)))
            begin
              reg281 <= {((|((reg245 ? reg242 : reg246) && $signed(reg235))) ?
                      (~&{(reg247 ? reg257 : reg271)}) : $signed(((^(8'hbb)) ?
                          (reg229 >= reg204) : (reg229 | wire181)))),
                  reg189};
            end
          else
            begin
              reg281 <= (^~reg251[(5'h1b):(5'h1b)]);
              reg282 <= ($signed($unsigned(reg265)) <= $signed((reg264[(4'h8):(3'h5)] ?
                  reg249 : reg226[(4'ha):(4'h9)])));
            end
          reg283 = ((7'h42) <= $unsigned($unsigned($signed((~|reg271)))));
          for (forvar284 = (1'h0); (forvar284 < (1'h1)); forvar284 = (forvar284 + (1'h1)))
            begin
              reg285 <= reg216[(3'h5):(3'h4)];
              reg286 = $unsigned(((~(!reg235)) ^~ {((forvar243 != reg271) - ((8'hbb) ?
                      reg203 : wire237))}));
              reg287 <= (8'h9e);
              reg288 = $signed((|reg196[(3'h4):(2'h2)]));
              reg289 <= $unsigned(reg222[(3'h5):(2'h3)]);
              reg290 <= $unsigned(reg282);
            end
          reg291 = $unsigned($unsigned($signed(reg234[(5'h1b):(5'h18)])));
          if ((~^{$signed(($unsigned(reg259) ~^ {forvar262, (8'hbd), reg222})),
              (reg278[(1'h0):(1'h0)] | (7'h49)),
              (((reg249 ?
                  (8'ha5) : reg196) || ((8'had) >> reg268)) <<< (8'hba))}))
            begin
              reg292 = ((wire237 ?
                      reg275[(4'he):(4'hd)] : reg273[(1'h1):(1'h0)]) ?
                  (reg220 > {(~|{reg187, reg212}),
                      reg213}) : $signed((((wire188 < reg212) - {reg218,
                      reg216}) ~^ (+$signed(wire237)))));
              reg293 <= $unsigned({(8'ha3)});
            end
          else
            begin
              reg293 <= $unsigned(forvar239[(3'h5):(3'h4)]);
              reg294 = ($unsigned(($signed($unsigned(wire183)) << reg250[(4'hd):(3'h6)])) || forvar279[(1'h1):(1'h0)]);
              reg295 <= ((7'h54) ?
                  reg270[(5'h11):(2'h2)] : ((({(8'ha9),
                      reg281} >>> reg277[(2'h2):(2'h2)]) - $signed(reg226[(1'h0):(1'h0)])) - (~forvar284)));
              reg296 <= (^~(reg226[(2'h3):(2'h3)] ?
                  reg227[(4'h8):(1'h0)] : $signed((~(~|reg276)))));
              reg297 <= reg241;
              reg298 <= {(reg222 <= (~|reg270)), reg277};
            end
        end
      for (forvar299 = (1'h0); (forvar299 < (1'h1)); forvar299 = (forvar299 + (1'h1)))
        begin
          if (($unsigned((reg253 - reg290[(3'h4):(2'h2)])) + reg217))
            begin
              reg300 <= (((+(^~{reg214, reg227})) ?
                  reg255[(2'h3):(1'h0)] : reg203) >>> reg230);
              reg301 = $signed(forvar284);
              reg302 = {(((~forvar279) != reg222[(2'h2):(1'h0)]) ?
                      {(8'h9c),
                          ((^reg278) * $signed(reg256)),
                          forvar243} : ((reg276[(1'h1):(1'h1)] ?
                              $signed(reg230) : reg267[(3'h7):(1'h1)]) ?
                          ($signed(forvar238) ~^ (reg186 ?
                              reg277 : reg270)) : {((8'ha5) ?
                                  reg283 : reg267)})),
                  reg240};
              reg303 <= (wire185[(1'h0):(1'h0)] ?
                  (&(~&$signed({reg256}))) : ((^~({reg186,
                      reg269} ~^ reg260[(1'h1):(1'h0)])) << $signed($signed((reg209 ?
                      wire236 : (8'hb3))))));
              reg304 <= $unsigned(reg204);
              reg305 <= {reg297};
            end
          else
            begin
              reg301 = $unsigned((~|$signed(({reg268} + ((7'h51) ?
                  reg266 : reg255)))));
              reg303 <= $signed((+(&(7'h45))));
              reg306 = reg274[(5'h13):(4'h9)];
              reg307 <= (&$signed($unsigned((reg230[(5'h14):(4'he)] ?
                  {reg245} : (reg274 ? reg189 : reg251)))));
              reg308 = $unsigned({(!reg264[(2'h2):(1'h0)]),
                  $unsigned((reg233[(5'h12):(4'ha)] >>> ((7'h4a) && reg282))),
                  (+((reg233 * reg282) ?
                      reg189[(1'h0):(1'h0)] : (reg296 > (7'h41))))});
              reg309 <= reg209;
            end
        end
    end
  assign wire310 = reg293[(5'h11):(5'h10)];
  assign wire311 = {$unsigned($unsigned($signed((wire185 != reg196))))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1961
#(parameter param2320 = (((~|((~(8'hac)) ? (^~(7'h54)) : (7'h54))) ? {((!(8'ha0)) ? (7'h4e) : {(8'ha7)}), {((8'hb6) ^~ (7'h50)), {(8'hbd), (7'h52)}}, (!(-(8'haf)))} : (!(((7'h4a) <= (8'hba)) == {(7'h55), (7'h4d), (8'hb6)}))) ? (~&((((8'hb3) > (8'h9e)) <<< {(7'h52), (7'h57)}) ? (~((7'h47) ? (8'ha4) : (8'hb0))) : {((8'h9e) >> (7'h49)), {(8'ha8), (8'haf)}})) : ((^~({(8'hbf), (8'h9f), (8'hb8)} || ((8'hbb) || (7'h4c)))) ? (!(!{(7'h55)})) : ((~{(8'hb1), (7'h57)}) != ({(7'h4b), (8'ha0), (7'h41)} ? {(8'ha7), (8'hb8), (7'h4c)} : ((8'hae) ? (7'h55) : (7'h54)))))))
(y, clk, wire1966, wire1965, wire1964, wire1963, wire1962);
  output wire [(32'h17ad):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire1966;
  input wire signed [(5'h18):(1'h0)] wire1965;
  input wire [(3'h6):(1'h0)] wire1964;
  input wire signed [(5'h18):(1'h0)] wire1963;
  input wire signed [(3'h7):(1'h0)] wire1962;
  wire [(2'h2):(1'h0)] wire2213;
  wire [(3'h4):(1'h0)] wire2212;
  wire [(4'hf):(1'h0)] wire2211;
  wire [(2'h3):(1'h0)] wire2210;
  wire signed [(5'h13):(1'h0)] wire2209;
  wire signed [(5'h15):(1'h0)] wire1967;
  reg [(5'h17):(1'h0)] reg2319 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2318 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2317 = (1'h0);
  reg [(4'h8):(1'h0)] reg2316 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2314 = (1'h0);
  reg [(3'h5):(1'h0)] reg2311 = (1'h0);
  reg [(4'h8):(1'h0)] reg2309 = (1'h0);
  reg [(5'h10):(1'h0)] reg2307 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2305 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2304 = (1'h0);
  reg [(5'h18):(1'h0)] reg2303 = (1'h0);
  reg [(2'h3):(1'h0)] reg2301 = (1'h0);
  reg [(4'h8):(1'h0)] reg2299 = (1'h0);
  reg [(4'hc):(1'h0)] reg2292 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2291 = (1'h0);
  reg [(5'h12):(1'h0)] reg2290 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2288 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2286 = (1'h0);
  reg [(5'h19):(1'h0)] reg2280 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2279 = (1'h0);
  reg [(5'h13):(1'h0)] reg2276 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2274 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2270 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2267 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2264 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2263 = (1'h0);
  reg [(4'hb):(1'h0)] reg2262 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2260 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2258 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2257 = (1'h0);
  reg [(4'h9):(1'h0)] reg2255 = (1'h0);
  reg [(5'h13):(1'h0)] reg2253 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2252 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2250 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2249 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2247 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2239 = (1'h0);
  reg [(5'h19):(1'h0)] reg2238 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2230 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2225 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2221 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2219 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2215 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2208 = (1'h0);
  reg [(5'h18):(1'h0)] reg2206 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2202 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2200 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2194 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2189 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2187 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2185 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2182 = (1'h0);
  reg [(3'h4):(1'h0)] reg2180 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2177 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2173 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2171 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2169 = (1'h0);
  reg [(4'h8):(1'h0)] reg2164 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2160 = (1'h0);
  reg [(5'h10):(1'h0)] reg2159 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2157 = (1'h0);
  reg [(4'h9):(1'h0)] reg2155 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2153 = (1'h0);
  reg [(4'hb):(1'h0)] reg2143 = (1'h0);
  reg [(5'h13):(1'h0)] reg2151 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2150 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2146 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2145 = (1'h0);
  reg [(4'hc):(1'h0)] reg2144 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2142 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2141 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2139 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2137 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2136 = (1'h0);
  reg [(3'h4):(1'h0)] reg2133 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2132 = (1'h0);
  reg [(4'h8):(1'h0)] reg2131 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2130 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2129 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2128 = (1'h0);
  reg [(4'h9):(1'h0)] reg2126 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2125 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2123 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2121 = (1'h0);
  reg [(3'h7):(1'h0)] reg2120 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2119 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2117 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2115 = (1'h0);
  reg [(4'h9):(1'h0)] reg2113 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2112 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2110 = (1'h0);
  reg [(3'h7):(1'h0)] reg2109 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2107 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2106 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2105 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2104 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2102 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2098 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2097 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2092 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2091 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2088 = (1'h0);
  reg [(4'h8):(1'h0)] reg2083 = (1'h0);
  reg [(4'hb):(1'h0)] reg2081 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2079 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2078 = (1'h0);
  reg [(5'h13):(1'h0)] reg2074 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2073 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2071 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2070 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2066 = (1'h0);
  reg [(5'h12):(1'h0)] reg2063 = (1'h0);
  reg [(5'h15):(1'h0)] reg2062 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2061 = (1'h0);
  reg [(4'ha):(1'h0)] reg2059 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2058 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2056 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2055 = (1'h0);
  reg [(5'h16):(1'h0)] reg2053 = (1'h0);
  reg [(3'h7):(1'h0)] reg2052 = (1'h0);
  reg [(5'h15):(1'h0)] reg2050 = (1'h0);
  reg [(5'h11):(1'h0)] reg2045 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2042 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2041 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2040 = (1'h0);
  reg [(5'h15):(1'h0)] reg2039 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2034 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2029 = (1'h0);
  reg [(3'h5):(1'h0)] reg2036 = (1'h0);
  reg [(3'h5):(1'h0)] reg2035 = (1'h0);
  reg [(5'h12):(1'h0)] reg2032 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2031 = (1'h0);
  reg [(5'h11):(1'h0)] reg2028 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2027 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2022 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2021 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2018 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2016 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2014 = (1'h0);
  reg [(4'hc):(1'h0)] reg2011 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2010 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1985 = (1'h0);
  reg [(5'h15):(1'h0)] reg2007 = (1'h0);
  reg [(2'h3):(1'h0)] reg2003 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2002 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1999 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1998 = (1'h0);
  reg [(4'hc):(1'h0)] reg1996 = (1'h0);
  reg [(5'h17):(1'h0)] reg1995 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1994 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1989 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1988 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1982 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1981 = (1'h0);
  reg [(5'h16):(1'h0)] reg1980 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1979 = (1'h0);
  reg [(4'he):(1'h0)] reg1978 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1976 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1973 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1971 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1970 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1969 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2312 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2315 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2313 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2312 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2310 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2308 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2306 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2302 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2300 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar2298 = (1'h0);
  reg [(5'h16):(1'h0)] reg2297 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2296 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2295 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2294 = (1'h0);
  reg [(4'hd):(1'h0)] reg2293 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2289 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2287 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2285 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2284 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2283 = (1'h0);
  reg [(2'h3):(1'h0)] reg2282 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2273 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2281 = (1'h0);
  reg [(3'h6):(1'h0)] reg2278 = (1'h0);
  reg [(4'hb):(1'h0)] reg2277 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2275 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2273 = (1'h0);
  reg [(5'h12):(1'h0)] reg2272 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2271 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2269 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2268 = (1'h0);
  reg [(3'h6):(1'h0)] reg2266 = (1'h0);
  reg [(5'h18):(1'h0)] reg2265 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2261 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2259 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2256 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2254 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2251 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2241 = (1'h0);
  reg [(3'h5):(1'h0)] reg2240 = (1'h0);
  reg [(5'h11):(1'h0)] reg2248 = (1'h0);
  reg [(5'h12):(1'h0)] reg2246 = (1'h0);
  reg [(5'h10):(1'h0)] reg2245 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2244 = (1'h0);
  reg [(5'h16):(1'h0)] reg2243 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2242 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2241 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2240 = (1'h0);
  reg [(4'h8):(1'h0)] reg2237 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2236 = (1'h0);
  reg [(2'h3):(1'h0)] reg2235 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2234 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2233 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2232 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2231 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2229 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2228 = (1'h0);
  reg [(3'h5):(1'h0)] reg2227 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2226 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2224 = (1'h0);
  reg [(5'h19):(1'h0)] reg2223 = (1'h0);
  reg [(5'h19):(1'h0)] reg2222 = (1'h0);
  reg [(5'h11):(1'h0)] reg2220 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2218 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar2217 = (1'h0);
  reg [(5'h18):(1'h0)] reg2216 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2214 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2207 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2205 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2204 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2203 = (1'h0);
  reg [(4'h9):(1'h0)] reg2201 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2199 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2198 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2197 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2196 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2195 = (1'h0);
  reg [(5'h11):(1'h0)] reg2193 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2192 = (1'h0);
  reg [(4'hd):(1'h0)] reg2191 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar2190 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2188 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2187 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2186 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2184 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2183 = (1'h0);
  reg [(4'hc):(1'h0)] reg2181 = (1'h0);
  reg [(4'hf):(1'h0)] reg2179 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2178 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2176 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2175 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2174 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2172 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2170 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2168 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2158 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2167 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2166 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2165 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2163 = (1'h0);
  reg [(2'h2):(1'h0)] reg2162 = (1'h0);
  reg [(5'h15):(1'h0)] reg2161 = (1'h0);
  reg [(5'h16):(1'h0)] reg2158 = (1'h0);
  reg [(4'hf):(1'h0)] reg2156 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2154 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2152 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2141 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2149 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2148 = (1'h0);
  reg [(4'ha):(1'h0)] reg2147 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2143 = (1'h0);
  reg [(3'h4):(1'h0)] reg2140 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2138 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2135 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2134 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2127 = (1'h0);
  reg [(4'h8):(1'h0)] reg2124 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2122 = (1'h0);
  reg [(5'h16):(1'h0)] reg2118 = (1'h0);
  reg [(3'h7):(1'h0)] reg2116 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2114 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2111 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2108 = (1'h0);
  reg [(5'h18):(1'h0)] reg2103 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2101 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2100 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2099 = (1'h0);
  reg [(4'h9):(1'h0)] reg2096 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2095 = (1'h0);
  reg [(5'h11):(1'h0)] reg2094 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2093 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2090 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2089 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2087 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar2086 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2085 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2084 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2082 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2069 = (1'h0);
  reg [(4'hd):(1'h0)] reg2080 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2077 = (1'h0);
  reg [(4'ha):(1'h0)] reg2076 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2075 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2072 = (1'h0);
  reg [(4'he):(1'h0)] reg2069 = (1'h0);
  reg [(4'h9):(1'h0)] reg2068 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2067 = (1'h0);
  reg [(4'hc):(1'h0)] reg2065 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2064 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2060 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2057 = (1'h0);
  reg [(3'h5):(1'h0)] reg2054 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2051 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2049 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2048 = (1'h0);
  reg [(5'h15):(1'h0)] reg2047 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2046 = (1'h0);
  reg [(3'h7):(1'h0)] reg2044 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2043 = (1'h0);
  reg [(4'ha):(1'h0)] reg2038 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2037 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2032 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2034 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2033 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2030 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2029 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2026 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2025 = (1'h0);
  reg [(3'h4):(1'h0)] reg2024 = (1'h0);
  reg [(2'h2):(1'h0)] reg2023 = (1'h0);
  reg [(4'ha):(1'h0)] reg2008 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2020 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2019 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2017 = (1'h0);
  reg [(4'h8):(1'h0)] reg2015 = (1'h0);
  reg [(2'h3):(1'h0)] reg2013 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2012 = (1'h0);
  reg [(5'h10):(1'h0)] reg2009 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2008 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2006 = (1'h0);
  reg [(3'h5):(1'h0)] reg2005 = (1'h0);
  reg [(4'h9):(1'h0)] reg2004 = (1'h0);
  reg [(2'h3):(1'h0)] reg2001 = (1'h0);
  reg [(5'h19):(1'h0)] reg2000 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1997 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1993 = (1'h0);
  reg [(3'h5):(1'h0)] reg1992 = (1'h0);
  reg [(5'h10):(1'h0)] reg1991 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1990 = (1'h0);
  reg [(5'h14):(1'h0)] reg1987 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1986 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1985 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1984 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1983 = (1'h0);
  reg [(5'h19):(1'h0)] reg1977 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1975 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1974 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1972 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1968 = (1'h0);
  assign y = {wire2213,
                 wire2212,
                 wire2211,
                 wire2210,
                 wire2209,
                 wire1967,
                 reg2319,
                 reg2318,
                 reg2317,
                 reg2316,
                 reg2314,
                 reg2311,
                 reg2309,
                 reg2307,
                 reg2305,
                 reg2304,
                 reg2303,
                 reg2301,
                 reg2299,
                 reg2292,
                 reg2291,
                 reg2290,
                 reg2288,
                 reg2286,
                 reg2280,
                 reg2279,
                 reg2276,
                 reg2274,
                 reg2270,
                 reg2267,
                 reg2264,
                 reg2263,
                 reg2262,
                 reg2260,
                 reg2258,
                 reg2257,
                 reg2255,
                 reg2253,
                 reg2252,
                 reg2250,
                 reg2249,
                 reg2247,
                 reg2239,
                 reg2238,
                 reg2230,
                 reg2225,
                 reg2221,
                 reg2219,
                 reg2215,
                 reg2208,
                 reg2206,
                 reg2202,
                 reg2200,
                 reg2194,
                 reg2189,
                 reg2187,
                 reg2185,
                 reg2182,
                 reg2180,
                 reg2177,
                 reg2173,
                 reg2171,
                 reg2169,
                 reg2164,
                 reg2160,
                 reg2159,
                 reg2157,
                 reg2155,
                 reg2153,
                 reg2143,
                 reg2151,
                 reg2150,
                 reg2146,
                 reg2145,
                 reg2144,
                 reg2142,
                 reg2141,
                 reg2139,
                 reg2137,
                 reg2136,
                 reg2133,
                 reg2132,
                 reg2131,
                 reg2130,
                 reg2129,
                 reg2128,
                 reg2126,
                 reg2125,
                 reg2123,
                 reg2121,
                 reg2120,
                 reg2119,
                 reg2117,
                 reg2115,
                 reg2113,
                 reg2112,
                 reg2110,
                 reg2109,
                 reg2107,
                 reg2106,
                 reg2105,
                 reg2104,
                 reg2102,
                 reg2098,
                 reg2097,
                 reg2092,
                 reg2091,
                 reg2088,
                 reg2083,
                 reg2081,
                 reg2079,
                 reg2078,
                 reg2074,
                 reg2073,
                 reg2071,
                 reg2070,
                 reg2066,
                 reg2063,
                 reg2062,
                 reg2061,
                 reg2059,
                 reg2058,
                 reg2056,
                 reg2055,
                 reg2053,
                 reg2052,
                 reg2050,
                 reg2045,
                 reg2042,
                 reg2041,
                 reg2040,
                 reg2039,
                 reg2034,
                 reg2029,
                 reg2036,
                 reg2035,
                 reg2032,
                 reg2031,
                 reg2028,
                 reg2027,
                 reg2022,
                 reg2021,
                 reg2018,
                 reg2016,
                 reg2014,
                 reg2011,
                 reg2010,
                 reg1985,
                 reg2007,
                 reg2003,
                 reg2002,
                 reg1999,
                 reg1998,
                 reg1996,
                 reg1995,
                 reg1994,
                 reg1989,
                 reg1988,
                 reg1982,
                 reg1981,
                 reg1980,
                 reg1979,
                 reg1978,
                 reg1976,
                 reg1973,
                 reg1971,
                 reg1970,
                 reg1969,
                 forvar2312,
                 reg2315,
                 reg2313,
                 reg2312,
                 reg2310,
                 reg2308,
                 reg2306,
                 reg2302,
                 reg2300,
                 forvar2298,
                 reg2297,
                 forvar2296,
                 reg2295,
                 reg2294,
                 reg2293,
                 reg2289,
                 reg2287,
                 reg2285,
                 forvar2284,
                 forvar2283,
                 reg2282,
                 reg2273,
                 reg2281,
                 reg2278,
                 reg2277,
                 reg2275,
                 forvar2273,
                 reg2272,
                 reg2271,
                 reg2269,
                 reg2268,
                 reg2266,
                 reg2265,
                 reg2261,
                 reg2259,
                 forvar2256,
                 reg2254,
                 reg2251,
                 forvar2241,
                 reg2240,
                 reg2248,
                 reg2246,
                 reg2245,
                 reg2244,
                 reg2243,
                 reg2242,
                 reg2241,
                 forvar2240,
                 reg2237,
                 reg2236,
                 reg2235,
                 forvar2234,
                 reg2233,
                 forvar2232,
                 forvar2231,
                 reg2229,
                 reg2228,
                 reg2227,
                 forvar2226,
                 reg2224,
                 reg2223,
                 reg2222,
                 reg2220,
                 reg2218,
                 forvar2217,
                 reg2216,
                 forvar2214,
                 reg2207,
                 forvar2205,
                 reg2204,
                 reg2203,
                 reg2201,
                 forvar2199,
                 forvar2198,
                 reg2197,
                 reg2196,
                 reg2195,
                 reg2193,
                 reg2192,
                 reg2191,
                 forvar2190,
                 reg2188,
                 forvar2187,
                 reg2186,
                 reg2184,
                 reg2183,
                 reg2181,
                 reg2179,
                 forvar2178,
                 reg2176,
                 reg2175,
                 reg2174,
                 reg2172,
                 reg2170,
                 forvar2168,
                 forvar2158,
                 reg2167,
                 reg2166,
                 reg2165,
                 reg2163,
                 reg2162,
                 reg2161,
                 reg2158,
                 reg2156,
                 reg2154,
                 reg2152,
                 forvar2141,
                 reg2149,
                 reg2148,
                 reg2147,
                 forvar2143,
                 reg2140,
                 reg2138,
                 reg2135,
                 forvar2134,
                 forvar2127,
                 reg2124,
                 reg2122,
                 reg2118,
                 reg2116,
                 forvar2114,
                 reg2111,
                 reg2108,
                 reg2103,
                 reg2101,
                 reg2100,
                 reg2099,
                 reg2096,
                 reg2095,
                 reg2094,
                 reg2093,
                 forvar2090,
                 reg2089,
                 reg2087,
                 forvar2086,
                 reg2085,
                 reg2084,
                 reg2082,
                 forvar2069,
                 reg2080,
                 reg2077,
                 reg2076,
                 reg2075,
                 reg2072,
                 reg2069,
                 reg2068,
                 reg2067,
                 reg2065,
                 reg2064,
                 reg2060,
                 reg2057,
                 reg2054,
                 reg2051,
                 reg2049,
                 reg2048,
                 reg2047,
                 reg2046,
                 reg2044,
                 reg2043,
                 reg2038,
                 reg2037,
                 forvar2032,
                 forvar2034,
                 reg2033,
                 reg2030,
                 forvar2029,
                 reg2026,
                 reg2025,
                 reg2024,
                 reg2023,
                 reg2008,
                 reg2020,
                 reg2019,
                 reg2017,
                 reg2015,
                 reg2013,
                 reg2012,
                 reg2009,
                 forvar2008,
                 reg2006,
                 reg2005,
                 reg2004,
                 reg2001,
                 reg2000,
                 reg1997,
                 reg1993,
                 reg1992,
                 reg1991,
                 reg1990,
                 reg1987,
                 reg1986,
                 forvar1985,
                 reg1984,
                 reg1983,
                 reg1977,
                 reg1975,
                 reg1974,
                 reg1972,
                 reg1968,
                 (1'h0)};
  assign wire1967 = wire1962;
  always
    @(posedge clk) begin
      if (wire1965[(3'h5):(2'h2)])
        begin
          if (wire1964[(1'h0):(1'h0)])
            begin
              reg1968 = (wire1962 ? wire1967 : wire1966);
              reg1969 <= $unsigned((+($unsigned(((7'h41) ?
                  wire1966 : reg1968)) >= {{wire1963},
                  (+wire1963),
                  (&wire1963)})));
              reg1970 <= {(wire1966[(1'h1):(1'h1)] == (wire1963 != (~&$unsigned(wire1966)))),
                  ($signed(((wire1967 ? wire1962 : wire1964) ^ wire1962)) ?
                      wire1963[(5'h13):(4'hf)] : (wire1967[(3'h7):(3'h7)] ?
                          (^~(wire1962 >> wire1965)) : $signed((reg1968 ?
                              reg1968 : reg1968)))),
                  wire1964};
              reg1971 <= {(8'ha9), reg1970, (7'h41)};
            end
          else
            begin
              reg1969 <= (~|$unsigned($unsigned($signed((reg1970 != reg1970)))));
              reg1970 <= (~^reg1968[(2'h3):(2'h3)]);
              reg1971 <= reg1970[(5'h1b):(5'h17)];
              reg1972 = (+({(reg1969[(5'h10):(5'h10)] != wire1967),
                  $signed($signed(reg1968))} << $signed(wire1967[(1'h1):(1'h0)])));
            end
          reg1973 <= $signed($signed((~|$signed((reg1970 ?
              reg1968 : reg1969)))));
        end
      else
        begin
          reg1969 <= reg1972[(3'h5):(3'h5)];
          reg1972 = ({reg1972[(3'h7):(1'h0)],
              $signed(reg1972[(4'h9):(3'h7)]),
              reg1970[(5'h12):(4'h8)]} >> (~|reg1970[(5'h16):(4'h9)]));
          if (((^reg1968) ?
              wire1962 : $unsigned(($unsigned((wire1965 & wire1964)) ?
                  (^~(reg1971 - wire1967)) : ((wire1965 - wire1965) ?
                      wire1963[(4'hd):(4'h8)] : {(8'hbb),
                          reg1970,
                          wire1965})))))
            begin
              reg1973 <= reg1968[(3'h4):(2'h2)];
              reg1974 = ($signed(reg1969[(3'h4):(2'h2)]) ^~ ((|wire1963[(4'hc):(2'h3)]) && (((|reg1969) <<< wire1965) <<< $signed((wire1964 - wire1967)))));
              reg1975 = {(!wire1963), reg1971};
            end
          else
            begin
              reg1973 <= ($signed($signed(wire1962)) ?
                  ((|$signed((|reg1974))) ?
                      wire1967[(5'h11):(3'h7)] : $signed((~reg1968))) : $signed((reg1968 <<< $signed((|wire1967)))));
              reg1976 <= (reg1969 ^ (~reg1970[(5'h1b):(4'hb)]));
              reg1977 = (wire1967 ^ $signed({reg1976,
                  reg1970[(5'h15):(2'h3)]}));
            end
          if ($signed((((reg1970[(4'hc):(4'hb)] > $unsigned(reg1975)) ?
                  (^~(8'hab)) : $signed(wire1964[(1'h0):(1'h0)])) ?
              reg1976[(1'h1):(1'h0)] : ($unsigned((reg1969 ?
                  reg1974 : (8'ha7))) - $unsigned((reg1971 ?
                  wire1966 : wire1963))))))
            begin
              reg1978 <= {((reg1974[(2'h3):(2'h3)] ?
                      (~&$unsigned(wire1964)) : $signed(wire1965[(3'h4):(2'h2)])) < ($signed(wire1965[(5'h11):(4'hc)]) ?
                      $unsigned((^(8'had))) : ({reg1974, wire1965} ?
                          reg1976[(5'h1d):(3'h5)] : (reg1971 == (8'ha1))))),
                  reg1971[(5'h15):(5'h15)],
                  ((&((wire1965 & reg1968) ?
                          $unsigned((7'h56)) : $signed((7'h54)))) ?
                      ((-(wire1963 | wire1965)) ?
                          (~wire1965) : (^$unsigned((8'hb1)))) : (reg1977[(5'h10):(1'h1)] ?
                          $signed($unsigned(wire1963)) : (reg1977 ?
                              (reg1973 ? wire1966 : reg1972) : (&reg1969))))};
              reg1979 <= (($signed(($unsigned(reg1978) ?
                      (|reg1978) : (8'hba))) ?
                  (((reg1978 ^~ reg1970) ?
                          wire1966[(4'ha):(4'h8)] : $unsigned(reg1972)) ?
                      reg1968 : $signed((reg1971 == reg1973))) : {{$signed(reg1972)},
                      reg1976}) + (reg1970 + (($signed(reg1977) <<< $signed(reg1976)) ?
                  reg1974 : (8'haf))));
              reg1980 <= ($signed(($signed({wire1964,
                  (8'ha8)}) >> $unsigned(reg1979[(4'he):(4'hc)]))) <<< reg1975);
              reg1981 <= reg1974;
              reg1982 <= $signed(reg1980[(3'h5):(1'h0)]);
              reg1983 = reg1981;
            end
          else
            begin
              reg1978 <= (reg1976 <<< {reg1974[(1'h0):(1'h0)],
                  ((reg1978 ^~ (~|reg1976)) ? (~&$signed(reg1969)) : wire1964),
                  $signed(wire1966[(1'h0):(1'h0)])});
            end
        end
      if (reg1974)
        begin
          reg1984 = reg1975;
          for (forvar1985 = (1'h0); (forvar1985 < (3'h6)); forvar1985 = (forvar1985 + (1'h1)))
            begin
              reg1986 = $signed((((~&forvar1985) >> {$unsigned(reg1968),
                      reg1974}) ?
                  wire1963[(3'h6):(3'h6)] : $signed(((reg1982 ?
                      wire1966 : reg1972) && reg1970[(4'he):(2'h3)]))));
              reg1987 = $signed(({(reg1976 <= reg1973),
                      ((reg1974 ? reg1976 : wire1962) ^~ $signed(reg1971))} ?
                  ($unsigned((wire1964 ?
                      reg1974 : reg1979)) - $signed((reg1976 <= wire1962))) : reg1979));
              reg1988 <= $unsigned($unsigned($signed({reg1976[(4'hc):(2'h2)],
                  $unsigned((7'h47))})));
              reg1989 <= (!(reg1971[(2'h3):(2'h3)] ?
                  wire1963[(4'h8):(3'h6)] : reg1983[(2'h3):(2'h3)]));
              reg1990 = $signed(((({reg1987} ? reg1971 : (wire1963 ^ reg1977)) ?
                  ((reg1980 << reg1980) <= (reg1978 ?
                      reg1974 : reg1989)) : $unsigned(reg1978[(3'h5):(3'h4)])) | wire1963[(4'h8):(4'h8)]));
              reg1991 = reg1989;
              reg1992 = $unsigned(($signed(($signed(reg1971) ?
                  {(7'h48), reg1970, (8'hb0)} : (~|reg1975))) >> ({(^reg1988),
                      $signed(reg1990)} ?
                  reg1970[(4'h8):(2'h2)] : reg1977)));
            end
          if ((+reg1972[(1'h1):(1'h0)]))
            begin
              reg1993 = wire1966;
              reg1994 <= {((reg1968[(1'h1):(1'h1)] ?
                      ($signed((8'hb8)) ?
                          (reg1972 ?
                              forvar1985 : reg1988) : (wire1967 >> reg1970)) : reg1991) ^ {(7'h55),
                      $unsigned((reg1976 | wire1964)),
                      reg1973})};
              reg1995 <= reg1978;
              reg1996 <= reg1980;
            end
          else
            begin
              reg1993 = reg1981[(5'h15):(4'h9)];
              reg1997 = $signed((reg1980[(5'h16):(3'h5)] && $unsigned(($unsigned(reg1990) ?
                  wire1967[(3'h5):(1'h0)] : ((7'h43) ? reg1979 : reg1980)))));
              reg1998 <= (((((forvar1985 ? reg1990 : reg1994) ?
                      reg1980[(3'h4):(2'h3)] : wire1962) ~^ $signed(wire1962)) == {(reg1995 ?
                          $signed(reg1974) : $unsigned(reg1974))}) ?
                  (~$unsigned((~^(reg1968 >= reg1993)))) : (^~(~^{reg1969})));
              reg1999 <= (reg1969[(5'h1c):(5'h12)] ?
                  (8'ha7) : (~^(({reg1989, reg1998} | (wire1965 - (8'had))) ?
                      (~^reg1979) : $unsigned((~|(8'h9f))))));
              reg2000 = $signed((~&(($unsigned(reg1974) >> (~^forvar1985)) >> ($unsigned(reg1994) | wire1963))));
            end
          if (reg1968)
            begin
              reg2001 = ((7'h4f) <= (reg1995 >> reg1992));
              reg2002 <= ((~|$signed({(wire1962 * wire1966),
                      $signed(reg1974)})) ?
                  {(wire1965[(4'ha):(1'h1)] != $unsigned($unsigned(reg1981)))} : (~&$signed({$unsigned(reg1991),
                      $unsigned(reg1996)})));
              reg2003 <= $unsigned((&$signed(((reg1994 || reg1981) ?
                  $unsigned(reg1986) : (reg1981 < reg1972)))));
              reg2004 = (!$signed((reg1993 ~^ $signed({wire1967,
                  (7'h4c),
                  reg1987}))));
              reg2005 = $signed({(((-reg1972) | ((8'ha3) >>> reg1984)) ?
                      $unsigned(reg2002) : $unsigned((reg1971 - reg1971)))});
              reg2006 = {reg1988[(5'h10):(3'h4)],
                  {(8'ha1), (+(|(reg1987 ? reg1999 : (8'ha5))))},
                  wire1963[(3'h7):(2'h2)]};
              reg2007 <= ((($signed($signed(reg1990)) << reg1992[(1'h1):(1'h0)]) || ($signed((reg1972 & reg1974)) ?
                  reg1974 : $unsigned(reg2006))) ~^ reg1980[(5'h15):(5'h10)]);
            end
          else
            begin
              reg2002 <= ($unsigned($unsigned($unsigned((reg1969 ?
                  wire1965 : reg1973)))) ^ $unsigned($signed(((&reg1997) ?
                  (reg2004 ? (8'ha0) : reg1994) : reg1996[(4'h8):(3'h5)]))));
            end
        end
      else
        begin
          reg1985 <= (~^(reg1968[(1'h0):(1'h0)] < {(reg1973[(5'h19):(4'hb)] ?
                  $signed(reg2002) : (reg2006 != reg1980)),
              (~&(reg1986 >= wire1965))}));
        end
      if (reg1993)
        begin
          for (forvar2008 = (1'h0); (forvar2008 < (1'h0)); forvar2008 = (forvar2008 + (1'h1)))
            begin
              reg2009 = $signed($signed($signed(({reg1976} ?
                  (reg2001 < wire1962) : (reg1968 || reg1972)))));
              reg2010 <= $unsigned(($signed(reg1985) * (((|wire1963) ?
                      (~(7'h51)) : reg1986[(4'ha):(3'h6)]) ?
                  (forvar1985[(4'h9):(3'h5)] ?
                      (reg1976 >>> reg1998) : $unsigned(reg2009)) : $signed($signed(wire1964)))));
              reg2011 <= reg1971[(5'h1b):(4'hf)];
              reg2012 = (^reg2011[(3'h7):(2'h2)]);
              reg2013 = (~^(wire1963[(4'hc):(1'h1)] < {$signed((reg1984 ?
                      reg1996 : reg1992)),
                  reg1991[(4'hf):(1'h0)],
                  reg1975}));
            end
          reg2014 <= reg2011[(3'h7):(3'h6)];
          if (reg2001)
            begin
              reg2015 = (($unsigned((^(reg2009 ?
                      reg1998 : wire1965))) > reg1989) ?
                  (((&(~&wire1963)) ?
                      (reg1971[(2'h2):(1'h0)] ?
                          (reg1976 ?
                              wire1962 : reg2012) : reg1983[(3'h6):(1'h0)]) : (reg2014 ?
                          (wire1963 ? reg1968 : reg1985) : (reg1997 ?
                              reg1983 : reg1996))) | $unsigned({(8'ha2)})) : forvar1985[(5'h13):(2'h2)]);
              reg2016 <= {(!{{reg1975, {reg1990}}}),
                  reg1982,
                  ($signed($unsigned((~|(8'hac)))) << (($signed(forvar1985) ?
                          forvar1985 : wire1967) ?
                      {reg1968, (reg2002 ? reg2004 : reg1984)} : (-{reg2002,
                          (8'hb1)})))};
              reg2017 = ({((^~(reg2015 != (8'h9e))) || ((!reg2006) ~^ $unsigned(reg1997))),
                  $signed(reg2011)} ^~ $signed($unsigned(reg1997)));
              reg2018 <= $signed(reg2013);
            end
          else
            begin
              reg2015 = $unsigned(reg2017[(3'h7):(3'h4)]);
              reg2017 = ({reg1981[(5'h16):(2'h3)],
                  {(~|$unsigned(wire1967))}} != (~(wire1965[(2'h2):(1'h1)] ?
                  (reg1984[(2'h3):(2'h3)] ?
                      (8'h9f) : reg1995[(2'h2):(2'h2)]) : (8'ha8))));
              reg2018 <= wire1963[(2'h2):(1'h0)];
              reg2019 = $signed($unsigned((reg1989 > (&reg1975[(3'h5):(2'h3)]))));
            end
          reg2020 = reg2016;
        end
      else
        begin
          if ((~(((8'ha2) ?
              $signed((reg2014 ?
                  reg1971 : reg2006)) : (|reg1978)) <= (($unsigned(reg1982) >> (reg2012 ~^ reg1993)) ?
              reg1982[(2'h2):(1'h0)] : $unsigned(reg1996[(4'h9):(3'h7)])))))
            begin
              reg2008 = {$signed($unsigned(wire1964[(3'h4):(3'h4)])),
                  ($unsigned({(-reg2011)}) ?
                      $signed(reg2004[(3'h6):(1'h1)]) : (8'hba))};
              reg2009 = ((~$signed($signed(reg1989))) ?
                  {$unsigned((reg2003 ?
                          (wire1962 ?
                              reg1984 : reg1978) : (8'ha7)))} : reg1971);
              reg2010 <= reg1980[(4'hd):(1'h1)];
            end
          else
            begin
              reg2010 <= reg1980;
              reg2012 = ((reg2010[(4'he):(1'h1)] ?
                  $unsigned($unsigned((reg1997 < reg1983))) : $unsigned(wire1965)) ^~ (~&((reg1993 ?
                      $signed(wire1966) : reg2011) ?
                  ($unsigned(reg1987) ?
                      (~wire1963) : (~^forvar1985)) : {(reg2005 * (8'hbf)),
                      (reg1979 ~^ reg2017),
                      reg1983})));
              reg2014 <= $unsigned($unsigned(reg1989[(3'h6):(1'h1)]));
              reg2016 <= $unsigned($unsigned((-$unsigned({reg2012,
                  (7'h57),
                  (7'h43)}))));
              reg2017 = ({reg1987} ?
                  $unsigned((-$unsigned(reg1978))) : reg1975);
              reg2019 = ($signed(($signed((^~reg1969)) < {$unsigned(wire1966)})) != forvar2008);
              reg2020 = (|reg2016);
            end
          if ((reg1987 ?
              ((!(reg1982 ?
                  (wire1962 ?
                      reg1977 : reg1989) : {(8'ha8)})) - (8'ha5)) : $signed((!(!reg1981)))))
            begin
              reg2021 <= reg1999[(5'h1c):(4'hb)];
              reg2022 <= reg1996;
              reg2023 = reg2000[(5'h19):(4'hc)];
              reg2024 = reg1979[(1'h1):(1'h1)];
              reg2025 = $signed((!reg1995));
              reg2026 = ((&(8'ha4)) || (~$unsigned(($signed(reg1997) > reg2000[(2'h2):(2'h2)]))));
            end
          else
            begin
              reg2021 <= (reg1978 > ((reg2000[(4'h8):(3'h5)] - {(reg2004 - reg2005),
                  (8'ha8)}) >>> reg2020[(3'h4):(1'h1)]));
              reg2023 = ((-$unsigned((((8'ha2) >= reg1976) << reg2018[(1'h1):(1'h0)]))) ~^ reg2016[(4'h9):(2'h3)]);
              reg2024 = (reg1996 >> (reg1977[(5'h12):(2'h3)] ?
                  (^~$signed((reg1987 > reg1982))) : $unsigned((~&$unsigned(reg2009)))));
              reg2025 = (~|$unsigned(reg1969));
            end
          reg2027 <= (!wire1965[(4'hc):(3'h6)]);
        end
      if (reg2023[(1'h1):(1'h0)])
        begin
          reg2028 <= $signed(reg2015[(3'h5):(3'h4)]);
          for (forvar2029 = (1'h0); (forvar2029 < (3'h6)); forvar2029 = (forvar2029 + (1'h1)))
            begin
              reg2030 = $unsigned(wire1965[(5'h17):(4'hb)]);
              reg2031 <= $unsigned(reg2025);
              reg2032 <= $signed(reg1992);
            end
          reg2033 = $unsigned(reg1983[(3'h5):(2'h2)]);
          for (forvar2034 = (1'h0); (forvar2034 < (1'h1)); forvar2034 = (forvar2034 + (1'h1)))
            begin
              reg2035 <= reg1982;
              reg2036 <= (~|(|$signed($unsigned(reg2004))));
            end
        end
      else
        begin
          reg2028 <= $signed({(~^(forvar2034 ?
                  $unsigned(reg1983) : (forvar1985 ? reg2000 : reg1996)))});
          if ((~^(|wire1965[(4'ha):(4'h8)])))
            begin
              reg2029 <= {(reg2001[(1'h0):(1'h0)] ?
                      reg2021[(1'h0):(1'h0)] : reg2005),
                  $unsigned(reg1978[(2'h3):(1'h1)])};
              reg2030 = (~^wire1965);
              reg2031 <= ($unsigned(reg1974[(5'h12):(4'he)]) ?
                  (7'h4e) : (reg2024 ?
                      ((7'h46) ?
                          reg1979 : reg1979[(3'h6):(3'h4)]) : (|reg1971)));
            end
          else
            begin
              reg2029 <= (8'hae);
            end
          for (forvar2032 = (1'h0); (forvar2032 < (1'h0)); forvar2032 = (forvar2032 + (1'h1)))
            begin
              reg2034 <= $unsigned($unsigned({$unsigned((~&reg1996)),
                  $unsigned($unsigned((7'h45)))}));
              reg2035 <= reg1998;
              reg2037 = (reg2015 ?
                  reg1994[(5'h15):(3'h5)] : $signed($unsigned(({reg2020,
                      reg2013,
                      wire1966} & (reg2019 ~^ (8'hb0))))));
              reg2038 = (!$unsigned((&$unsigned(reg2016))));
              reg2039 <= reg1988[(4'ha):(4'h9)];
              reg2040 <= reg1970[(4'ha):(3'h6)];
            end
          reg2041 <= $unsigned($signed(reg2036));
          if ({((~reg2027[(2'h2):(1'h1)]) ?
                  (((reg1988 ? reg2008 : reg2013) >> ((8'hbb) ?
                          reg1972 : reg1991)) ?
                      ((reg2001 != reg1986) ?
                          (reg1977 ?
                              reg1984 : reg2013) : (-reg1998)) : {((7'h46) ?
                              reg1998 : (8'hb5)),
                          (|reg1982),
                          reg1986[(5'h16):(3'h4)]}) : ((reg1982 ^ (forvar2008 ?
                      reg2004 : wire1965)) ^ ($unsigned(reg2017) ?
                      reg1973[(3'h6):(3'h5)] : $signed(reg2039))))})
            begin
              reg2042 <= reg1998;
              reg2043 = reg1976;
              reg2044 = (((~&(reg1976[(4'h9):(2'h3)] && $unsigned(forvar2034))) <= reg1992[(3'h4):(2'h3)]) ?
                  (reg1973[(4'h9):(3'h4)] ?
                      $unsigned(($signed(wire1965) ?
                          $unsigned((8'hba)) : $signed(reg1972))) : (~|(reg2039 ?
                          $signed(reg2029) : $signed((7'h47))))) : ((^~reg1993[(4'h9):(3'h5)]) == $signed($signed(reg1974))));
            end
          else
            begin
              reg2042 <= (~^reg1977[(3'h6):(3'h6)]);
              reg2043 = reg1981;
              reg2045 <= ($signed(((^(reg1975 == forvar2008)) ?
                  reg2013 : $unsigned((~^reg2021)))) != ((&reg1992) ?
                  ((|reg2001[(2'h3):(1'h0)]) >= $unsigned((wire1967 >= reg1996))) : reg1979));
              reg2046 = reg2040;
            end
          if (reg2016[(4'he):(3'h6)])
            begin
              reg2047 = $signed($unsigned(reg2011));
              reg2048 = $signed(($unsigned(($signed(reg2012) ^ $signed((8'hb6)))) ?
                  (8'h9c) : reg1990[(1'h1):(1'h0)]));
              reg2049 = (({$unsigned(reg1985[(5'h1b):(3'h5)])} ?
                  $unsigned((7'h49)) : (~{$signed((7'h41))})) >= (reg1980[(3'h7):(3'h7)] <= ($signed(reg1999) ?
                  {$signed(reg2015),
                      reg1975,
                      $unsigned(reg2018)} : reg2009[(4'h8):(2'h3)])));
              reg2050 <= reg2028;
              reg2051 = forvar1985;
              reg2052 <= $unsigned(reg1979[(5'h15):(4'ha)]);
            end
          else
            begin
              reg2047 = (reg2006[(3'h6):(1'h0)] ?
                  reg1990 : ((~^{{reg2008, (8'ha5), reg1988},
                          (reg2039 ? (8'ha4) : (8'hb8)),
                          reg1989[(3'h5):(1'h0)]}) ?
                      reg1982[(4'h9):(4'h8)] : {({reg2004, reg2025, reg2044} ?
                              $signed(reg2028) : (~reg2051)),
                          reg1975[(5'h18):(4'h8)],
                          ($unsigned(reg2015) ?
                              reg1992[(2'h3):(2'h3)] : (reg2031 && (7'h55)))}));
              reg2050 <= ($signed(reg1989) ^ reg1998[(3'h5):(3'h5)]);
              reg2051 = $unsigned({(^{$unsigned(reg1969)}),
                  $unsigned(((wire1964 ? reg1969 : reg1976) ?
                      (7'h53) : (reg2032 ? reg1987 : reg1979)))});
            end
        end
      reg2053 <= (({(~^reg1980),
                  ((^reg2034) ? $signed(reg2013) : forvar2032),
                  $signed(reg1993[(3'h5):(1'h0)])} ?
              {$signed($signed(reg2049))} : (+$unsigned(reg2016))) ?
          reg1994[(5'h14):(4'hf)] : (&reg2023));
      if (((7'h47) != reg2033))
        begin
          if ((~^($unsigned(((reg2004 ? reg2020 : reg1984) ?
              (&(8'hb7)) : (~&reg2013))) < reg1994[(5'h10):(4'h9)])))
            begin
              reg2054 = (-(~&($signed(reg2053) || ($unsigned(reg1976) + ((7'h44) ?
                  reg2009 : reg2048)))));
              reg2055 <= $signed($signed((reg2022[(5'h13):(4'hd)] + (7'h48))));
              reg2056 <= $unsigned({(((^~(7'h44)) ?
                          $signed(reg2038) : $unsigned(reg1975)) ?
                      {((8'hb7) ? wire1964 : reg2043),
                          $unsigned(reg2006),
                          (^(7'h56))} : {$signed(reg1985), $signed(reg2032)}),
                  ((((8'ha0) ? reg2040 : forvar2008) >>> reg2019) ?
                      ((reg2038 != reg1979) & reg2009[(4'hb):(3'h7)]) : (~^$unsigned(reg2024))),
                  $signed($signed(reg1999[(1'h1):(1'h0)]))});
              reg2057 = (&{(wire1967 ?
                      (|{(7'h57), reg2007}) : $signed((reg2031 == (7'h45)))),
                  $signed(((reg2019 ? reg1988 : reg2027) ?
                      wire1963[(5'h10):(4'h8)] : reg2027)),
                  (reg2035 ? (!reg2010) : ($signed(reg1986) ~^ (^~reg2045)))});
              reg2058 <= reg2042;
              reg2059 <= (reg2014 < ((reg2010 ^~ (+(~(8'h9d)))) > (+forvar1985)));
            end
          else
            begin
              reg2055 <= (|$signed($unsigned(wire1966[(1'h1):(1'h0)])));
              reg2056 <= {$unsigned({$signed($unsigned((7'h48))),
                      $unsigned($signed(reg2023))}),
                  (~^(^~$signed(reg2041))),
                  reg2047};
              reg2058 <= (~&$signed($unsigned(reg1986[(5'h13):(4'h8)])));
              reg2059 <= reg1975;
              reg2060 = $signed($signed({($unsigned(reg2024) ?
                      forvar2032 : (reg2043 | reg1998)),
                  reg1981[(5'h19):(4'h9)]}));
            end
          reg2061 <= reg2036[(3'h5):(3'h4)];
        end
      else
        begin
          if ((+(reg1998[(3'h5):(3'h4)] ^ $unsigned({reg1983[(3'h5):(3'h4)],
              reg2034}))))
            begin
              reg2054 = ($unsigned(reg1970) | (|{(~$unsigned(reg2005))}));
              reg2055 <= wire1967[(5'h10):(3'h7)];
            end
          else
            begin
              reg2055 <= $signed($unsigned($unsigned($unsigned({reg2023}))));
            end
          reg2056 <= $signed($signed(reg2042));
          if ((~&(($signed(reg2025[(2'h2):(1'h1)]) ?
                  (((7'h42) ~^ (8'hb2)) ?
                      $unsigned(reg2025) : reg2047[(5'h13):(5'h11)]) : $signed((|wire1966))) ?
              ($signed(((8'hab) >>> reg1979)) - {reg2028,
                  reg2042,
                  $unsigned((7'h58))}) : reg2045[(4'hb):(3'h7)])))
            begin
              reg2058 <= (reg2017[(3'h7):(2'h3)] ?
                  reg2012[(1'h0):(1'h0)] : wire1967);
              reg2059 <= (((wire1965 ?
                  reg1972[(2'h2):(1'h1)] : (|reg2037[(3'h7):(3'h4)])) | (&$signed($unsigned(reg2009)))) ~^ reg1988[(4'h8):(1'h1)]);
              reg2061 <= ((&$signed({(!reg1974),
                  $signed(wire1963),
                  reg1988})) <= (|reg2026));
              reg2062 <= (reg2058 ^ (^reg2053));
              reg2063 <= (+$signed($unsigned($signed($signed(forvar2029)))));
            end
          else
            begin
              reg2057 = $signed((forvar2029 ?
                  (7'h43) : $unsigned({reg1982[(4'h9):(3'h6)],
                      reg2014,
                      (reg1991 ? reg1976 : (8'h9c))})));
              reg2060 = $signed($unsigned(reg2053[(4'he):(1'h1)]));
              reg2064 = forvar2029[(5'h13):(4'ha)];
              reg2065 = reg2042[(4'hc):(4'hb)];
            end
          reg2066 <= $signed(reg2041[(3'h7):(1'h1)]);
          reg2067 = $unsigned($signed((-(7'h4b))));
        end
    end
  always
    @(posedge clk) begin
      reg2068 = ((-(~$unsigned((reg2061 ? reg1999 : reg2007)))) ^ wire1966);
      if ($signed((wire1965 * reg2032)))
        begin
          if ($unsigned((reg2058[(2'h2):(2'h2)] >> $signed(($signed(reg2056) | {reg2031,
              reg2029,
              (8'hb4)})))))
            begin
              reg2069 = reg2022[(5'h10):(4'hf)];
            end
          else
            begin
              reg2069 = ($unsigned(reg2021[(4'h8):(2'h2)]) ?
                  $unsigned(($unsigned($unsigned(reg1980)) > reg2055[(1'h1):(1'h1)])) : {$signed($unsigned($unsigned(reg2053))),
                      (reg1989[(2'h3):(1'h0)] <<< reg2022[(5'h12):(3'h7)])});
              reg2070 <= $unsigned((~&reg2069));
              reg2071 <= (8'ha7);
              reg2072 = (($signed($unsigned(wire1966)) ^ (!reg2028[(5'h11):(1'h0)])) && (&$unsigned($signed($unsigned(reg2016)))));
              reg2073 <= ((~^reg2070[(5'h1a):(4'ha)]) && $signed($signed({(8'hb7),
                  ((8'ha3) ~^ reg1970),
                  $unsigned(reg2018)})));
            end
          if ((($signed((reg1978 & $unsigned(reg1995))) ?
                  (^$signed((~^reg1980))) : (reg1989[(1'h1):(1'h0)] ?
                      ((reg2016 ? reg1971 : reg2035) ?
                          (reg2072 ?
                              reg1985 : wire1965) : wire1965[(5'h13):(3'h6)]) : wire1966[(1'h1):(1'h0)])) ?
              $signed((reg2028[(4'hd):(3'h6)] ?
                  ($unsigned(reg2036) ?
                      $signed(reg1985) : reg1973[(4'h9):(3'h5)]) : $unsigned(reg2007[(4'h9):(2'h3)]))) : {reg2052,
                  wire1964[(3'h4):(3'h4)]}))
            begin
              reg2074 <= reg2062[(4'ha):(4'h8)];
            end
          else
            begin
              reg2075 = $unsigned(reg1996[(3'h6):(1'h1)]);
              reg2076 = reg2069;
              reg2077 = {reg1981, reg2011};
              reg2078 <= (-(^~{reg2039[(5'h12):(4'hb)],
                  ((^~reg1969) >> (reg2002 >= (8'ha5))),
                  wire1964}));
              reg2079 <= (^~$signed((+reg2021)));
              reg2080 = (~(^~(($signed(reg1985) * ((7'h55) ?
                  (8'hbf) : reg2027)) <= $unsigned($unsigned(reg2078)))));
              reg2081 <= (((^$unsigned({reg2042, reg1998, reg1996})) ?
                  (^reg2058[(1'h1):(1'h1)]) : (^$signed($signed(reg1973)))) && {$signed(reg1980),
                  ($unsigned({wire1965}) ^~ {(~reg2075),
                      reg2071[(3'h4):(2'h2)]}),
                  $signed((7'h45))});
            end
        end
      else
        begin
          for (forvar2069 = (1'h0); (forvar2069 < (3'h4)); forvar2069 = (forvar2069 + (1'h1)))
            begin
              reg2072 = (-reg2068);
              reg2075 = reg2072[(4'ha):(2'h3)];
              reg2076 = ($signed(reg1985) | reg1996);
              reg2078 <= $unsigned(reg1976);
            end
          reg2080 = $unsigned({($unsigned(reg2071[(4'h8):(2'h3)]) ?
                  {(^(7'h4b))} : reg2040[(3'h7):(1'h0)]),
              $signed(reg2040[(2'h3):(2'h2)])});
          reg2081 <= $unsigned((|$unsigned(((reg2069 ?
              reg2002 : reg1998) < {wire1962, reg2031, reg2002}))));
          if ({((reg2058[(3'h4):(1'h0)] & $signed($unsigned(reg2081))) ?
                  {reg2016[(3'h4):(2'h2)],
                      reg1995[(4'hb):(3'h5)],
                      $signed((-reg2074))} : (-(!((7'h50) == reg2056))))})
            begin
              reg2082 = $unsigned(reg2075);
              reg2083 <= (7'h56);
            end
          else
            begin
              reg2082 = reg1970;
              reg2084 = reg2011[(4'h8):(4'h8)];
              reg2085 = $signed((({$unsigned(reg1973),
                      (reg2018 >> reg2039),
                      (reg2028 != wire1964)} == {(wire1963 ?
                          reg2032 : wire1965),
                      reg2061,
                      reg2062[(3'h7):(3'h5)]}) ?
                  (reg2036 ?
                      $unsigned((-reg2032)) : {$unsigned(reg2070),
                          reg2031,
                          (reg2039 & reg1994)}) : {reg1995[(5'h15):(4'hf)]}));
            end
          for (forvar2086 = (1'h0); (forvar2086 < (2'h3)); forvar2086 = (forvar2086 + (1'h1)))
            begin
              reg2087 = $unsigned($unsigned(reg2076));
            end
          reg2088 <= ($unsigned((7'h55)) ?
              ((^~(reg2039[(5'h10):(4'hd)] ^~ reg2068)) ?
                  $signed(((~|reg1971) ?
                      reg2077[(3'h5):(3'h4)] : (|reg2035))) : $unsigned(((wire1965 ^~ reg2056) ?
                      $signed(wire1966) : (forvar2086 >> wire1963)))) : reg2003[(1'h0):(1'h0)]);
        end
      reg2089 = {(+(^$signed($signed(reg2028)))),
          ((-$signed(reg2002[(1'h1):(1'h0)])) ~^ (~^(+reg1980)))};
      for (forvar2090 = (1'h0); (forvar2090 < (1'h0)); forvar2090 = (forvar2090 + (1'h1)))
        begin
          reg2091 <= reg2014;
          reg2092 <= (reg2076[(3'h6):(2'h3)] ?
              (((~^{reg2073, (8'hba), reg2071}) ?
                      $unsigned(reg2085[(5'h1e):(5'h14)]) : forvar2069[(3'h7):(3'h5)]) ?
                  (((7'h4c) >>> reg1998[(4'hb):(3'h7)]) ?
                      (~reg2041[(5'h1c):(5'h10)]) : reg1985[(3'h5):(1'h1)]) : reg1980[(1'h1):(1'h1)]) : reg2050);
          if (reg2070)
            begin
              reg2093 = $signed(wire1962);
              reg2094 = (($unsigned(($signed(reg2059) ?
                          $signed(reg2002) : reg2010)) ?
                      $signed(((~reg1969) & reg2083[(3'h5):(3'h5)])) : (&$signed($signed(reg2071)))) ?
                  {$signed(reg2031[(2'h2):(1'h0)])} : $signed((+$signed((reg2016 ?
                      forvar2086 : reg2084)))));
              reg2095 = reg2016;
              reg2096 = (8'hbf);
              reg2097 <= reg2077[(5'h18):(4'hd)];
            end
          else
            begin
              reg2093 = $signed(($unsigned(reg2032[(3'h5):(2'h3)]) < (($unsigned(reg2076) || wire1965[(4'he):(2'h2)]) ?
                  ($signed(reg2092) & {(7'h47), reg2042}) : reg2093)));
              reg2097 <= (reg1970[(1'h1):(1'h1)] * (({$signed(reg2053),
                  {reg2088, wire1962},
                  {reg2036,
                      reg2092}} >= $signed((8'hb0))) * (~|{(~|reg2052)})));
              reg2098 <= $signed(reg2094);
              reg2099 = reg2056;
              reg2100 = (8'haa);
              reg2101 = ($signed(reg2080[(4'h9):(3'h4)]) * (!((wire1966 ~^ (reg2029 ?
                      reg2088 : reg2056)) ?
                  (((7'h4f) | reg2039) ?
                      (~reg1971) : reg1988) : $unsigned((7'h4a)))));
            end
          reg2102 <= $unsigned((~&$signed($unsigned($unsigned(reg2091)))));
          if ($unsigned(($unsigned((~^reg1973)) ?
              $signed($unsigned($unsigned(reg2101))) : ($unsigned((reg2071 ?
                  reg2085 : reg2007)) ^~ $signed((reg2088 ?
                  reg1994 : reg2088))))))
            begin
              reg2103 = reg2042;
              reg2104 <= (~&(($signed((reg2070 >= reg2097)) ?
                  $signed($signed(reg2092)) : $signed((reg2059 ?
                      reg2098 : reg2014))) + $unsigned($signed($signed(reg2078)))));
              reg2105 <= (^reg2072[(5'h1d):(5'h1b)]);
              reg2106 <= {(((~&reg2101[(4'h8):(2'h3)]) + $signed((-reg1981))) - (reg2003 ~^ reg2099)),
                  (-$signed(reg2098)),
                  $signed({$unsigned($unsigned(reg2029)),
                      $signed($signed(reg2061)),
                      $unsigned((+reg2045))})};
              reg2107 <= {$signed(reg2103),
                  $signed(reg1988),
                  {$signed(reg2035),
                      $signed((+(reg2085 ? reg2078 : reg1978))),
                      (&((~&reg2073) ? (^~reg2099) : $signed(reg2085)))}};
              reg2108 = reg2103[(5'h17):(1'h1)];
              reg2109 <= (($unsigned(reg2098) > {{(8'hb3),
                      (forvar2090 - reg2094),
                      (7'h43)}}) >> $signed((|($signed(reg2032) ?
                  (reg2089 ? reg2077 : reg2056) : (&reg1973)))));
            end
          else
            begin
              reg2103 = ({$unsigned(({wire1965, (7'h56)} ?
                          $signed(reg2085) : $signed(reg2082))),
                      reg2089} ?
                  ($signed((8'hb6)) ^~ reg2003) : wire1962);
              reg2104 <= ((reg1999[(4'h9):(3'h4)] & $signed(($unsigned(reg1988) << (^~(8'ha5))))) << (~&$unsigned(reg1973[(5'h19):(5'h14)])));
            end
          reg2110 <= (~|reg2062[(5'h11):(4'hd)]);
        end
    end
  always
    @(posedge clk) begin
      reg2111 = reg1994;
      reg2112 <= (reg2070[(5'h1d):(5'h18)] ?
          reg2036 : ($signed((~^$signed(wire1962))) ?
              {$unsigned({reg1995, reg2078, reg2045}), reg2105} : (!reg2018)));
    end
  always
    @(posedge clk) begin
      reg2113 <= {(8'hb8), {reg2059}};
      for (forvar2114 = (1'h0); (forvar2114 < (2'h2)); forvar2114 = (forvar2114 + (1'h1)))
        begin
          if ((|reg2109[(2'h3):(1'h0)]))
            begin
              reg2115 <= (reg2056[(3'h6):(3'h4)] >>> (7'h52));
              reg2116 = $signed(reg2092[(4'hc):(1'h1)]);
            end
          else
            begin
              reg2115 <= reg1999;
              reg2117 <= (7'h40);
            end
          if ($unsigned((reg2071 >= {(((8'hba) - reg1973) && (~&reg1994)),
              $unsigned(reg2039[(2'h3):(2'h3)])})))
            begin
              reg2118 = reg1973;
              reg2119 <= ($unsigned($unsigned(reg2056)) ?
                  (^(reg2118 | {{reg2106,
                          (8'haa),
                          reg2106}})) : (~^$signed((reg2059[(3'h6):(2'h3)] ?
                      reg2117[(2'h2):(2'h2)] : {reg2042, reg1999, (7'h57)}))));
              reg2120 <= $unsigned($unsigned((^reg1994[(5'h14):(4'hf)])));
              reg2121 <= ({$signed(reg2106),
                      $signed(((+reg2105) ~^ $unsigned(reg2061))),
                      $signed((7'h56))} ?
                  reg1970 : $signed({$unsigned((forvar2114 | reg2071)),
                      (!(&reg2066))}));
              reg2122 = (+reg2109);
            end
          else
            begin
              reg2118 = reg2021[(3'h6):(1'h0)];
              reg2119 <= {$signed(((!reg2070[(3'h6):(1'h1)]) != $unsigned((^~reg1998)))),
                  $unsigned(reg2063)};
              reg2120 <= (({reg2120,
                      ($signed(reg2035) ?
                          (reg1999 + reg2120) : $signed((8'ha6))),
                      ({reg2058} > reg2029[(3'h4):(1'h0)])} ?
                  $unsigned(reg2070[(1'h0):(1'h0)]) : $unsigned(reg2040)) | ($unsigned({(reg2088 ?
                      reg2071 : reg2105),
                  $unsigned(reg2042),
                  $signed(reg1985)}) > $unsigned({$signed(reg2041),
                  (reg2063 ~^ reg2040)})));
              reg2121 <= reg2062[(5'h13):(3'h7)];
              reg2123 <= (~&$signed((^~$unsigned((reg1981 <= reg2119)))));
            end
          reg2124 = (reg1971[(4'h9):(2'h3)] ?
              reg1976[(5'h19):(3'h5)] : (reg2014[(5'h12):(5'h11)] ?
                  reg2040[(1'h1):(1'h0)] : (!(((8'ha0) ^~ reg2073) * $signed(reg1998)))));
          reg2125 <= (reg2091[(3'h5):(3'h4)] ?
              (~|reg2121) : ($signed($signed((reg1988 << wire1964))) <= (&(reg2016[(3'h5):(1'h1)] >= (^~reg2061)))));
        end
      reg2126 <= $signed(reg2066[(4'h8):(2'h2)]);
      for (forvar2127 = (1'h0); (forvar2127 < (2'h2)); forvar2127 = (forvar2127 + (1'h1)))
        begin
          if (reg2010)
            begin
              reg2128 <= (&$signed(((8'hb6) ?
                  (reg2042[(3'h7):(3'h5)] >>> $signed(reg2018)) : {((7'h44) ?
                          (8'haa) : reg2081),
                      reg1970})));
            end
          else
            begin
              reg2128 <= reg1976;
              reg2129 <= $unsigned({$signed($signed(reg2115[(4'hc):(3'h6)])),
                  $unsigned((^(~^reg2014)))});
              reg2130 <= ((|reg2063[(3'h5):(1'h0)]) * {forvar2127[(5'h15):(3'h4)],
                  reg2010[(5'h16):(4'hf)],
                  (((!(8'haf)) ? reg1970 : reg2078) | $signed((~^reg2062)))});
              reg2131 <= $signed($signed(reg2088[(3'h5):(3'h5)]));
              reg2132 <= reg2107;
              reg2133 <= (reg2116 == $signed(((~&(+reg2063)) && $unsigned((reg2123 >= reg2016)))));
            end
          for (forvar2134 = (1'h0); (forvar2134 < (3'h5)); forvar2134 = (forvar2134 + (1'h1)))
            begin
              reg2135 = ($signed(reg2059[(1'h1):(1'h0)]) << {$unsigned((+reg2109))});
              reg2136 <= ({$unsigned((!$unsigned((7'h55)))),
                  $signed(reg1994[(5'h18):(4'ha)])} ^ (wire1964 ?
                  $signed((~&(reg2112 << reg2050))) : ($signed({reg2124}) ?
                      (7'h45) : $signed(reg2050))));
              reg2137 <= (reg2074 ?
                  $signed($signed({reg2029,
                      reg1989})) : reg1976[(4'hf):(4'h8)]);
              reg2138 = reg2061[(3'h4):(3'h4)];
              reg2139 <= $signed($unsigned($unsigned(($signed(reg2014) ?
                  $unsigned(reg2035) : reg1971[(5'h18):(5'h11)]))));
              reg2140 = (~^((!{(reg2120 ? wire1965 : (8'h9f)),
                      (reg1981 ? (7'h4d) : reg1978)}) ?
                  reg2106[(4'hd):(4'h9)] : ($unsigned(((8'h9d) ?
                          reg2039 : reg2135)) ?
                      $signed($unsigned(reg2098)) : $unsigned(reg1994[(5'h1b):(3'h7)]))));
            end
        end
      if (reg2056[(5'h14):(4'hc)])
        begin
          reg2141 <= $signed(wire1963[(4'he):(1'h1)]);
          reg2142 <= ((!reg2061) && $unsigned($signed((~{(8'h9e), reg2091}))));
          for (forvar2143 = (1'h0); (forvar2143 < (3'h4)); forvar2143 = (forvar2143 + (1'h1)))
            begin
              reg2144 <= (~(~&((~&reg2118) ?
                  reg2011[(1'h1):(1'h1)] : (~&(reg1996 ? reg2133 : reg2061)))));
              reg2145 <= reg2141;
            end
          reg2146 <= ({$unsigned(((~&reg2121) ? reg2107 : reg2116)),
              {reg2010},
              reg2081} != reg2035[(2'h3):(1'h1)]);
          if ($signed($unsigned((forvar2114[(4'hf):(2'h2)] ?
              $unsigned($unsigned(reg2139)) : $signed($unsigned(reg2144))))))
            begin
              reg2147 = reg2055[(1'h1):(1'h0)];
              reg2148 = $signed($signed($unsigned((reg2071 ?
                  {reg2133, reg2078, reg2031} : (reg1999 ?
                      reg1969 : reg2055)))));
              reg2149 = $unsigned({reg2131});
              reg2150 <= $signed($unsigned(reg2034[(5'h18):(5'h11)]));
            end
          else
            begin
              reg2150 <= reg2102[(3'h5):(1'h0)];
            end
          reg2151 <= (&$signed($unsigned((-(reg2021 ? reg2137 : reg2002)))));
        end
      else
        begin
          for (forvar2141 = (1'h0); (forvar2141 < (2'h2)); forvar2141 = (forvar2141 + (1'h1)))
            begin
              reg2142 <= ($signed(reg1973[(5'h19):(4'hf)]) ?
                  (reg2092 ?
                      ((8'hab) ?
                          (~$signed((7'h48))) : ($unsigned((7'h50)) ?
                              ((7'h56) ?
                                  reg2055 : reg2129) : reg2132[(3'h6):(2'h3)])) : (^~{$unsigned(reg2123),
                          reg2027[(2'h2):(1'h0)]})) : ((~^($unsigned((8'haa)) ?
                      $signed(reg1978) : (reg2036 ?
                          reg1981 : reg2003))) << ($unsigned((reg1979 ?
                          reg1979 : reg2040)) ?
                      {$signed(reg2132)} : $unsigned($unsigned(reg2119)))));
              reg2143 <= forvar2127[(5'h19):(3'h6)];
              reg2144 <= reg1979[(4'he):(1'h1)];
            end
          if (reg2035[(2'h2):(2'h2)])
            begin
              reg2147 = ((&$signed((^~$unsigned(reg2070)))) <<< $signed(reg2018[(4'h8):(2'h2)]));
              reg2150 <= reg2059[(1'h0):(1'h0)];
              reg2152 = {reg2032, forvar2134};
              reg2153 <= (reg2145 ?
                  {(-(^(8'ha8))),
                      reg2112[(5'h19):(1'h0)]} : ($unsigned($signed((reg2131 != reg2007))) <= (({reg2122,
                              reg2097,
                              reg2123} ?
                          (8'ha1) : $unsigned(reg2144)) ?
                      ({(7'h4d), reg2058} ?
                          (^~reg2106) : $signed(reg2050)) : (reg2125 ?
                          reg2148[(1'h1):(1'h0)] : reg2035[(3'h4):(2'h3)]))));
              reg2154 = $signed({$signed(reg2062), reg1979});
              reg2155 <= (+$unsigned(($unsigned(reg1989[(3'h4):(3'h4)]) ?
                  $unsigned(((7'h4e) >> reg2136)) : (-$unsigned(reg1981)))));
            end
          else
            begin
              reg2145 <= reg2107;
              reg2146 <= ($unsigned((&({(7'h50), reg2081, reg2091} ?
                  reg2113 : (reg2138 * reg2055)))) <<< reg2133[(1'h0):(1'h0)]);
              reg2150 <= (&((((7'h57) < $unsigned(reg2002)) <<< (&(reg2106 ?
                      reg2022 : reg2010))) ?
                  $unsigned($unsigned($unsigned(reg2061))) : ((~^(reg2021 & reg2079)) + (8'h9d))));
              reg2151 <= $unsigned((!((~^reg2113) ?
                  (reg2131 >>> (&reg2027)) : $signed((reg2074 || reg2052)))));
              reg2153 <= $signed(reg2011[(3'h6):(1'h0)]);
              reg2154 = (+(8'ha6));
              reg2156 = $signed((7'h41));
            end
          reg2157 <= $unsigned((8'ha2));
        end
      if ({($unsigned($signed((-reg2092))) * $signed($unsigned(reg2104))),
          $unsigned(reg2116)})
        begin
          reg2158 = (reg2056 || $unsigned($unsigned($unsigned((reg2074 ?
              reg2039 : reg2052)))));
          reg2159 <= (~&$signed($unsigned(((forvar2127 <<< reg2125) ?
              {reg2140, (7'h4e)} : (reg2063 ? reg2061 : reg2125)))));
          reg2160 <= (($signed($unsigned((^~reg2131))) - reg2063[(3'h5):(1'h1)]) ?
              (($unsigned(reg2016) ~^ reg2028) ?
                  (reg2041[(1'h1):(1'h0)] ?
                      reg1985 : ((reg2151 < reg2129) ?
                          reg2148 : reg2154[(4'h9):(4'h8)])) : reg2143) : ((((reg2131 ?
                      reg1971 : (7'h44)) & $signed(reg2156)) <= $signed(reg2159)) ?
                  (8'hb6) : (reg2014[(5'h17):(4'ha)] ?
                      (!{reg1976}) : ((reg2027 >> (7'h41)) ?
                          (reg2092 >>> wire1964) : $signed(reg2109)))));
          if ($signed(reg2036))
            begin
              reg2161 = (~&$signed(wire1964));
              reg2162 = (^~reg2137[(5'h12):(4'hb)]);
              reg2163 = ($signed(reg2136) ?
                  reg2157[(1'h1):(1'h0)] : (~&$unsigned(($signed(reg2073) ?
                      $signed(reg2156) : $unsigned(reg2045)))));
              reg2164 <= $signed(reg2147[(1'h1):(1'h0)]);
              reg2165 = $unsigned($unsigned({((-forvar2134) < reg2131),
                  (7'h47),
                  (!wire1965[(5'h18):(5'h14)])}));
            end
          else
            begin
              reg2161 = $signed({$signed(((reg2011 ?
                      forvar2143 : (7'h4a)) <= (~&reg2158))),
                  ({$signed((8'h9d))} || {$signed((8'had))}),
                  {$signed((reg2022 != reg2078)),
                      (|reg2083),
                      (reg2074 ^ (~^forvar2143))}});
              reg2162 = (&reg2040);
              reg2164 <= $unsigned(reg2050[(5'h10):(1'h0)]);
              reg2165 = $signed((-(reg2157[(2'h3):(2'h2)] ?
                  $unsigned((^~(7'h4c))) : reg2016)));
              reg2166 = $unsigned({$signed(reg2144[(4'h9):(1'h1)]),
                  reg1971[(5'h10):(5'h10)]});
            end
          reg2167 = {reg2098[(4'h9):(2'h3)]};
        end
      else
        begin
          for (forvar2158 = (1'h0); (forvar2158 < (3'h5)); forvar2158 = (forvar2158 + (1'h1)))
            begin
              reg2159 <= $unsigned(reg2027);
            end
          reg2161 = {$signed({(+$signed(reg2053)),
                  $unsigned((+(8'hb0))),
                  $unsigned((~&reg2061))}),
              (($signed(((7'h51) <<< reg1980)) > ($unsigned((7'h4d)) ?
                  reg2036 : $unsigned(forvar2134))) << $unsigned($unsigned(reg2061))),
              {reg2107, reg1988[(1'h1):(1'h0)]}};
        end
      for (forvar2168 = (1'h0); (forvar2168 < (3'h6)); forvar2168 = (forvar2168 + (1'h1)))
        begin
          reg2169 <= $signed({reg2142});
          if (($signed((($unsigned(reg2160) ? (reg2091 < (7'h51)) : reg2031) ?
              reg1996[(4'ha):(2'h2)] : $unsigned(reg2014))) & ((&$unsigned(reg2003[(1'h0):(1'h0)])) ?
              $unsigned((!reg2118[(5'h11):(2'h3)])) : ($signed($unsigned(reg2143)) ?
                  ($signed(reg2137) != {reg2128,
                      reg2070,
                      reg1996}) : (+(reg2145 ? reg2056 : reg2148))))))
            begin
              reg2170 = ((7'h4a) + ($unsigned($unsigned((reg2034 >> reg1978))) ?
                  $signed({forvar2141,
                      (reg2139 >> (8'ha8))}) : $unsigned($unsigned($unsigned(reg2122)))));
              reg2171 <= (^~$unsigned($unsigned(reg2055)));
            end
          else
            begin
              reg2171 <= $unsigned((~^$signed($signed(reg2063))));
            end
          if (wire1964[(3'h4):(1'h1)])
            begin
              reg2172 = $signed($unsigned(($unsigned((reg2083 ?
                      reg2045 : reg2014)) ?
                  ((reg2119 ? reg2150 : (8'ha1)) & reg2079) : {reg1985,
                      reg2144,
                      (forvar2141 - reg1982)})));
              reg2173 <= (&(~|wire1963[(5'h15):(2'h3)]));
              reg2174 = (|(|(((^~(7'h50)) == $unsigned(reg2058)) && ($unsigned(reg2031) ?
                  $unsigned(forvar2134) : reg1995))));
              reg2175 = $signed($signed($signed(wire1962[(3'h7):(2'h3)])));
              reg2176 = $unsigned((&reg2133));
              reg2177 <= $unsigned(((|(reg1989[(3'h7):(3'h5)] || (-(8'hb9)))) ?
                  (($signed(reg2174) >= {reg2040,
                      reg2116}) ~^ {$unsigned(reg2139),
                      (reg2078 ? reg2027 : forvar2141),
                      $signed(reg2091)}) : {{(+reg2118),
                          reg2151[(4'hb):(1'h0)]},
                      {$signed(reg2149), reg2066}}));
            end
          else
            begin
              reg2172 = ((-($unsigned(reg2021[(1'h1):(1'h0)]) ?
                  reg2056[(5'h1b):(5'h12)] : ((reg2121 || reg2053) ^~ reg2098))) <= (~reg2113[(2'h2):(2'h2)]));
              reg2173 <= $signed((~((+((8'ha0) ?
                  reg2173 : reg2153)) + {(~|reg2088), reg2088})));
              reg2174 = {reg2105};
              reg2175 = {((~|(forvar2127 >> $signed(reg1998))) << ((~&reg2170) ?
                      (^reg1988) : $signed($signed((8'ha1))))),
                  reg2133[(2'h3):(2'h2)]};
            end
          for (forvar2178 = (1'h0); (forvar2178 < (1'h1)); forvar2178 = (forvar2178 + (1'h1)))
            begin
              reg2179 = (8'ha4);
              reg2180 <= (reg2083[(1'h1):(1'h0)] ?
                  reg2029 : $unsigned($unsigned(reg1985[(5'h15):(4'he)])));
            end
          if (reg2135[(4'hd):(4'h8)])
            begin
              reg2181 = reg2162[(1'h1):(1'h1)];
              reg2182 <= $signed(reg2029);
              reg2183 = {reg2130[(2'h3):(2'h3)],
                  ((|(7'h4b)) + (-$unsigned(reg2126[(2'h3):(1'h0)])))};
            end
          else
            begin
              reg2182 <= (~|$unsigned((({reg2150} ?
                      reg2112[(4'he):(4'hc)] : (reg2126 & reg2097)) ?
                  reg2031[(1'h0):(1'h0)] : ($unsigned(reg2028) ?
                      (reg1981 ? reg2133 : reg1996) : reg2119))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg2184 = $signed(((+($signed(wire1966) < (-reg2027))) ^ $unsigned((^~(reg2110 ?
          (8'hb2) : reg2042)))));
      reg2185 <= $signed($signed($unsigned(((reg2011 ^~ reg1985) * $signed(reg2171)))));
      if ($unsigned($unsigned((^~(~|{reg2142, (7'h4e)})))))
        begin
          reg2186 = $signed(reg2123);
          for (forvar2187 = (1'h0); (forvar2187 < (2'h3)); forvar2187 = (forvar2187 + (1'h1)))
            begin
              reg2188 = reg2182;
            end
        end
      else
        begin
          reg2187 <= (!reg2011);
          if (((reg2083[(2'h3):(2'h3)] - $signed((reg2153 ?
                  reg2055 : (reg2066 ? reg2129 : forvar2187)))) ?
              $unsigned(($unsigned((reg2039 ^~ (8'hbc))) ?
                  (reg2106[(3'h4):(1'h1)] ^~ (wire1964 ?
                      reg2018 : (7'h4e))) : ((reg2169 != reg2061) >= (reg1998 ?
                      reg2112 : reg2106)))) : $signed($unsigned($signed({reg2169,
                  reg2073,
                  reg2137})))))
            begin
              reg2188 = $signed(($unsigned($unsigned(reg2091[(4'h8):(1'h0)])) >= (~|$signed({reg2117}))));
            end
          else
            begin
              reg2189 <= $signed((($signed(reg2133[(2'h3):(1'h1)]) | $signed((~|reg2039))) ^ $signed({$unsigned((7'h47)),
                  $signed(wire1966),
                  $signed(reg2155)})));
            end
          for (forvar2190 = (1'h0); (forvar2190 < (1'h1)); forvar2190 = (forvar2190 + (1'h1)))
            begin
              reg2191 = (~(~$signed(reg2029)));
              reg2192 = reg1971;
              reg2193 = $unsigned(reg2040[(3'h7):(1'h1)]);
            end
          reg2194 <= $unsigned(reg1994[(3'h6):(3'h4)]);
          reg2195 = (^$unsigned((8'hbd)));
          reg2196 = (-reg2066[(3'h7):(1'h1)]);
        end
      reg2197 = $unsigned($signed(reg2196[(5'h18):(4'hb)]));
      for (forvar2198 = (1'h0); (forvar2198 < (1'h1)); forvar2198 = (forvar2198 + (1'h1)))
        begin
          for (forvar2199 = (1'h0); (forvar2199 < (3'h6)); forvar2199 = (forvar2199 + (1'h1)))
            begin
              reg2200 <= $signed($signed(($unsigned((reg2153 && reg2120)) ?
                  $signed((7'h4a)) : $signed((+(7'h49))))));
              reg2201 = reg1996;
              reg2202 <= $unsigned((reg2022 <<< ($signed((~|reg2125)) ?
                  (reg2003[(2'h2):(1'h0)] << reg2059) : reg2137)));
              reg2203 = reg2035;
              reg2204 = reg2112;
            end
          for (forvar2205 = (1'h0); (forvar2205 < (3'h4)); forvar2205 = (forvar2205 + (1'h1)))
            begin
              reg2206 <= $unsigned(({(~{(7'h4a)}),
                  (reg2169 >>> (~|(8'ha5))),
                  {$unsigned(reg2151)}} ~^ $unsigned((^(reg2002 ?
                  reg2061 : wire1965)))));
              reg2207 = $unsigned((reg2110 ? reg2059 : $signed((|reg2171))));
            end
          reg2208 <= reg2119;
        end
    end
  assign wire2209 = $signed($unsigned((~|((reg2055 ^ reg2125) ?
                        (reg2107 == reg2018) : reg2035[(2'h3):(2'h2)]))));
  assign wire2210 = ((((^~reg2052[(3'h7):(3'h7)]) > $unsigned({reg2206,
                            reg2145,
                            reg1969})) ?
                        $unsigned((&(reg2208 ~^ reg2145))) : $unsigned(reg2115)) >>> {{($unsigned(reg2028) ?
                                reg2141[(3'h5):(2'h2)] : (-reg2177)),
                            reg1981}});
  assign wire2211 = $unsigned(((~^$signed(reg2132)) << ($unsigned((reg2109 ?
                            (8'hac) : reg1995)) ?
                        $unsigned({reg2155, reg2022}) : $unsigned((8'hb5)))));
  assign wire2212 = $unsigned(({$unsigned({reg1976}),
                        $unsigned(reg2041[(5'h1a):(5'h15)])} >>> ((^~(^~reg2208)) ^~ (+(reg2119 + reg2081)))));
  assign wire2213 = (wire1967 <= (~^$signed($signed($unsigned(reg2132)))));
  always
    @(posedge clk) begin
      for (forvar2214 = (1'h0); (forvar2214 < (3'h6)); forvar2214 = (forvar2214 + (1'h1)))
        begin
          reg2215 <= (reg2177[(5'h14):(4'hb)] ?
              ($signed((8'ha7)) <= $unsigned($unsigned((+reg2031)))) : $unsigned($signed(reg2056)));
          reg2216 = $unsigned(((wire1967[(4'h9):(3'h7)] ^~ ($unsigned(wire1965) ?
                  ((8'ha7) ? reg2208 : reg2059) : (reg2056 == wire1966))) ?
              (~reg2110) : ($signed((reg2189 ?
                  reg1982 : reg2137)) <= (!$signed(reg2117)))));
          for (forvar2217 = (1'h0); (forvar2217 < (3'h4)); forvar2217 = (forvar2217 + (1'h1)))
            begin
              reg2218 = reg2109[(2'h2):(1'h1)];
              reg2219 <= reg2121[(2'h2):(1'h0)];
              reg2220 = (~(reg2022 ?
                  $signed(reg2173[(4'hb):(2'h2)]) : ($signed((~|wire2211)) | (^~$signed(reg2151)))));
              reg2221 <= reg2078;
              reg2222 = $unsigned($unsigned($unsigned({$unsigned(reg1985)})));
              reg2223 = $signed((~(reg2061 ? (~reg2105) : reg2022)));
              reg2224 = (!$signed((reg2053[(1'h1):(1'h1)] || reg2061)));
            end
          reg2225 <= {reg2121, reg2041};
          for (forvar2226 = (1'h0); (forvar2226 < (1'h0)); forvar2226 = (forvar2226 + (1'h1)))
            begin
              reg2227 = (+(|reg1985[(4'ha):(3'h6)]));
              reg2228 = {({((reg2002 ? reg2117 : reg2053) >= reg2225),
                      reg2218[(4'hc):(3'h7)]} >>> $unsigned(($signed(reg2126) ?
                      reg2146 : reg2097))),
                  ((8'hb5) < {($signed(reg1973) != reg2131),
                      (^~$signed((8'ha1))),
                      $unsigned($signed(reg2007))}),
                  forvar2214};
              reg2229 = ($signed($signed({(reg2007 ? reg2169 : (7'h4a))})) ?
                  ($signed(reg2003) ?
                      reg2177[(3'h6):(3'h5)] : (~|reg2202)) : (7'h41));
            end
        end
      reg2230 <= ($unsigned((^~(+(~|reg1979)))) ?
          $unsigned($signed($unsigned($unsigned(reg2180)))) : (~{(^~(reg2224 | (8'hb6)))}));
      for (forvar2231 = (1'h0); (forvar2231 < (3'h4)); forvar2231 = (forvar2231 + (1'h1)))
        begin
          for (forvar2232 = (1'h0); (forvar2232 < (1'h1)); forvar2232 = (forvar2232 + (1'h1)))
            begin
              reg2233 = ($signed((((wire2211 ? reg2053 : reg2063) ^ (wire1966 ?
                          wire1962 : wire2210)) ?
                      reg2073 : (&{reg2220, wire1962}))) ?
                  $signed((wire2213 ?
                      $unsigned($signed(reg2045)) : ((reg2117 + reg2189) ?
                          $signed(reg2136) : $signed(reg2137)))) : (reg2137[(4'hc):(4'hb)] ?
                      ((reg2123 << (8'h9d)) ?
                          {reg2106[(2'h2):(1'h0)],
                              (reg2131 ?
                                  reg1998 : reg2218)} : $signed(reg2132[(1'h0):(1'h0)])) : $signed(($unsigned(reg2007) >>> (8'hbd)))));
            end
          for (forvar2234 = (1'h0); (forvar2234 < (2'h3)); forvar2234 = (forvar2234 + (1'h1)))
            begin
              reg2235 = (($signed($signed(((8'hb7) || reg2110))) ?
                      (reg2157 <<< $signed($unsigned(reg2208))) : reg1971[(4'hb):(4'hb)]) ?
                  (reg2130 ?
                      $unsigned(((reg2200 * (8'h9f)) ?
                          reg2202 : $signed(reg2027))) : {(~|(reg2128 ?
                              reg2157 : reg2042)),
                          (7'h46)}) : reg2187[(3'h7):(3'h5)]);
              reg2236 = (~|(reg2202[(4'ha):(3'h7)] ?
                  $signed(reg2150) : $unsigned(reg2029)));
            end
          reg2237 = reg2180;
        end
      reg2238 <= $unsigned(reg1981[(5'h1b):(1'h1)]);
      if ((reg2151[(4'h9):(1'h1)] ? (^(-reg2227)) : forvar2217))
        begin
          reg2239 <= reg2173;
          for (forvar2240 = (1'h0); (forvar2240 < (3'h4)); forvar2240 = (forvar2240 + (1'h1)))
            begin
              reg2241 = ($signed((({reg2151,
                  reg2173,
                  reg2224} * reg2219[(3'h6):(3'h6)]) <<< ((reg2078 | reg2092) ?
                  (reg2115 - reg2180) : (-reg2120)))) || reg2113[(2'h3):(1'h0)]);
              reg2242 = $signed({(!$signed($unsigned(reg2235)))});
              reg2243 = {reg2225[(4'hd):(3'h5)],
                  $signed($signed((-$signed(reg1994)))),
                  (~&$unsigned(($signed((8'hbb)) || reg2018[(1'h1):(1'h0)])))};
              reg2244 = ($signed($unsigned((~$unsigned(reg2010)))) - reg2141[(5'h15):(4'he)]);
            end
          reg2245 = reg2036[(3'h4):(1'h1)];
          reg2246 = $unsigned((&{{{reg2121, reg2052}}}));
          reg2247 <= (reg2014[(5'h17):(5'h12)] ?
              reg2125[(4'hb):(4'h9)] : (8'ha8));
          reg2248 = (reg1989[(3'h6):(1'h0)] << $signed((-$unsigned(reg1998))));
          reg2249 <= ({(~|((~reg2238) ?
                      ((7'h41) ? reg2002 : reg2115) : (+reg2224)))} ?
              (reg1981 ?
                  ((reg1985 | $unsigned(reg2062)) ?
                      $signed(reg2224[(5'h19):(5'h14)]) : (&(reg2107 + reg2247))) : $signed($unsigned($unsigned(reg2206)))) : reg2014[(5'h18):(1'h0)]);
        end
      else
        begin
          reg2240 = $signed(((&$unsigned($unsigned(reg2219))) >> (wire2210[(2'h2):(2'h2)] ?
              reg2246[(4'he):(4'h8)] : ($signed(reg2189) > reg2102))));
          for (forvar2241 = (1'h0); (forvar2241 < (3'h4)); forvar2241 = (forvar2241 + (1'h1)))
            begin
              reg2247 <= $signed((^reg1979));
            end
          reg2249 <= ($unsigned($unsigned($unsigned($signed(reg2078)))) & ($signed(reg2056) > ($unsigned({(8'hbf)}) | $signed($unsigned(reg2177)))));
          reg2250 <= (^~($signed($unsigned(reg2074)) ?
              {$unsigned(reg2230), (~(^~(7'h45)))} : reg1976[(5'h10):(1'h0)]));
          if ({((forvar2214[(2'h3):(1'h1)] ^~ reg2141[(2'h2):(1'h0)]) ?
                  $unsigned($unsigned(reg2123[(4'he):(3'h4)])) : reg1969[(5'h11):(4'h9)]),
              ($signed(($signed(reg2092) <= $signed(reg2132))) ?
                  $signed(reg2041[(5'h1b):(1'h0)]) : ($unsigned($signed(reg2200)) ?
                      reg2032[(3'h7):(3'h5)] : reg2031))})
            begin
              reg2251 = (&({($signed((8'hbf)) ^ (reg1978 ?
                      (8'haf) : (8'hbe)))} != ($unsigned(forvar2241[(4'h8):(4'h8)]) < ($unsigned((7'h46)) > (reg2239 | forvar2231)))));
              reg2252 <= (wire2212[(3'h4):(1'h0)] ?
                  (reg2115 & ($unsigned(reg2045[(3'h5):(3'h4)]) ?
                      reg2224 : $signed($unsigned(reg2225)))) : reg1973[(5'h13):(4'hc)]);
              reg2253 <= reg2145[(4'he):(3'h4)];
              reg2254 = reg2142;
              reg2255 <= (^~((!(^~reg2246[(3'h6):(3'h5)])) ^~ reg2078));
            end
          else
            begin
              reg2251 = ((!forvar2226) != (|(~|$unsigned((+reg2243)))));
            end
          for (forvar2256 = (1'h0); (forvar2256 < (3'h5)); forvar2256 = (forvar2256 + (1'h1)))
            begin
              reg2257 <= reg2223[(5'h12):(5'h11)];
              reg2258 <= (reg2142 & $signed(((8'hb0) ?
                  reg2074[(4'hc):(2'h3)] : ($signed(reg2215) < reg1998[(4'ha):(4'h8)]))));
              reg2259 = reg2235;
              reg2260 <= {reg2222};
              reg2261 = (!reg2222[(4'hf):(2'h3)]);
              reg2262 <= (~$unsigned(reg1994));
            end
          reg2263 <= ((~|reg2259[(4'hd):(4'hb)]) <= {reg2153[(2'h2):(1'h1)]});
        end
    end
  always
    @(posedge clk) begin
      if ($signed($signed(reg2253)))
        begin
          reg2264 <= {(~|reg2003[(2'h2):(1'h0)]),
              {(+reg1973[(1'h1):(1'h1)]),
                  $unsigned((reg2031[(2'h3):(1'h1)] > (reg2145 ^~ reg2164)))},
              {$unsigned(reg1985),
                  ((|reg2079) ?
                      ($unsigned(reg2157) ?
                          reg2088[(4'he):(3'h5)] : reg2258[(1'h1):(1'h1)]) : ($signed(reg2257) ?
                          $signed(reg1999) : wire2212[(2'h2):(1'h0)])),
                  reg2081[(3'h4):(2'h2)]}};
          if ($unsigned((~&(!reg2144))))
            begin
              reg2265 = (((((~^reg2083) ?
                      $unsigned(reg2011) : reg2264) > (reg2202[(5'h12):(1'h1)] >= reg2250[(3'h5):(1'h1)])) ?
                  (reg2206[(5'h12):(1'h1)] >= (7'h4b)) : ($signed($unsigned(reg2042)) == $unsigned(((7'h4e) ?
                      wire1967 : reg2239)))) >>> reg2107);
              reg2266 = ((reg2031[(2'h3):(1'h0)] ?
                      (7'h43) : reg2230[(5'h1a):(4'hd)]) ?
                  ((((~^reg2153) ? {reg2252, reg2014} : $signed(reg2119)) ?
                      reg2219[(4'h9):(1'h1)] : wire1965) != ({(wire1967 | wire1962)} || reg2066[(3'h6):(3'h5)])) : (({$unsigned((7'h4c)),
                          $signed(reg2189)} ?
                      reg2169 : {(reg2128 ? (8'hbd) : reg2164),
                          reg2257[(4'hd):(4'hb)]}) ~^ reg2074[(5'h11):(5'h11)]));
              reg2267 <= $unsigned(reg2206[(5'h18):(5'h10)]);
            end
          else
            begin
              reg2267 <= $unsigned($signed((reg2249[(3'h4):(3'h4)] ?
                  reg2164[(3'h7):(1'h1)] : reg1988[(3'h7):(1'h0)])));
              reg2268 = (~|reg2117[(3'h4):(2'h2)]);
              reg2269 = (reg2252 ?
                  {{$signed(reg1969[(5'h18):(4'hd)]),
                          reg2070[(3'h5):(3'h5)],
                          $signed((reg2032 != reg2131))}} : (wire1962[(1'h0):(1'h0)] ?
                      wire2211 : (~|$signed(reg2185))));
              reg2270 <= {$signed($unsigned(reg2056[(4'h8):(3'h7)]))};
              reg2271 = $unsigned((wire2211[(2'h3):(1'h0)] * $unsigned($signed((reg2066 ?
                  reg1969 : reg2265)))));
              reg2272 = $signed((($unsigned(((8'hb4) || (8'hb4))) + ($unsigned(reg2269) ?
                      {reg2206} : (wire2213 ? (8'hb0) : (7'h4f)))) ?
                  (^(+{reg2144})) : {$signed((&reg2126))}));
            end
          for (forvar2273 = (1'h0); (forvar2273 < (3'h4)); forvar2273 = (forvar2273 + (1'h1)))
            begin
              reg2274 <= reg2070;
              reg2275 = ($unsigned($signed(reg1988)) ?
                  (reg2264[(4'hf):(3'h6)] ^ ((reg2265 > $unsigned((7'h53))) - reg2071)) : reg2056[(5'h13):(4'hd)]);
              reg2276 <= (reg2045[(5'h10):(3'h5)] <<< reg2185);
            end
          if ((^{$unsigned(({reg1985, (8'ha7), wire2211} != {reg1970,
                  reg2107,
                  reg2253})),
              reg2031[(1'h1):(1'h0)]}))
            begin
              reg2277 = (!{$unsigned(((&wire2210) ? reg2136 : (&reg2010))),
                  ((^~{reg2056, reg2113}) ?
                      {reg2052[(3'h5):(3'h5)]} : (~(reg2145 ?
                          reg2249 : wire1963)))});
              reg2278 = reg2056[(1'h1):(1'h1)];
            end
          else
            begin
              reg2277 = ((|$signed(reg2105)) >> (^(!{(reg1978 ?
                      reg2045 : reg2164)})));
              reg2278 = (-reg2268[(4'hb):(3'h5)]);
              reg2279 <= {({(~|reg2150), $signed(reg2265)} ?
                      (~$unsigned((reg2142 ?
                          reg2056 : (7'h43)))) : $unsigned($signed({reg2056,
                          reg1979}))),
                  $signed(wire1967[(4'hf):(3'h4)])};
              reg2280 <= (({reg1980[(4'hf):(4'hb)]} ?
                  (+reg2185) : reg2055[(3'h4):(2'h2)]) ^~ (reg1976 << (~^reg2187)));
              reg2281 = ($signed((~^(-(~&reg2081)))) ?
                  $signed($signed({(reg2059 ? wire1965 : reg2202),
                      wire2209})) : (7'h4f));
            end
        end
      else
        begin
          reg2264 <= (|((-{$signed(reg2260)}) ?
              ($signed($unsigned((8'hbf))) ?
                  reg2275[(1'h1):(1'h1)] : (~&(reg1969 || (8'haa)))) : (^{reg2050[(2'h3):(2'h2)]})));
          if ((reg2045 ?
              (($signed((reg2133 ?
                  reg2131 : (7'h50))) ^ (^~(&reg2052))) <<< forvar2273) : $signed((~|$signed(reg2221[(2'h3):(2'h2)])))))
            begin
              reg2267 <= (($unsigned(reg2022[(5'h17):(4'h8)]) >>> $unsigned(((reg2247 >> wire1962) ^ $signed((8'ha1))))) ?
                  $unsigned($signed((7'h40))) : $signed(reg2144[(4'ha):(2'h3)]));
              reg2268 = (~(~&((~^{reg2097, reg1976, reg2061}) ?
                  reg2136[(3'h7):(2'h2)] : $signed({(8'haa),
                      reg2258,
                      (7'h46)}))));
              reg2269 = reg2055[(1'h0):(1'h0)];
              reg2271 = (reg2250[(4'ha):(2'h2)] | (~|(~|reg2169)));
            end
          else
            begin
              reg2267 <= {reg2129, $signed($unsigned(reg2265[(5'h14):(4'hc)]))};
              reg2270 <= (~^$signed((8'hb4)));
              reg2271 = ($unsigned(($signed((8'ha9)) - $unsigned($unsigned(reg2032)))) * reg2050);
              reg2272 = $unsigned(((($signed(reg1995) && (reg2119 ?
                      reg2056 : (8'hac))) >> reg2263[(4'hd):(4'ha)]) ?
                  wire2213 : reg2121));
              reg2273 = $signed((~reg2271[(5'h16):(4'hb)]));
            end
          reg2275 = $unsigned($unsigned(((!(~&reg2271)) <<< reg2098[(4'hb):(3'h6)])));
          reg2276 <= (8'hbb);
        end
      reg2282 = $signed((($unsigned($unsigned(reg2081)) ?
          $signed(wire2213) : ((~^(8'ha9)) == $unsigned((7'h4c)))) > (((reg2281 ?
              reg2171 : reg2018) >= (reg2219 | reg2225)) ?
          ({reg2252,
              reg2115,
              reg2276} + reg2150[(4'hf):(4'hd)]) : reg2265[(5'h13):(1'h0)])));
    end
  always
    @(posedge clk) begin
      for (forvar2283 = (1'h0); (forvar2283 < (1'h0)); forvar2283 = (forvar2283 + (1'h1)))
        begin
          for (forvar2284 = (1'h0); (forvar2284 < (1'h0)); forvar2284 = (forvar2284 + (1'h1)))
            begin
              reg2285 = ($signed($unsigned((^reg2185))) && reg2088[(5'h16):(5'h16)]);
              reg2286 <= (~reg1985);
            end
          reg2287 = $signed(($signed(wire1965) << $unsigned(forvar2284[(2'h2):(1'h1)])));
          reg2288 <= reg2253;
          if ((~|$unsigned((($signed(reg1971) ? $signed((8'ha1)) : reg2219) ?
              (~reg1973[(4'hb):(3'h4)]) : ({reg2157,
                  (8'ha1),
                  reg2159} <<< (reg2062 & reg1998))))))
            begin
              reg2289 = {{(reg2036[(1'h0):(1'h0)] <<< $signed(reg2034)),
                      reg2045[(5'h10):(4'hd)],
                      (^$signed(wire1962))}};
            end
          else
            begin
              reg2290 <= reg2035;
              reg2291 <= (7'h46);
              reg2292 <= $unsigned((($unsigned((forvar2284 ?
                      reg1969 : wire1963)) >= $unsigned((reg2066 >> reg2200))) ?
                  (7'h4a) : ((&$signed(reg2133)) + $unsigned($signed(reg2092)))));
              reg2293 = (((reg2106 ?
                      $signed((-(8'hb6))) : (wire1963[(1'h1):(1'h0)] + reg2189)) * (&{(-reg2022),
                      reg2219[(4'h9):(3'h6)],
                      (^~reg2010)})) ?
                  {(|$signed(reg2119)),
                      ({{reg2208}} ?
                          ((reg2098 ?
                              (8'ha8) : reg2120) || (reg2061 >> reg2014)) : (reg2027[(3'h5):(2'h2)] ?
                              wire1964 : $signed(reg2262))),
                      $signed((wire1964 ?
                          reg2021 : reg2291[(3'h6):(3'h6)]))} : reg2073);
              reg2294 = ($unsigned((-(((8'hb5) << reg2078) + $unsigned(reg2010)))) >> $signed(((reg2062 != $signed(reg2066)) ?
                  reg2145[(5'h12):(4'hc)] : reg2142)));
            end
          reg2295 = reg2206;
        end
      for (forvar2296 = (1'h0); (forvar2296 < (3'h5)); forvar2296 = (forvar2296 + (1'h1)))
        begin
          reg2297 = $signed((^$signed($signed($signed(wire1967)))));
          for (forvar2298 = (1'h0); (forvar2298 < (2'h2)); forvar2298 = (forvar2298 + (1'h1)))
            begin
              reg2299 <= (reg2053[(5'h12):(3'h7)] && (~^reg2169));
              reg2300 = $signed(((wire2212[(1'h1):(1'h1)] ?
                  {$unsigned(reg2255),
                      reg2153[(1'h1):(1'h1)]} : ((reg2260 > reg2003) && (~|reg1976))) ~^ (^~$signed(reg2066))));
              reg2301 <= (reg2144 ?
                  (+{$signed(reg2032)}) : (reg2066[(4'hb):(1'h1)] ?
                      (((reg2039 ?
                          reg2123 : reg1969) != (+reg2276)) * (((8'hb2) < reg2299) ?
                          (reg2113 ?
                              reg2027 : reg2300) : $signed((7'h4b)))) : reg2238[(5'h10):(4'hc)]));
              reg2302 = reg2270;
            end
          if (reg2221)
            begin
              reg2303 <= $signed(reg2297[(4'hd):(2'h2)]);
              reg2304 <= (+$signed((({reg1980, reg2079} ?
                  (8'had) : ((7'h42) * reg2098)) & reg2297[(4'he):(4'hd)])));
              reg2305 <= (~|($signed(reg2091[(4'h9):(4'h8)]) == $unsigned(((reg2303 ?
                      reg2129 : reg2131) ?
                  (reg2136 >> reg2295) : (7'h41)))));
              reg2306 = $unsigned(reg2035);
            end
          else
            begin
              reg2303 <= reg1980[(2'h3):(1'h1)];
              reg2306 = (8'h9f);
              reg2307 <= ($unsigned((reg2230[(1'h0):(1'h0)] >>> (wire2212[(1'h1):(1'h1)] & $unsigned(reg2032)))) ?
                  reg1989 : reg2238[(5'h18):(3'h4)]);
              reg2308 = reg2189;
              reg2309 <= $signed($signed($unsigned((8'hbe))));
              reg2310 = reg2133;
            end
        end
      reg2311 <= reg2255;
      if ((8'had))
        begin
          if (reg2221[(1'h0):(1'h0)])
            begin
              reg2312 = ((&reg1981) ?
                  reg2189 : (reg2305[(4'he):(1'h0)] << reg2301[(1'h0):(1'h0)]));
              reg2313 = ($unsigned(reg2007) ? (~^reg2042) : $unsigned(reg1982));
              reg2314 <= (reg2219[(2'h2):(1'h1)] ?
                  reg2083[(3'h7):(1'h0)] : ($signed($signed(reg2088)) ?
                      reg2003[(2'h2):(1'h1)] : ($signed((^reg2303)) ?
                          {(reg2070 ? reg2257 : reg2249),
                              reg2070[(4'h8):(2'h2)]} : $unsigned((reg1982 ?
                              reg1982 : (8'hb6))))));
              reg2315 = (((((|reg2303) ?
                      (~|reg2120) : reg2286) > ($unsigned((8'ha8)) <= (reg2027 ?
                      wire1963 : (8'hbb)))) ?
                  ((|$unsigned(wire1966)) ?
                      reg1989 : {$unsigned((8'hac))}) : forvar2284[(1'h1):(1'h0)]) << $unsigned(reg1970));
              reg2316 <= $unsigned(reg2215[(1'h1):(1'h0)]);
              reg2317 <= (reg2091 ?
                  {(^$signed(reg2136[(3'h4):(2'h3)])),
                      ((reg2260 ? reg2153[(1'h1):(1'h1)] : reg1976) ~^ reg2104),
                      $unsigned($signed((reg2007 <= reg2267)))} : reg2262);
            end
          else
            begin
              reg2312 = $unsigned(reg2102);
              reg2314 <= $signed((($signed(reg2053[(5'h10):(4'h9)]) ?
                      reg2088[(4'hf):(4'he)] : $unsigned($signed((7'h52)))) ?
                  reg2098[(4'h8):(3'h4)] : $signed({reg1978})));
            end
          reg2318 <= $unsigned($unsigned((7'h50)));
        end
      else
        begin
          for (forvar2312 = (1'h0); (forvar2312 < (3'h5)); forvar2312 = (forvar2312 + (1'h1)))
            begin
              reg2313 = (~^{(!reg2185),
                  $unsigned((^~(reg2299 ? reg2293 : (8'hb5)))),
                  {reg2150}});
            end
        end
      reg2319 <= ($unsigned((reg2307 ?
              ((forvar2283 ?
                  reg2097 : reg2200) * ((8'ha5) > reg2239)) : reg2002[(2'h2):(1'h1)])) ?
          (($unsigned($unsigned(reg2062)) | ((reg2189 & reg2239) ?
                  reg2055[(3'h6):(3'h5)] : (reg2157 ? reg2305 : reg2106))) ?
              $unsigned(reg2126) : (($signed(wire2213) >> reg2253[(4'hd):(3'h4)]) ^ (|{reg1994,
                  (8'ha1),
                  (8'hae)}))) : reg2091[(4'ha):(4'h8)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1686  (y, clk, wire1691, wire1690, wire1689, wire1688, wire1687);
  output wire [(32'hde2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire1691;
  input wire [(5'h14):(1'h0)] wire1690;
  input wire [(5'h1d):(1'h0)] wire1689;
  input wire [(5'h1d):(1'h0)] wire1688;
  input wire signed [(4'hb):(1'h0)] wire1687;
  wire [(5'h1a):(1'h0)] wire1905;
  wire [(4'h9):(1'h0)] wire1833;
  wire signed [(4'hb):(1'h0)] wire1832;
  wire [(5'h1c):(1'h0)] wire1814;
  wire [(4'he):(1'h0)] wire1810;
  wire signed [(5'h1c):(1'h0)] wire1809;
  wire [(5'h13):(1'h0)] wire1693;
  wire signed [(4'hb):(1'h0)] wire1692;
  reg [(3'h7):(1'h0)] reg1903 = (1'h0);
  reg [(3'h5):(1'h0)] reg1902 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1900 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1892 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1890 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1888 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1887 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1885 = (1'h0);
  reg [(4'hb):(1'h0)] reg1884 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1880 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1879 = (1'h0);
  reg [(5'h12):(1'h0)] reg1874 = (1'h0);
  reg [(4'ha):(1'h0)] reg1873 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1869 = (1'h0);
  reg [(5'h11):(1'h0)] reg1862 = (1'h0);
  reg [(5'h17):(1'h0)] reg1861 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1857 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1856 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1855 = (1'h0);
  reg [(4'h8):(1'h0)] reg1834 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1852 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1850 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1846 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1843 = (1'h0);
  reg [(2'h3):(1'h0)] reg1842 = (1'h0);
  reg [(5'h19):(1'h0)] reg1835 = (1'h0);
  reg [(5'h17):(1'h0)] reg1831 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1829 = (1'h0);
  reg [(4'hd):(1'h0)] reg1828 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1827 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1826 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1825 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1820 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1819 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1818 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1817 = (1'h0);
  reg [(3'h6):(1'h0)] reg1812 = (1'h0);
  reg [(5'h16):(1'h0)] reg1811 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1808 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1804 = (1'h0);
  reg [(4'hc):(1'h0)] reg1803 = (1'h0);
  reg [(3'h4):(1'h0)] reg1799 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1795 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1794 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1791 = (1'h0);
  reg [(4'hb):(1'h0)] reg1786 = (1'h0);
  reg [(5'h12):(1'h0)] reg1785 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1784 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1782 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1781 = (1'h0);
  reg [(4'h8):(1'h0)] reg1780 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1778 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1776 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1774 = (1'h0);
  reg [(5'h12):(1'h0)] reg1773 = (1'h0);
  reg [(3'h5):(1'h0)] reg1768 = (1'h0);
  reg [(3'h5):(1'h0)] reg1766 = (1'h0);
  reg [(3'h4):(1'h0)] reg1765 = (1'h0);
  reg [(4'hb):(1'h0)] reg1764 = (1'h0);
  reg [(5'h16):(1'h0)] reg1762 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1761 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1756 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1753 = (1'h0);
  reg [(4'hb):(1'h0)] reg1750 = (1'h0);
  reg [(5'h14):(1'h0)] reg1748 = (1'h0);
  reg [(3'h7):(1'h0)] reg1747 = (1'h0);
  reg [(5'h16):(1'h0)] reg1746 = (1'h0);
  reg [(3'h4):(1'h0)] reg1744 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1743 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1739 = (1'h0);
  reg [(3'h6):(1'h0)] reg1738 = (1'h0);
  reg [(5'h14):(1'h0)] reg1736 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1735 = (1'h0);
  reg [(2'h2):(1'h0)] reg1734 = (1'h0);
  reg [(5'h11):(1'h0)] reg1732 = (1'h0);
  reg [(5'h15):(1'h0)] reg1730 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1728 = (1'h0);
  reg [(4'hb):(1'h0)] reg1719 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1716 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1714 = (1'h0);
  reg [(5'h18):(1'h0)] reg1711 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1710 = (1'h0);
  reg [(5'h13):(1'h0)] reg1707 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1706 = (1'h0);
  reg [(4'hb):(1'h0)] reg1705 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1704 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1703 = (1'h0);
  reg [(5'h17):(1'h0)] reg1702 = (1'h0);
  reg [(4'hf):(1'h0)] reg1701 = (1'h0);
  reg [(3'h4):(1'h0)] reg1699 = (1'h0);
  reg [(5'h11):(1'h0)] reg1904 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1901 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1899 = (1'h0);
  reg [(5'h17):(1'h0)] reg1898 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1897 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1896 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1895 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1894 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1893 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1891 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1889 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1886 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1883 = (1'h0);
  reg [(5'h10):(1'h0)] reg1882 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1881 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1878 = (1'h0);
  reg [(4'ha):(1'h0)] reg1877 = (1'h0);
  reg [(5'h10):(1'h0)] reg1876 = (1'h0);
  reg [(4'ha):(1'h0)] reg1875 = (1'h0);
  reg [(2'h2):(1'h0)] reg1872 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1871 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1870 = (1'h0);
  reg [(5'h18):(1'h0)] reg1868 = (1'h0);
  reg [(2'h3):(1'h0)] reg1867 = (1'h0);
  reg [(4'hf):(1'h0)] reg1866 = (1'h0);
  reg [(5'h18):(1'h0)] reg1865 = (1'h0);
  reg [(4'hf):(1'h0)] reg1864 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1863 = (1'h0);
  reg [(5'h13):(1'h0)] reg1860 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1859 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1858 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1854 = (1'h0);
  reg [(5'h15):(1'h0)] reg1853 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1851 = (1'h0);
  reg [(3'h5):(1'h0)] reg1849 = (1'h0);
  reg [(2'h3):(1'h0)] reg1848 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1847 = (1'h0);
  reg [(4'ha):(1'h0)] reg1845 = (1'h0);
  reg [(3'h5):(1'h0)] reg1844 = (1'h0);
  reg [(4'ha):(1'h0)] reg1841 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1840 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1839 = (1'h0);
  reg [(2'h2):(1'h0)] reg1838 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1837 = (1'h0);
  reg [(4'ha):(1'h0)] reg1836 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1834 = (1'h0);
  reg [(5'h16):(1'h0)] reg1830 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1824 = (1'h0);
  reg [(4'hf):(1'h0)] reg1823 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1822 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1821 = (1'h0);
  reg [(3'h6):(1'h0)] reg1816 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1815 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1813 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1797 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1796 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1807 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1806 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1805 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1802 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1801 = (1'h0);
  reg [(2'h2):(1'h0)] reg1800 = (1'h0);
  reg [(3'h4):(1'h0)] reg1798 = (1'h0);
  reg [(4'h9):(1'h0)] reg1797 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1796 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1793 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1792 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1772 = (1'h0);
  reg [(4'ha):(1'h0)] reg1771 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1790 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1789 = (1'h0);
  reg [(5'h16):(1'h0)] reg1788 = (1'h0);
  reg [(4'ha):(1'h0)] reg1787 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1783 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1779 = (1'h0);
  reg [(5'h18):(1'h0)] reg1777 = (1'h0);
  reg [(3'h6):(1'h0)] reg1775 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1772 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1771 = (1'h0);
  reg [(3'h5):(1'h0)] reg1770 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1769 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1767 = (1'h0);
  reg [(5'h13):(1'h0)] reg1763 = (1'h0);
  reg [(4'hd):(1'h0)] reg1760 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1759 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1758 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1757 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1755 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1754 = (1'h0);
  reg [(3'h5):(1'h0)] reg1752 = (1'h0);
  reg [(2'h3):(1'h0)] reg1751 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1749 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1745 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1742 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1741 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1740 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1737 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1733 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1731 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1729 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1727 = (1'h0);
  reg [(5'h16):(1'h0)] reg1726 = (1'h0);
  reg [(3'h7):(1'h0)] reg1725 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1724 = (1'h0);
  reg [(5'h15):(1'h0)] reg1723 = (1'h0);
  reg [(3'h7):(1'h0)] reg1722 = (1'h0);
  reg [(5'h14):(1'h0)] reg1721 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1720 = (1'h0);
  reg [(5'h17):(1'h0)] reg1718 = (1'h0);
  reg [(4'hb):(1'h0)] reg1717 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1715 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1713 = (1'h0);
  reg [(4'h8):(1'h0)] reg1712 = (1'h0);
  reg [(5'h10):(1'h0)] reg1709 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1708 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1700 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1698 = (1'h0);
  reg [(3'h6):(1'h0)] reg1697 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1696 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar1695 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1694 = (1'h0);
  assign y = {wire1905,
                 wire1833,
                 wire1832,
                 wire1814,
                 wire1810,
                 wire1809,
                 wire1693,
                 wire1692,
                 reg1903,
                 reg1902,
                 reg1900,
                 reg1892,
                 reg1890,
                 reg1888,
                 reg1887,
                 reg1885,
                 reg1884,
                 reg1880,
                 reg1879,
                 reg1874,
                 reg1873,
                 reg1869,
                 reg1862,
                 reg1861,
                 reg1857,
                 reg1856,
                 reg1855,
                 reg1834,
                 reg1852,
                 reg1850,
                 reg1846,
                 reg1843,
                 reg1842,
                 reg1835,
                 reg1831,
                 reg1829,
                 reg1828,
                 reg1827,
                 reg1826,
                 reg1825,
                 reg1820,
                 reg1819,
                 reg1818,
                 reg1817,
                 reg1812,
                 reg1811,
                 reg1808,
                 reg1804,
                 reg1803,
                 reg1799,
                 reg1795,
                 reg1794,
                 reg1791,
                 reg1786,
                 reg1785,
                 reg1784,
                 reg1782,
                 reg1781,
                 reg1780,
                 reg1778,
                 reg1776,
                 reg1774,
                 reg1773,
                 reg1768,
                 reg1766,
                 reg1765,
                 reg1764,
                 reg1762,
                 reg1761,
                 reg1756,
                 reg1753,
                 reg1750,
                 reg1748,
                 reg1747,
                 reg1746,
                 reg1744,
                 reg1743,
                 reg1739,
                 reg1738,
                 reg1736,
                 reg1735,
                 reg1734,
                 reg1732,
                 reg1730,
                 reg1728,
                 reg1719,
                 reg1716,
                 reg1714,
                 reg1711,
                 reg1710,
                 reg1707,
                 reg1706,
                 reg1705,
                 reg1704,
                 reg1703,
                 reg1702,
                 reg1701,
                 reg1699,
                 reg1904,
                 reg1901,
                 forvar1899,
                 reg1898,
                 forvar1897,
                 reg1896,
                 reg1895,
                 reg1894,
                 reg1893,
                 reg1891,
                 forvar1889,
                 forvar1886,
                 reg1883,
                 reg1882,
                 reg1881,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1875,
                 reg1872,
                 reg1871,
                 reg1870,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1864,
                 forvar1863,
                 reg1860,
                 reg1859,
                 reg1858,
                 reg1854,
                 reg1853,
                 reg1851,
                 reg1849,
                 reg1848,
                 reg1847,
                 reg1845,
                 reg1844,
                 reg1841,
                 reg1840,
                 reg1839,
                 reg1838,
                 reg1837,
                 reg1836,
                 forvar1834,
                 reg1830,
                 reg1824,
                 reg1823,
                 reg1822,
                 reg1821,
                 reg1816,
                 forvar1815,
                 reg1813,
                 forvar1797,
                 reg1796,
                 reg1807,
                 reg1806,
                 reg1805,
                 forvar1802,
                 reg1801,
                 reg1800,
                 reg1798,
                 reg1797,
                 forvar1796,
                 reg1793,
                 reg1792,
                 forvar1772,
                 reg1771,
                 reg1790,
                 reg1789,
                 reg1788,
                 reg1787,
                 reg1783,
                 reg1779,
                 reg1777,
                 reg1775,
                 reg1772,
                 forvar1771,
                 reg1770,
                 reg1769,
                 forvar1767,
                 reg1763,
                 reg1760,
                 reg1759,
                 reg1758,
                 reg1757,
                 forvar1755,
                 reg1754,
                 reg1752,
                 reg1751,
                 reg1749,
                 reg1745,
                 reg1742,
                 forvar1741,
                 forvar1740,
                 reg1737,
                 reg1733,
                 reg1731,
                 reg1729,
                 reg1727,
                 reg1726,
                 reg1725,
                 reg1724,
                 reg1723,
                 reg1722,
                 reg1721,
                 forvar1720,
                 reg1718,
                 reg1717,
                 reg1715,
                 reg1713,
                 reg1712,
                 reg1709,
                 reg1708,
                 reg1700,
                 forvar1698,
                 reg1697,
                 reg1696,
                 forvar1695,
                 reg1694,
                 (1'h0)};
  assign wire1692 = $signed($unsigned(($unsigned($unsigned(wire1688)) ?
                        (^~wire1690[(2'h2):(1'h0)]) : {(wire1689 ?
                                (8'haa) : wire1689),
                            (!wire1690)})));
  assign wire1693 = $signed((($unsigned((wire1690 ?
                        wire1690 : wire1688)) ^ (~|$signed(wire1687))) >= $signed(wire1687)));
  always
    @(posedge clk) begin
      reg1694 = $signed((~|wire1687[(2'h2):(2'h2)]));
    end
  always
    @(posedge clk) begin
      for (forvar1695 = (1'h0); (forvar1695 < (1'h0)); forvar1695 = (forvar1695 + (1'h1)))
        begin
          reg1696 = (((wire1690[(4'ha):(2'h2)] >>> $signed((wire1688 ~^ wire1693))) ?
              ($signed($unsigned(wire1691)) ?
                  (~(forvar1695 | wire1687)) : wire1690) : wire1689[(4'hd):(4'h8)]) ~^ wire1687[(3'h5):(3'h4)]);
          reg1697 = (!{$signed($unsigned($unsigned(wire1687))),
              $unsigned(wire1692[(3'h7):(1'h1)]),
              (~|((+reg1696) != (^~wire1687)))});
          for (forvar1698 = (1'h0); (forvar1698 < (2'h2)); forvar1698 = (forvar1698 + (1'h1)))
            begin
              reg1699 <= wire1690[(4'hf):(2'h2)];
              reg1700 = wire1688;
              reg1701 <= $signed(reg1697[(1'h1):(1'h1)]);
              reg1702 <= $unsigned((&(^~$signed(wire1691[(4'h8):(3'h7)]))));
              reg1703 <= ((({reg1699[(1'h1):(1'h0)]} ?
                      ((reg1702 != wire1692) - (~wire1689)) : reg1696[(4'h8):(3'h5)]) ?
                  wire1689 : (8'haa)) ^~ ($unsigned(wire1691) ^ wire1690));
              reg1704 <= wire1692;
            end
          if (reg1703[(3'h4):(2'h2)])
            begin
              reg1705 <= (forvar1695[(5'h13):(5'h11)] ?
                  $unsigned($signed((^~(!(8'ha6))))) : ($unsigned($unsigned((reg1703 & forvar1695))) == $signed((!forvar1698))));
              reg1706 <= $unsigned({(~^$signed($unsigned((8'hbd)))),
                  {$signed((forvar1698 == wire1689))},
                  $signed(reg1703)});
              reg1707 <= wire1687;
              reg1708 = (forvar1695 ?
                  (+reg1701[(4'ha):(3'h6)]) : $signed((~((forvar1695 ?
                      wire1692 : reg1703) ~^ (|wire1691)))));
              reg1709 = ($unsigned((({(8'hb9), (7'h58), (8'ha3)} ?
                      wire1693[(5'h11):(4'h8)] : (reg1697 == reg1702)) == wire1692)) ?
                  $unsigned($unsigned(reg1702[(5'h15):(4'hf)])) : ($unsigned((^~$unsigned(wire1692))) * (~|$unsigned((~^reg1706)))));
              reg1710 <= ((&forvar1698[(4'he):(4'hb)]) ?
                  $unsigned(reg1707[(4'ha):(4'h9)]) : reg1701[(4'hd):(3'h6)]);
            end
          else
            begin
              reg1705 <= ((($signed((reg1696 ? reg1696 : reg1710)) ?
                      (!wire1688) : (reg1697 >> (reg1706 ?
                          forvar1698 : reg1706))) >= $signed(((reg1697 - wire1688) <<< forvar1695[(2'h2):(1'h0)]))) ?
                  (((reg1706[(1'h0):(1'h0)] ?
                          reg1701 : {(8'hb6),
                              reg1707,
                              wire1688}) << $signed((reg1709 ?
                          reg1696 : wire1690))) ?
                      (~{{wire1692, reg1705},
                          reg1703,
                          $unsigned(reg1701)}) : ($unsigned(reg1701[(4'h9):(4'h8)]) - (|reg1701))) : (7'h41));
            end
          if ($signed(reg1703[(4'h8):(3'h4)]))
            begin
              reg1711 <= ({($signed((-reg1705)) < (reg1702 + $signed(reg1696)))} ?
                  (8'hac) : reg1709);
              reg1712 = $unsigned(wire1692);
              reg1713 = reg1699[(1'h1):(1'h1)];
            end
          else
            begin
              reg1712 = $unsigned(reg1713);
              reg1714 <= {reg1705, reg1702, wire1689};
              reg1715 = (^((&$signed(wire1687)) >= reg1703[(3'h5):(3'h4)]));
              reg1716 <= ((&(((reg1708 != reg1697) ? reg1711 : (~reg1699)) ?
                  ($unsigned(reg1715) ?
                      $unsigned(reg1697) : reg1699) : ((reg1706 ^ reg1709) < reg1705[(1'h0):(1'h0)]))) - reg1700[(3'h4):(1'h1)]);
              reg1717 = (-{{wire1691[(3'h5):(1'h1)],
                      reg1696[(3'h4):(1'h1)],
                      (((8'ha4) <<< reg1715) ?
                          {reg1716, wire1687} : (wire1693 ?
                              reg1704 : wire1690))}});
              reg1718 = (reg1701 ?
                  {(7'h55)} : $signed((reg1702[(4'ha):(3'h7)] ?
                      (-reg1709[(3'h6):(2'h2)]) : $signed(((8'ha7) >= reg1708)))));
            end
          reg1719 <= $unsigned((~(($signed(wire1687) ?
              $signed(reg1699) : {reg1708,
                  (8'hb9),
                  reg1708}) != $signed({reg1711, reg1713, (7'h58)}))));
          for (forvar1720 = (1'h0); (forvar1720 < (2'h2)); forvar1720 = (forvar1720 + (1'h1)))
            begin
              reg1721 = ((($unsigned($signed(reg1709)) * reg1697) ?
                  wire1692[(3'h4):(3'h4)] : $signed((|$unsigned((7'h46))))) << {$signed(reg1715),
                  (~(~|(reg1699 ? reg1706 : (7'h46)))),
                  reg1705[(3'h6):(3'h4)]});
              reg1722 = $signed($signed((|((reg1711 | wire1690) <= $unsigned(reg1718)))));
              reg1723 = $unsigned(((8'ha2) ?
                  (reg1712 && $signed($unsigned((8'ha7)))) : reg1717[(3'h5):(2'h2)]));
              reg1724 = ((^reg1718) ?
                  $unsigned($unsigned($signed($unsigned(reg1722)))) : forvar1720[(5'h10):(4'hb)]);
              reg1725 = $unsigned((-{((reg1702 ? forvar1698 : (7'h4a)) ?
                      $signed(forvar1695) : reg1717[(4'h8):(4'h8)]),
                  ($signed(wire1693) >> (reg1716 ? reg1716 : reg1701)),
                  (^~$signed(reg1708))}));
              reg1726 = ((-$signed($signed($unsigned(reg1724)))) <<< {(reg1721[(3'h5):(2'h2)] ^ (~(~reg1705))),
                  wire1687,
                  (~^{{reg1700, (8'ha6), reg1705},
                      ((8'hb0) || forvar1695),
                      {reg1701, reg1714}})});
            end
        end
      if ({reg1721,
          $unsigned($unsigned((wire1689[(5'h12):(4'h8)] ?
              {(7'h4a)} : reg1718)))})
        begin
          reg1727 = {(~^{reg1705, reg1726, reg1717})};
          reg1728 <= $signed(($unsigned($unsigned((&reg1718))) ?
              $unsigned($unsigned(reg1727)) : (reg1712[(3'h7):(3'h4)] | reg1717[(3'h7):(1'h0)])));
        end
      else
        begin
          if ($unsigned(reg1710[(1'h0):(1'h0)]))
            begin
              reg1727 = ({reg1699,
                  (reg1728[(3'h7):(3'h7)] ?
                      ((wire1690 == reg1726) == $unsigned(forvar1720)) : $signed(wire1688[(5'h13):(4'hf)])),
                  {reg1704,
                      (reg1703 ? forvar1698[(4'he):(4'hc)] : (~&reg1719)),
                      (+$signed(wire1692))}} <<< ($unsigned($unsigned(forvar1695[(5'h12):(2'h3)])) > {forvar1695[(3'h6):(3'h6)],
                  forvar1695,
                  $unsigned($unsigned((7'h41)))}));
              reg1729 = ($unsigned($unsigned(($unsigned(reg1706) ?
                  $signed(wire1690) : (reg1715 <= reg1713)))) && (+(^~(8'hb5))));
            end
          else
            begin
              reg1727 = {{$unsigned((8'hb5)), reg1715}};
              reg1729 = (wire1692 ?
                  {{reg1696[(4'h9):(1'h0)],
                          $unsigned(forvar1695[(5'h1c):(5'h1b)]),
                          ($signed(reg1712) ?
                              {reg1725,
                                  reg1724} : ((8'ha4) * (8'ha9)))}} : (~reg1728));
              reg1730 <= reg1728;
              reg1731 = $unsigned(wire1687[(3'h5):(1'h1)]);
              reg1732 <= (&reg1722);
              reg1733 = ({$signed(($unsigned(reg1721) ?
                          $signed((8'ha9)) : {(8'h9f), reg1717}))} ?
                  wire1687[(1'h1):(1'h0)] : $signed($unsigned(reg1718[(1'h1):(1'h0)])));
              reg1734 <= $unsigned((8'ha7));
            end
          reg1735 <= ($signed($signed(wire1687[(2'h2):(2'h2)])) || reg1700[(2'h3):(2'h3)]);
          reg1736 <= reg1724;
          reg1737 = reg1730[(5'h12):(4'h8)];
          reg1738 <= (((|($unsigned(reg1734) >>> (&reg1724))) ?
              (~reg1731) : (|(reg1701 ?
                  $signed(reg1733) : {reg1730}))) ^ reg1734[(1'h1):(1'h0)]);
          reg1739 <= reg1721;
        end
      for (forvar1740 = (1'h0); (forvar1740 < (2'h3)); forvar1740 = (forvar1740 + (1'h1)))
        begin
          for (forvar1741 = (1'h0); (forvar1741 < (2'h3)); forvar1741 = (forvar1741 + (1'h1)))
            begin
              reg1742 = $signed(reg1722);
              reg1743 <= $unsigned($signed((((reg1733 + forvar1698) ?
                      (reg1702 ? reg1725 : reg1699) : $signed(reg1725)) ?
                  $signed(reg1701[(4'ha):(2'h2)]) : (&reg1712))));
              reg1744 <= $signed($unsigned(reg1723));
              reg1745 = {reg1711[(4'h9):(2'h2)], reg1702[(4'hd):(4'hc)]};
              reg1746 <= {reg1701,
                  (|{(^~wire1692[(3'h4):(2'h2)]),
                      $signed((~wire1690)),
                      wire1688[(3'h6):(3'h4)]}),
                  $unsigned($unsigned(reg1730))};
              reg1747 <= (reg1726[(2'h2):(1'h0)] ?
                  {reg1727} : (reg1730[(3'h5):(3'h5)] || $unsigned($unsigned((+(8'hb7))))));
            end
          if ({reg1703[(2'h3):(1'h1)], reg1722[(1'h1):(1'h1)]})
            begin
              reg1748 <= reg1743[(3'h5):(1'h0)];
              reg1749 = ((reg1706 ?
                  $unsigned(reg1735[(4'hc):(4'h9)]) : $unsigned((reg1727 ?
                      (!forvar1740) : reg1726[(4'hc):(3'h5)]))) >> $unsigned($unsigned((^reg1702[(4'h8):(3'h7)]))));
              reg1750 <= wire1692[(4'ha):(1'h1)];
              reg1751 = (~&{((reg1699[(2'h3):(2'h3)] <= reg1749) ?
                      (reg1724[(3'h5):(1'h0)] ^ reg1710) : ((~&reg1710) <<< wire1691)),
                  reg1737,
                  reg1746[(5'h16):(4'h9)]});
              reg1752 = reg1749;
            end
          else
            begin
              reg1748 <= (&$unsigned(reg1750));
              reg1749 = reg1700[(3'h5):(1'h1)];
            end
          reg1753 <= reg1708[(5'h18):(5'h11)];
          reg1754 = reg1709;
          for (forvar1755 = (1'h0); (forvar1755 < (3'h4)); forvar1755 = (forvar1755 + (1'h1)))
            begin
              reg1756 <= {((((reg1724 != reg1730) << reg1737) ^ (&(wire1691 ^~ reg1738))) != $unsigned($unsigned(((8'hb6) < reg1749))))};
              reg1757 = $signed($unsigned(reg1738[(3'h5):(2'h3)]));
              reg1758 = $signed((((reg1757 ? (~&(8'hb2)) : reg1717) ?
                      reg1719 : {wire1693[(3'h4):(2'h2)], (&forvar1720)}) ?
                  $signed($unsigned({reg1704,
                      reg1712,
                      reg1719})) : (&($signed(reg1744) | $unsigned((8'hbc))))));
              reg1759 = (reg1731 ?
                  ($signed((wire1693 >>> reg1701)) && $signed((~|(reg1753 - reg1746)))) : (-(~&($signed(reg1757) ^ $signed(forvar1695)))));
              reg1760 = (reg1704 ?
                  reg1713[(3'h4):(3'h4)] : $unsigned((~|($signed(reg1699) ^~ (+reg1739)))));
              reg1761 <= reg1723[(5'h10):(1'h1)];
              reg1762 <= reg1723;
            end
          reg1763 = reg1696;
        end
      reg1764 <= $signed($unsigned({{$signed(reg1754)},
          $signed($unsigned(reg1752))}));
      reg1765 <= reg1746[(3'h6):(2'h2)];
    end
  always
    @(posedge clk) begin
      reg1766 <= (wire1690 ? reg1750 : {reg1728[(3'h5):(1'h0)]});
      for (forvar1767 = (1'h0); (forvar1767 < (2'h3)); forvar1767 = (forvar1767 + (1'h1)))
        begin
          reg1768 <= {(reg1711 ? reg1748 : (~&$signed((|(8'had)))))};
        end
      reg1769 = ((reg1702 <<< (~&{(~(8'hab))})) >> reg1705[(2'h3):(2'h3)]);
      reg1770 = forvar1767;
    end
  always
    @(posedge clk) begin
      if ({$unsigned((~&(8'hbc))),
          {(~&$signed($unsigned(wire1689)))},
          $unsigned({((reg1728 ? (7'h53) : reg1746) ?
                  (&reg1735) : reg1711[(5'h12):(3'h7)]),
              $signed((reg1728 << reg1739)),
              $unsigned($unsigned(reg1701))})})
        begin
          for (forvar1771 = (1'h0); (forvar1771 < (3'h6)); forvar1771 = (forvar1771 + (1'h1)))
            begin
              reg1772 = ((wire1688[(4'he):(3'h6)] ?
                  (!$unsigned((reg1739 >= (8'ha5)))) : reg1765) ^~ ($unsigned(reg1738[(3'h5):(2'h2)]) ?
                  (-($signed(reg1701) ?
                      $unsigned(reg1704) : (reg1747 ~^ wire1691))) : ((~^$unsigned(reg1719)) ?
                      ((reg1739 >>> reg1703) + {wire1690}) : wire1690)));
              reg1773 <= reg1716[(1'h0):(1'h0)];
              reg1774 <= ($signed($signed(((reg1703 | reg1701) ^ (reg1739 ?
                  reg1711 : reg1753)))) <<< $signed($signed((reg1765[(2'h3):(1'h0)] >>> {reg1744,
                  wire1691,
                  (8'h9d)}))));
              reg1775 = reg1748;
              reg1776 <= wire1693[(4'hf):(1'h1)];
            end
          if ($unsigned(($unsigned((reg1761[(5'h16):(4'hd)] ?
              wire1688[(5'h16):(3'h4)] : {reg1735,
                  reg1747,
                  reg1734})) <<< (reg1705[(2'h2):(1'h0)] ?
              (8'hb7) : $signed(reg1762)))))
            begin
              reg1777 = $unsigned(((wire1693 ?
                  reg1716 : $unsigned((~reg1736))) + $unsigned((^~(reg1773 + reg1701)))));
              reg1778 <= (|(reg1735[(1'h1):(1'h1)] ~^ $unsigned((^wire1692))));
              reg1779 = ($signed(reg1728[(4'h9):(4'h9)]) ~^ $signed(reg1774));
              reg1780 <= reg1766[(2'h3):(1'h0)];
              reg1781 <= wire1689;
              reg1782 <= $signed(($signed(reg1711[(5'h17):(4'hc)]) | $unsigned(reg1710[(4'hf):(4'hf)])));
              reg1783 = reg1702[(2'h2):(1'h0)];
            end
          else
            begin
              reg1778 <= ((reg1735[(4'hb):(2'h3)] && ($unsigned(reg1768) == $unsigned((reg1781 ~^ reg1719)))) ?
                  (-reg1746[(4'hd):(2'h3)]) : $unsigned(reg1702[(4'hf):(2'h3)]));
              reg1780 <= $signed((reg1730 == (reg1780[(3'h5):(2'h3)] || $unsigned(reg1732))));
              reg1781 <= $signed($signed($unsigned(reg1732[(3'h5):(3'h5)])));
              reg1782 <= $unsigned((+$signed(wire1688)));
              reg1784 <= ((((&$signed(reg1756)) ?
                      wire1687[(4'h8):(2'h2)] : reg1704) >= reg1716[(3'h7):(3'h6)]) ?
                  wire1691[(3'h6):(3'h6)] : ($unsigned(wire1689[(4'hd):(4'h9)]) ?
                      (|(reg1719[(1'h0):(1'h0)] ?
                          (reg1744 | reg1777) : (wire1693 >>> reg1707))) : (|$unsigned((reg1748 ?
                          reg1710 : reg1773)))));
              reg1785 <= reg1782[(2'h3):(2'h3)];
              reg1786 <= $signed($signed((((reg1746 ~^ reg1711) >>> reg1784[(4'h9):(4'h9)]) >= reg1703)));
            end
          reg1787 = reg1699[(1'h1):(1'h0)];
          if ((-{reg1732[(4'he):(4'hd)],
              ({(+(8'h9c)),
                  wire1690[(1'h0):(1'h0)],
                  (reg1756 ? reg1702 : reg1738)} <= $signed((reg1738 ?
                  reg1739 : reg1776)))}))
            begin
              reg1788 = reg1707;
              reg1789 = (reg1739 ?
                  $unsigned(reg1773) : $signed((-$signed((^~(8'hb4))))));
            end
          else
            begin
              reg1788 = (($signed(($signed(reg1761) >>> (reg1736 ?
                      reg1774 : reg1714))) ?
                  reg1702 : reg1762) <<< ({(!$signed((8'ha0)))} > (^~$unsigned((~&reg1781)))));
              reg1789 = (~&{$unsigned(reg1730)});
            end
          reg1790 = $signed(wire1687[(4'ha):(2'h2)]);
          reg1791 <= (-$unsigned(((^$signed(reg1732)) ?
              (-reg1789) : (!{reg1732, wire1689, reg1764}))));
        end
      else
        begin
          reg1771 = reg1784[(3'h4):(1'h0)];
          for (forvar1772 = (1'h0); (forvar1772 < (1'h0)); forvar1772 = (forvar1772 + (1'h1)))
            begin
              reg1775 = reg1702[(2'h3):(2'h2)];
              reg1777 = ($signed($unsigned($signed((~&reg1732)))) + ((-($unsigned(reg1735) ?
                  (reg1776 == reg1766) : reg1703)) < ($unsigned((reg1773 ?
                  forvar1772 : wire1689)) >= reg1705)));
              reg1778 <= reg1784[(4'h9):(3'h5)];
            end
          if (reg1789)
            begin
              reg1780 <= (((8'ha3) ?
                      $signed($unsigned($signed(reg1753))) : ((7'h47) < {$unsigned(reg1743),
                          (wire1691 ~^ reg1730)})) ?
                  ((reg1789[(5'h11):(5'h11)] ?
                          reg1766 : reg1705[(1'h1):(1'h1)]) ?
                      (((reg1775 < reg1777) ?
                          $unsigned(reg1738) : (reg1778 ?
                              wire1691 : reg1702)) | reg1790) : $signed($signed(((8'ha0) ^~ forvar1772)))) : $unsigned($unsigned(($unsigned(reg1701) << $signed(reg1744)))));
              reg1783 = (+reg1732);
              reg1784 <= reg1734[(1'h0):(1'h0)];
              reg1785 <= $signed(reg1766);
            end
          else
            begin
              reg1779 = wire1691[(1'h1):(1'h0)];
              reg1780 <= $unsigned($unsigned({reg1771[(1'h1):(1'h0)],
                  reg1714,
                  ((~^reg1707) ~^ reg1787[(1'h0):(1'h0)])}));
              reg1781 <= reg1736[(5'h11):(3'h6)];
              reg1782 <= ((reg1747[(1'h1):(1'h1)] ?
                      {reg1734,
                          ((reg1719 == reg1748) >>> (+wire1689)),
                          $unsigned(reg1773)} : $unsigned(reg1743)) ?
                  (~^$signed({(|reg1764),
                      (8'hbf),
                      (reg1776 >= wire1692)})) : ($unsigned($signed($unsigned((8'ha8)))) ?
                      {(!(reg1704 < (8'hb6))),
                          ({reg1736,
                              reg1710} >= reg1707)} : (reg1711 * (reg1744 && ((7'h45) && wire1689)))));
            end
          if ({$signed($signed(reg1773)),
              (~&(&((wire1687 ? reg1704 : (7'h41)) ?
                  (reg1762 ? reg1768 : reg1738) : reg1784[(4'hd):(4'hc)])))})
            begin
              reg1786 <= reg1734[(1'h1):(1'h0)];
              reg1787 = reg1771;
            end
          else
            begin
              reg1787 = reg1771[(3'h7):(3'h6)];
              reg1788 = reg1786[(3'h5):(2'h2)];
              reg1789 = {{(~|$unsigned($signed((8'h9d)))),
                      $signed($signed($unsigned(reg1705)))},
                  $signed($unsigned((~$signed((7'h49)))))};
              reg1791 <= (~^($signed((+(reg1785 ?
                  reg1773 : reg1736))) <= ($unsigned(forvar1771) ?
                  ((reg1736 == reg1766) ?
                      {(8'h9d), reg1777} : {reg1778,
                          (8'hbd),
                          reg1761}) : $signed(reg1714))));
              reg1792 = ($signed((^$unsigned(reg1719))) >>> forvar1772[(4'hc):(3'h6)]);
              reg1793 = reg1787;
              reg1794 <= (reg1747 ?
                  ((~&(!(~^reg1783))) ?
                      (reg1784[(4'hc):(3'h5)] ?
                          reg1748 : reg1785) : (~^(wire1693 == reg1791))) : {(~&reg1719)});
            end
          reg1795 <= ((forvar1772[(4'hb):(4'hb)] ?
              (~^reg1736[(5'h14):(2'h2)]) : $unsigned($signed(((8'ha6) * reg1706)))) && reg1734[(1'h0):(1'h0)]);
        end
      if ({(|(^($unsigned(reg1778) | (7'h42))))})
        begin
          for (forvar1796 = (1'h0); (forvar1796 < (3'h5)); forvar1796 = (forvar1796 + (1'h1)))
            begin
              reg1797 = reg1768[(1'h0):(1'h0)];
              reg1798 = reg1739;
              reg1799 <= reg1771[(2'h2):(1'h0)];
              reg1800 = (~&((reg1773 ?
                  $signed(((8'hb3) > (8'hb2))) : (7'h4e)) && (reg1795[(5'h1c):(1'h0)] ?
                  (8'h9f) : (~|(reg1785 ? reg1799 : reg1795)))));
              reg1801 = ((7'h4f) < {(8'hb7),
                  (((reg1784 != reg1795) ?
                      reg1728[(3'h6):(3'h6)] : (reg1736 ?
                          reg1719 : wire1693)) << (!reg1773)),
                  {(~&(~&reg1787))}});
            end
          for (forvar1802 = (1'h0); (forvar1802 < (3'h4)); forvar1802 = (forvar1802 + (1'h1)))
            begin
              reg1803 <= $signed((&$signed((reg1707[(5'h10):(1'h1)] ?
                  $unsigned(reg1738) : reg1703))));
              reg1804 <= ($unsigned(reg1788[(5'h10):(4'he)]) >> (reg1738[(3'h4):(3'h4)] ?
                  (($unsigned(reg1732) ?
                      reg1743 : {reg1756,
                          (8'ha8)}) < $signed(wire1688[(5'h12):(5'h12)])) : $signed((^~reg1705))));
              reg1805 = $unsigned(($unsigned(reg1762[(4'hb):(2'h2)]) ^~ (&reg1794)));
              reg1806 = (^$signed(($signed(reg1784) ?
                  reg1775[(3'h4):(2'h3)] : (~^reg1711))));
              reg1807 = ((reg1777[(5'h14):(1'h1)] - $signed(reg1785[(3'h6):(3'h4)])) ?
                  (reg1728 < reg1710[(4'h8):(3'h7)]) : ((!reg1793) ?
                      wire1693 : (~$unsigned(reg1768))));
            end
        end
      else
        begin
          reg1796 = reg1805[(3'h7):(3'h5)];
          for (forvar1797 = (1'h0); (forvar1797 < (3'h5)); forvar1797 = (forvar1797 + (1'h1)))
            begin
              reg1798 = ((reg1719 >>> $signed($unsigned((~|reg1739)))) ?
                  reg1707 : (reg1800 ?
                      ((7'h47) ?
                          reg1750 : ((~^(8'hae)) ?
                              $unsigned(reg1711) : ((7'h4c) ?
                                  reg1711 : wire1693))) : (($unsigned((8'ha0)) ?
                          reg1703 : (reg1801 ?
                              (8'ha6) : reg1764)) || reg1766)));
              reg1799 <= $unsigned($signed(((-(reg1753 << (7'h49))) ?
                  $signed((~reg1772)) : (reg1747[(1'h0):(1'h0)] ?
                      wire1690 : (reg1699 ? reg1799 : reg1728)))));
            end
        end
      reg1808 <= $signed($unsigned(reg1738));
    end
  assign wire1809 = $unsigned((|$signed(reg1701)));
  assign wire1810 = ((+$signed(reg1703)) ?
                        $unsigned(reg1706[(4'h9):(4'h9)]) : $unsigned($signed(((!reg1716) >>> $unsigned(reg1701)))));
  always
    @(posedge clk) begin
      reg1811 <= $signed((($signed((-wire1693)) <= ((reg1784 == reg1711) ?
              $unsigned(reg1699) : {(8'h9d), reg1768, reg1799})) ?
          ($signed((reg1781 ? reg1778 : (8'hb4))) ?
              (wire1810[(4'h8):(2'h2)] == reg1706) : reg1701) : $unsigned((+(reg1748 - reg1756)))));
      if ((7'h56))
        begin
          reg1812 <= (((!$unsigned({(7'h54)})) ?
              (~^(reg1738[(2'h2):(1'h1)] ^~ reg1795)) : reg1743[(2'h2):(2'h2)]) >>> ($unsigned($unsigned((reg1808 ?
              reg1795 : reg1766))) >>> (-(wire1809 ? reg1738 : reg1778))));
        end
      else
        begin
          reg1812 <= reg1710[(4'hd):(4'hd)];
        end
      reg1813 = reg1732[(5'h10):(1'h1)];
    end
  assign wire1814 = reg1804[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar1815 = (1'h0); (forvar1815 < (1'h0)); forvar1815 = (forvar1815 + (1'h1)))
        begin
          if ((^$unsigned((^reg1785))))
            begin
              reg1816 = (~|(reg1784 && $signed(reg1732)));
              reg1817 <= {$unsigned($unsigned({(~|reg1774), reg1701})),
                  ((~^(reg1753[(5'h19):(5'h12)] ^ {wire1690,
                          reg1816,
                          wire1691})) ?
                      $unsigned(reg1710) : reg1781)};
              reg1818 <= $signed($signed($unsigned(reg1746)));
              reg1819 <= {$signed({(~|reg1799[(3'h4):(1'h0)]),
                      ($signed(wire1687) >= $unsigned(reg1704)),
                      reg1707[(5'h11):(3'h5)]})};
              reg1820 <= $signed($unsigned(($unsigned(reg1716) ?
                  $unsigned((reg1764 <= reg1784)) : $unsigned(reg1799[(2'h2):(1'h0)]))));
            end
          else
            begin
              reg1816 = $unsigned((~|$signed((^$signed(reg1778)))));
              reg1817 <= reg1794;
              reg1818 <= (reg1803[(4'h9):(3'h7)] ?
                  ((({reg1780, reg1716} ? ((8'hbd) * reg1711) : reg1699) ?
                      (wire1689[(5'h1b):(5'h12)] ?
                          $signed(reg1768) : $signed(reg1750)) : reg1739[(3'h7):(3'h6)]) + $signed(reg1812)) : $signed((~|$unsigned((reg1699 ?
                      reg1750 : reg1703)))));
              reg1821 = ($unsigned($unsigned(((|reg1753) || reg1808[(3'h7):(3'h5)]))) ^~ reg1816);
              reg1822 = $unsigned(wire1810);
            end
          if (wire1810[(3'h4):(2'h2)])
            begin
              reg1823 = $unsigned(reg1735[(4'ha):(1'h0)]);
              reg1824 = (^$signed(($unsigned($signed(reg1773)) == $signed((^reg1739)))));
            end
          else
            begin
              reg1825 <= wire1814;
              reg1826 <= (wire1687 > $signed({{(reg1764 ? reg1728 : (7'h49)),
                      {reg1819, reg1703, reg1750},
                      (reg1730 ? reg1710 : wire1687)},
                  {reg1761[(3'h6):(3'h6)]}}));
              reg1827 <= (~(+$unsigned(wire1809)));
              reg1828 <= wire1693[(1'h1):(1'h0)];
            end
          reg1829 <= $signed(({(7'h57),
                  ((reg1817 ? reg1750 : reg1786) ^~ reg1817),
                  $unsigned((forvar1815 >>> reg1819))} ?
              {reg1794[(5'h12):(2'h2)]} : $signed(({reg1827} ?
                  $unsigned(reg1828) : {reg1794, reg1699, wire1687}))));
          reg1830 = (($signed(((reg1746 ? reg1773 : reg1746) ?
                  (reg1773 ?
                      reg1748 : (8'hb4)) : reg1716)) < reg1732[(3'h4):(2'h3)]) ?
              $unsigned((~|(-$signed(reg1762)))) : ((^$signed(reg1728[(4'ha):(4'h8)])) & {reg1820[(1'h0):(1'h0)],
                  $signed($signed(reg1702))}));
          reg1831 <= (reg1743 >>> (&$signed($signed((reg1748 ?
              wire1687 : reg1819)))));
        end
    end
  assign wire1832 = $signed($signed((-(reg1761[(5'h10):(4'hb)] & wire1690[(4'hf):(4'he)]))));
  assign wire1833 = ((~&{{$unsigned(reg1735)}}) != reg1827[(2'h2):(1'h0)]);
  always
    @(posedge clk) begin
      if (((((reg1703[(3'h6):(3'h6)] ? (7'h44) : reg1812[(3'h5):(3'h5)]) ?
                  ((wire1693 ?
                      wire1690 : (8'ha1)) * reg1784[(4'h9):(2'h2)]) : {(reg1702 ?
                          reg1747 : (8'hac)),
                      $unsigned(reg1786)}) ?
              (+(&reg1781)) : (^~((~^wire1688) ?
                  ((8'hbc) >>> reg1773) : reg1829[(4'hf):(4'hf)]))) ?
          (+(($unsigned(reg1831) ? wire1692 : $signed(reg1764)) ?
              ({reg1739, reg1703, (8'hbb)} ?
                  $signed(reg1831) : (+reg1706)) : (reg1702[(3'h4):(1'h0)] ?
                  (reg1826 ?
                      reg1711 : reg1773) : (reg1780 * reg1719)))) : {reg1762[(2'h2):(1'h0)],
              reg1768}))
        begin
          for (forvar1834 = (1'h0); (forvar1834 < (3'h4)); forvar1834 = (forvar1834 + (1'h1)))
            begin
              reg1835 <= $unsigned({$signed(reg1780), $signed(reg1761)});
              reg1836 = $signed((wire1832 ?
                  {$unsigned((reg1820 <= reg1803)),
                      reg1812} : wire1688[(5'h1c):(4'h9)]));
              reg1837 = {$unsigned((reg1705 ?
                      ((^reg1812) ?
                          (~&wire1689) : wire1814[(5'h10):(4'hb)]) : reg1766[(2'h3):(1'h0)]))};
              reg1838 = (reg1818[(5'h18):(1'h1)] != (reg1714 < ($unsigned((^~reg1812)) ?
                  reg1748[(3'h4):(2'h3)] : reg1744[(1'h0):(1'h0)])));
              reg1839 = (~|$unsigned(reg1773));
              reg1840 = (reg1719[(1'h1):(1'h0)] ?
                  ($signed(reg1739) ?
                      (|{reg1828[(3'h5):(2'h3)],
                          reg1825}) : reg1817) : reg1766[(3'h5):(3'h4)]);
              reg1841 = $unsigned({{(|reg1819), (~|$signed(reg1753))},
                  $unsigned(($unsigned(reg1839) ?
                      (reg1785 ? (8'hb6) : reg1744) : ((8'ha0) ~^ reg1739)))});
            end
          reg1842 <= ((($signed($unsigned(reg1703)) << ($unsigned(wire1688) ?
                  (wire1809 ? reg1794 : (8'hbf)) : wire1687)) ?
              reg1738[(1'h0):(1'h0)] : ($unsigned((reg1732 <<< reg1795)) || $signed((reg1714 ?
                  reg1744 : reg1838)))) != ($unsigned($unsigned((~&reg1782))) ?
              $signed(reg1799[(2'h3):(1'h1)]) : (7'h47)));
          if (forvar1834[(4'h9):(3'h5)])
            begin
              reg1843 <= $unsigned($unsigned($unsigned($unsigned({(8'ha6),
                  reg1756}))));
              reg1844 = (~^reg1841);
              reg1845 = $unsigned(reg1786);
              reg1846 <= $unsigned((reg1839 ~^ ($unsigned((&reg1812)) ?
                  $unsigned(reg1836[(1'h1):(1'h0)]) : {(^reg1835),
                      $unsigned(reg1804),
                      (reg1828 ? reg1719 : reg1845)})));
              reg1847 = (reg1836[(2'h2):(1'h1)] ?
                  $unsigned(reg1778) : (^~reg1819));
              reg1848 = (8'ha8);
              reg1849 = (&(&{(reg1728 ? $signed((7'h49)) : wire1689),
                  reg1703,
                  reg1706}));
            end
          else
            begin
              reg1844 = ((|reg1748[(3'h4):(1'h0)]) ?
                  reg1840 : reg1811[(5'h12):(3'h7)]);
              reg1846 <= {$signed((reg1828[(3'h5):(1'h1)] ?
                      {reg1753} : ($signed((8'ha8)) << (~^reg1702)))),
                  $signed(reg1736)};
              reg1847 = (8'hac);
              reg1850 <= ((&{reg1785}) + (~^{{(^reg1776), (!wire1688)}}));
              reg1851 = (($signed((~|$unsigned(wire1688))) ?
                      reg1818 : ((~&$unsigned(reg1734)) - reg1835[(4'hc):(2'h3)])) ?
                  $signed((reg1841[(2'h2):(1'h1)] ~^ reg1838[(2'h2):(1'h0)])) : (^(7'h52)));
            end
          reg1852 <= (~|({{reg1780[(3'h4):(1'h0)],
                      $unsigned(reg1838),
                      reg1773[(2'h2):(1'h0)]},
                  {(reg1704 ? reg1848 : reg1730), reg1761[(5'h11):(4'h8)]}} ?
              (reg1743[(2'h3):(2'h2)] * $unsigned((+reg1764))) : ((!(8'hb1)) * reg1778[(3'h4):(1'h0)])));
          reg1853 = (~|reg1746);
        end
      else
        begin
          reg1834 <= $signed($unsigned(reg1808));
        end
      if (reg1743[(3'h4):(1'h1)])
        begin
          if ($signed($signed(reg1710)))
            begin
              reg1854 = reg1795[(4'hf):(1'h0)];
              reg1855 <= $signed(($unsigned(((~reg1827) >= (reg1719 | reg1719))) ?
                  reg1704 : ({$unsigned(reg1825)} < $unsigned({wire1691,
                      reg1736}))));
              reg1856 <= $unsigned((~^reg1702));
              reg1857 <= ((!(reg1707 && ($unsigned(reg1819) | wire1832))) >> (reg1736[(5'h10):(3'h5)] > reg1747));
              reg1858 = (reg1811 & (reg1837 != (~^((|reg1743) << (reg1705 << reg1748)))));
              reg1859 = (((reg1826 ?
                      $unsigned((7'h40)) : (!(+reg1838))) > $signed(($unsigned(reg1702) == ((8'ha7) ?
                      reg1773 : wire1810)))) ?
                  reg1811 : reg1735);
              reg1860 = {(&$signed(forvar1834[(4'hb):(2'h2)])),
                  reg1811,
                  reg1811[(4'hf):(4'h9)]};
            end
          else
            begin
              reg1855 <= $signed((reg1728[(1'h1):(1'h1)] ?
                  reg1773[(2'h3):(1'h0)] : reg1850));
              reg1856 <= $unsigned($unsigned(((8'had) ?
                  ($signed((7'h51)) ?
                      reg1829[(5'h13):(2'h2)] : $unsigned(reg1860)) : (-((7'h41) == reg1780)))));
              reg1857 <= {(^(|reg1854)), (~|reg1716[(3'h5):(3'h4)])};
              reg1858 = {reg1703[(3'h7):(2'h3)],
                  wire1692[(4'h9):(4'h9)],
                  (reg1795 ?
                      $unsigned({$unsigned(reg1856),
                          reg1753[(4'hb):(1'h1)],
                          $signed(wire1690)}) : $signed(((^reg1837) ?
                          reg1857 : reg1826[(1'h0):(1'h0)])))};
            end
        end
      else
        begin
          if ($signed(reg1846[(1'h0):(1'h0)]))
            begin
              reg1855 <= (reg1804[(2'h2):(1'h1)] ?
                  reg1781[(5'h17):(1'h1)] : $unsigned(((reg1711[(5'h12):(4'hf)] & $unsigned(reg1706)) + $signed((wire1687 <<< reg1716)))));
              reg1858 = $signed($signed((((~&reg1705) ^ reg1730[(1'h0):(1'h0)]) ?
                  {reg1852[(5'h19):(3'h5)]} : (~|$unsigned((7'h53))))));
              reg1861 <= wire1810;
              reg1862 <= ((8'hae) ?
                  $unsigned((reg1838[(1'h1):(1'h0)] > {((7'h41) >> (8'hab)),
                      $signed(reg1811)})) : wire1814);
            end
          else
            begin
              reg1854 = reg1780[(3'h4):(1'h0)];
            end
          for (forvar1863 = (1'h0); (forvar1863 < (3'h6)); forvar1863 = (forvar1863 + (1'h1)))
            begin
              reg1864 = reg1781[(5'h18):(5'h14)];
              reg1865 = reg1854[(3'h7):(3'h7)];
              reg1866 = $signed((+reg1837));
              reg1867 = $signed($unsigned($unsigned(reg1852[(5'h17):(4'hd)])));
              reg1868 = (~|reg1827[(2'h2):(1'h1)]);
              reg1869 <= (reg1747 ?
                  $signed((({(8'hb7), (8'h9f), reg1699} ?
                          $unsigned(reg1716) : (8'hb8)) ?
                      (8'h9e) : reg1791)) : reg1719[(4'h8):(2'h3)]);
            end
          if ($unsigned((^~(7'h51))))
            begin
              reg1870 = $unsigned({$unsigned(reg1705),
                  $unsigned(reg1851),
                  (reg1799[(3'h4):(2'h3)] ?
                      (reg1748 ?
                          (reg1705 ?
                              reg1738 : reg1825) : (^reg1743)) : $signed({reg1765,
                          wire1810}))});
              reg1871 = (reg1773[(1'h1):(1'h0)] ?
                  ($unsigned(reg1778) <= (reg1841 ?
                      reg1860 : ((reg1829 >>> reg1746) ?
                          $unsigned(reg1710) : reg1852))) : (~^($unsigned({(7'h40),
                          reg1784}) ?
                      $unsigned(reg1811) : $signed($unsigned(reg1786)))));
              reg1872 = reg1768;
            end
          else
            begin
              reg1870 = reg1820[(4'hb):(3'h7)];
              reg1871 = ($unsigned(reg1852[(5'h19):(1'h1)]) ?
                  reg1867[(2'h2):(2'h2)] : reg1766);
              reg1872 = $unsigned((~|(~^($unsigned(reg1861) >> (reg1736 & reg1869)))));
              reg1873 <= reg1836;
              reg1874 <= reg1861;
              reg1875 = reg1845;
              reg1876 = reg1762[(4'hc):(4'hb)];
            end
          if (($signed((reg1784[(1'h0):(1'h0)] << $unsigned(reg1765))) ?
              $signed((^((reg1773 ?
                  reg1819 : (8'ha1)) == $unsigned(reg1719)))) : ({$signed((reg1704 ?
                          reg1780 : reg1828)),
                      wire1833[(4'h8):(3'h6)]} ?
                  reg1747[(1'h0):(1'h0)] : ($unsigned((reg1851 & wire1814)) ?
                      $signed($unsigned(reg1835)) : reg1795))))
            begin
              reg1877 = {(^~(((reg1858 ?
                      reg1773 : (8'hb9)) <= {reg1703}) <<< (((7'h51) >> reg1710) ?
                      reg1855 : wire1688)))};
              reg1878 = ($unsigned((~(7'h48))) >> {reg1876[(5'h10):(4'hc)],
                  ((-reg1828) ?
                      ((reg1704 ? (8'hb7) : (8'ha9)) ?
                          (reg1856 < reg1705) : reg1876) : $unsigned((reg1836 ?
                          reg1842 : reg1819)))});
              reg1879 <= {$unsigned($signed($unsigned(reg1719)))};
              reg1880 <= reg1774[(5'h13):(3'h7)];
              reg1881 = (({reg1878,
                  (reg1858[(5'h17):(5'h10)] ?
                      wire1809[(5'h1a):(5'h1a)] : (reg1781 ?
                          reg1728 : reg1817))} && $unsigned((~$signed(reg1808)))) ^ (~&{($unsigned(reg1753) <<< $signed(reg1831))}));
              reg1882 = {reg1850, reg1876[(2'h3):(2'h2)]};
              reg1883 = ($signed(({(reg1870 ^ wire1810),
                      ((8'hac) | reg1756)} && $signed((reg1711 ?
                      reg1866 : (7'h46))))) ?
                  ({$unsigned((&reg1704)),
                          $unsigned($unsigned(reg1865)),
                          $signed({reg1706})} ?
                      reg1835[(4'he):(4'hb)] : ((((8'hba) ^~ reg1761) << ((8'ha6) ?
                              reg1808 : reg1730)) ?
                          reg1864 : $signed((~^(8'hb4))))) : $unsigned({(|reg1774)}));
            end
          else
            begin
              reg1879 <= $signed((~&({(8'hb6),
                  (+reg1837),
                  reg1707[(4'hd):(3'h7)]} >>> reg1875)));
              reg1881 = (|$unsigned($signed($signed($signed(reg1706)))));
              reg1884 <= (reg1849 == ($unsigned(((reg1875 <= reg1869) ?
                      reg1762[(3'h4):(1'h1)] : reg1738[(1'h0):(1'h0)])) ?
                  reg1843[(5'h19):(3'h7)] : (!((~|(7'h4b)) ?
                      $unsigned(reg1781) : reg1786))));
            end
          reg1885 <= $signed(({(wire1691 > $signed(forvar1834))} + (reg1874[(3'h7):(3'h7)] ^ $signed((|reg1876)))));
          for (forvar1886 = (1'h0); (forvar1886 < (1'h1)); forvar1886 = (forvar1886 + (1'h1)))
            begin
              reg1887 <= reg1826[(2'h2):(2'h2)];
              reg1888 <= reg1836;
            end
          for (forvar1889 = (1'h0); (forvar1889 < (3'h6)); forvar1889 = (forvar1889 + (1'h1)))
            begin
              reg1890 <= (wire1814[(5'h19):(4'h8)] ?
                  {$signed($unsigned(reg1732[(4'hf):(4'hd)]))} : reg1882);
              reg1891 = $unsigned(reg1859);
              reg1892 <= ({$unsigned(((reg1890 | reg1846) ?
                      $unsigned(reg1804) : reg1840[(5'h11):(4'he)]))} > ((-$signed((^~wire1688))) != $unsigned((reg1865[(5'h13):(5'h13)] ?
                  (+reg1843) : reg1881))));
              reg1893 = (!$unsigned($unsigned($unsigned($unsigned(reg1880)))));
              reg1894 = ((|reg1876) - $unsigned($signed($unsigned(((8'hab) ?
                  reg1744 : reg1880)))));
              reg1895 = reg1710;
              reg1896 = $unsigned(($unsigned((wire1814 ^ {(8'hb9),
                  reg1891,
                  reg1702})) ^~ $signed((reg1744 & (wire1814 ?
                  reg1865 : wire1693)))));
            end
        end
      for (forvar1897 = (1'h0); (forvar1897 < (3'h4)); forvar1897 = (forvar1897 + (1'h1)))
        begin
          reg1898 = (-(-$unsigned($signed(reg1744[(2'h2):(2'h2)]))));
          for (forvar1899 = (1'h0); (forvar1899 < (3'h5)); forvar1899 = (forvar1899 + (1'h1)))
            begin
              reg1900 <= reg1882;
              reg1901 = (~|$signed($unsigned($unsigned($signed(reg1799)))));
              reg1902 <= (|reg1875[(1'h0):(1'h0)]);
            end
          reg1903 <= (~|({$signed($signed((8'hb8)))} ? reg1699 : reg1714));
          reg1904 = {$signed($signed(($unsigned(wire1809) ^ (reg1812 ?
                  reg1845 : (8'hb8)))))};
        end
    end
  assign wire1905 = reg1747;
endmodule