(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param776 = (|((((^(8'hbe)) < ((8'hb4) ~^ (7'h40))) && ((^(8'hb7)) ? ((8'hbf) ? (8'hae) : (8'hbb)) : ((8'h9e) ? (8'hb6) : (8'hb7)))) <<< (&(-(~|(8'hb6)))))))
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h33a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire4;
  input wire [(5'h11):(1'h0)] wire3;
  input wire [(4'hb):(1'h0)] wire2;
  input wire signed [(3'h5):(1'h0)] wire1;
  input wire signed [(4'ha):(1'h0)] wire0;
  wire [(3'h5):(1'h0)] wire775;
  wire [(5'h10):(1'h0)] wire774;
  wire signed [(3'h7):(1'h0)] wire773;
  wire signed [(5'h15):(1'h0)] wire772;
  wire [(3'h4):(1'h0)] wire771;
  wire signed [(3'h5):(1'h0)] wire770;
  wire signed [(2'h2):(1'h0)] wire769;
  wire signed [(4'hd):(1'h0)] wire768;
  wire signed [(2'h3):(1'h0)] wire767;
  wire signed [(2'h2):(1'h0)] wire766;
  wire signed [(3'h7):(1'h0)] wire765;
  wire [(5'h11):(1'h0)] wire764;
  wire signed [(5'h11):(1'h0)] wire709;
  wire signed [(4'h8):(1'h0)] wire708;
  wire [(4'he):(1'h0)] wire707;
  wire signed [(5'h15):(1'h0)] wire706;
  wire signed [(4'hd):(1'h0)] wire705;
  wire [(4'hd):(1'h0)] wire704;
  wire signed [(4'h9):(1'h0)] wire703;
  wire [(4'he):(1'h0)] wire702;
  wire [(5'h13):(1'h0)] wire700;
  reg signed [(5'h13):(1'h0)] reg761 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg759 = (1'h0);
  reg [(3'h7):(1'h0)] reg758 = (1'h0);
  reg [(4'he):(1'h0)] reg756 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg752 = (1'h0);
  reg [(4'h8):(1'h0)] reg750 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg748 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg747 = (1'h0);
  reg [(4'hb):(1'h0)] reg744 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg742 = (1'h0);
  reg [(4'hf):(1'h0)] reg741 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg739 = (1'h0);
  reg [(3'h4):(1'h0)] reg737 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg735 = (1'h0);
  reg [(4'he):(1'h0)] reg734 = (1'h0);
  reg [(3'h7):(1'h0)] reg733 = (1'h0);
  reg [(3'h7):(1'h0)] reg730 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg726 = (1'h0);
  reg [(5'h13):(1'h0)] reg725 = (1'h0);
  reg [(2'h2):(1'h0)] reg722 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg721 = (1'h0);
  reg [(2'h3):(1'h0)] reg719 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg717 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg714 = (1'h0);
  reg [(2'h3):(1'h0)] reg710 = (1'h0);
  reg [(3'h6):(1'h0)] reg711 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg763 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg762 = (1'h0);
  reg [(3'h4):(1'h0)] reg760 = (1'h0);
  reg [(3'h6):(1'h0)] forvar757 = (1'h0);
  reg [(5'h14):(1'h0)] reg755 = (1'h0);
  reg [(4'he):(1'h0)] reg754 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg753 = (1'h0);
  reg [(5'h12):(1'h0)] forvar751 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg749 = (1'h0);
  reg [(5'h13):(1'h0)] forvar746 = (1'h0);
  reg [(5'h15):(1'h0)] reg745 = (1'h0);
  reg [(3'h4):(1'h0)] reg743 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar740 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg738 = (1'h0);
  reg signed [(4'he):(1'h0)] reg736 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg732 = (1'h0);
  reg [(4'he):(1'h0)] reg731 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg729 = (1'h0);
  reg [(4'h8):(1'h0)] reg728 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg727 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg724 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg723 = (1'h0);
  reg [(4'h8):(1'h0)] reg720 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar718 = (1'h0);
  reg [(5'h10):(1'h0)] reg716 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg713 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg712 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar710 = (1'h0);
  assign y = {wire775,
                 wire774,
                 wire773,
                 wire772,
                 wire771,
                 wire770,
                 wire769,
                 wire768,
                 wire767,
                 wire766,
                 wire765,
                 wire764,
                 wire709,
                 wire708,
                 wire707,
                 wire706,
                 wire705,
                 wire704,
                 wire703,
                 wire702,
                 wire700,
                 reg761,
                 reg759,
                 reg758,
                 reg756,
                 reg752,
                 reg750,
                 reg748,
                 reg747,
                 reg744,
                 reg742,
                 reg741,
                 reg739,
                 reg737,
                 reg735,
                 reg734,
                 reg733,
                 reg730,
                 reg726,
                 reg725,
                 reg722,
                 reg721,
                 reg719,
                 reg717,
                 reg715,
                 reg714,
                 reg710,
                 reg711,
                 reg763,
                 reg762,
                 reg760,
                 forvar757,
                 reg755,
                 reg754,
                 reg753,
                 forvar751,
                 reg749,
                 forvar746,
                 reg745,
                 reg743,
                 forvar740,
                 reg738,
                 reg736,
                 reg732,
                 reg731,
                 reg729,
                 reg728,
                 reg727,
                 reg724,
                 reg723,
                 reg720,
                 forvar718,
                 reg716,
                 reg713,
                 reg712,
                 forvar710,
                 (1'h0)};
  module5 #() modinst701 (.wire9(wire0), .y(wire700), .clk(clk), .wire7(wire2), .wire6(wire3), .wire8(wire4));
  assign wire702 = $unsigned({wire1[(2'h2):(1'h1)], wire1});
  assign wire703 = (({wire0[(1'h0):(1'h0)], wire4[(4'h8):(1'h1)]} ?
                           $unsigned(wire702[(4'hd):(4'hb)]) : (+wire4[(4'h8):(1'h0)])) ?
                       $signed((wire702[(2'h2):(1'h0)] ?
                           (8'hb6) : ($signed(wire702) ?
                               wire3[(3'h6):(3'h6)] : (wire4 | wire3)))) : $signed($unsigned((wire4[(3'h5):(2'h2)] ?
                           (wire3 * (7'h40)) : {wire2, wire700}))));
  assign wire704 = $unsigned($unsigned(($signed((wire702 ? wire1 : wire1)) ?
                       $unsigned(wire4[(4'ha):(2'h2)]) : (~$signed(wire700)))));
  assign wire705 = $unsigned(wire700[(5'h12):(5'h12)]);
  assign wire706 = (wire705 ?
                       ((wire702 ?
                           {(wire704 ? wire700 : wire702),
                               wire4[(3'h7):(3'h6)]} : (wire0[(3'h5):(1'h0)] && (~|wire700))) | (wire705 || $signed((&wire702)))) : (8'ha8));
  assign wire707 = $signed({(wire705 ?
                           wire0[(4'h8):(3'h6)] : {wire704[(4'h8):(1'h0)],
                               (~&wire3)})});
  assign wire708 = wire702;
  assign wire709 = wire702[(3'h7):(1'h1)];
  always
    @(posedge clk) begin
      if ($signed($unsigned(wire2[(3'h5):(1'h1)])))
        begin
          for (forvar710 = (1'h0); (forvar710 < (2'h3)); forvar710 = (forvar710 + (1'h1)))
            begin
              reg711 <= $signed(wire3);
            end
        end
      else
        begin
          if ((($signed(($unsigned(forvar710) ?
              (wire1 >= wire704) : {wire1})) <= ((~^(wire703 - (8'hb5))) + ((wire707 & wire703) <<< $unsigned(wire2)))) || $unsigned((((wire705 + (8'hb4)) == $unsigned(wire2)) ?
              $unsigned(wire708) : wire702))))
            begin
              reg710 <= (!$unsigned($signed((wire706[(4'hb):(3'h7)] + ((8'hb2) ?
                  forvar710 : wire702)))));
              reg711 <= {$unsigned($unsigned($unsigned(((8'h9f) ?
                      wire702 : wire709))))};
              reg712 = $signed(wire4[(4'h9):(3'h6)]);
              reg713 = $signed((8'hb2));
              reg714 <= (reg712[(3'h7):(3'h4)] | (~|(wire1[(2'h2):(1'h1)] <<< {wire707})));
            end
          else
            begin
              reg710 <= $signed($unsigned(($unsigned(wire704[(4'ha):(4'ha)]) ?
                  ((8'hba) || (wire706 ?
                      reg712 : wire704)) : $unsigned(reg714))));
            end
          if (($unsigned((reg711[(1'h0):(1'h0)] ?
              wire707[(2'h3):(1'h1)] : ((8'hb2) ?
                  $unsigned(wire708) : $unsigned(reg711)))) > ($signed((+(wire709 ^~ wire708))) ?
              wire703[(3'h7):(1'h0)] : ((wire704[(4'h8):(3'h5)] >> {(8'hbc),
                  reg714}) >= (reg713 < (wire707 & wire709))))))
            begin
              reg715 <= wire708[(3'h7):(1'h1)];
              reg716 = $signed((~(~|((~&wire702) > (reg714 < reg713)))));
              reg717 <= $signed($signed($signed($unsigned($signed(wire709)))));
            end
          else
            begin
              reg715 <= $signed((-forvar710));
            end
          for (forvar718 = (1'h0); (forvar718 < (2'h2)); forvar718 = (forvar718 + (1'h1)))
            begin
              reg719 <= ({(~&wire706[(3'h7):(2'h3)]),
                  {((wire706 < reg714) || (wire700 >= wire3))}} << $unsigned($unsigned(($signed(forvar710) & (reg716 < wire3)))));
              reg720 = wire1;
              reg721 <= {(reg713[(1'h1):(1'h1)] ?
                      wire702[(4'hd):(3'h7)] : $unsigned($unsigned((~reg710)))),
                  wire703};
            end
          if ($unsigned(wire702[(4'h9):(3'h5)]))
            begin
              reg722 <= (~&{(8'hb5)});
            end
          else
            begin
              reg723 = $unsigned(reg717[(1'h1):(1'h1)]);
              reg724 = reg719;
              reg725 <= ($unsigned(reg722) ^~ $signed(((~|((8'hb6) ?
                  (8'hb8) : wire3)) <= ((reg711 ?
                  wire709 : reg711) ^~ wire0[(1'h1):(1'h0)]))));
              reg726 <= wire703[(2'h3):(1'h0)];
              reg727 = (+$unsigned(reg714[(3'h5):(1'h1)]));
            end
        end
      if ((wire4[(4'h8):(3'h4)] * (wire707 ?
          $signed($signed(reg726)) : (((wire703 ? reg723 : (8'ha4)) ?
              $signed(reg710) : (~^reg719)) ^ (^(~^reg723))))))
        begin
          if (($signed(((8'hbe) ?
                  ((!reg725) ?
                      (wire702 ?
                          (8'ha2) : wire702) : (~|reg723)) : $unsigned($unsigned(wire709)))) ?
              reg717[(1'h0):(1'h0)] : (reg716 ^ reg714)))
            begin
              reg728 = (wire706 || reg717[(1'h1):(1'h1)]);
              reg729 = (8'ha7);
            end
          else
            begin
              reg728 = reg713[(3'h5):(2'h3)];
              reg730 <= {(~|(~($unsigned(reg717) ?
                      (~(8'hb0)) : (reg724 ? (8'hac) : reg722))))};
              reg731 = reg714[(1'h0):(1'h0)];
              reg732 = $signed((((wire705[(4'hc):(4'h9)] == reg711) >= (^wire2[(2'h2):(1'h1)])) ?
                  $unsigned(reg728) : {($unsigned((8'ha6)) ?
                          $unsigned((7'h42)) : wire4)}));
              reg733 <= reg732[(2'h2):(1'h0)];
            end
          reg734 <= ($signed($unsigned({$unsigned(reg720),
              ((8'ha7) != (8'h9c))})) != $signed((($unsigned(reg725) ?
                  (wire1 ^ reg714) : reg722) ?
              wire706[(5'h15):(5'h11)] : ($signed(reg710) << (wire703 << (8'h9c))))));
        end
      else
        begin
          if ({{(((wire706 ? reg732 : reg726) ?
                          (~^reg716) : (wire0 < wire702)) ?
                      $signed((reg722 ? reg725 : wire703)) : ((reg727 ?
                          reg715 : reg727) << reg716)),
                  wire707[(4'he):(4'hb)]}})
            begin
              reg728 = (((!$signed((reg720 ?
                  wire709 : wire1))) >> reg722) == ((~|wire4[(4'h9):(1'h1)]) != ($unsigned({wire705}) && reg717)));
              reg730 <= reg717;
              reg733 <= {wire706[(4'he):(3'h7)]};
              reg734 <= ($unsigned($signed(reg726)) ?
                  (^(^~(reg711 >>> (reg723 ?
                      reg728 : reg723)))) : (-{$signed((wire708 + reg729)),
                      wire1[(1'h0):(1'h0)]}));
              reg735 <= reg712;
            end
          else
            begin
              reg728 = ($unsigned((wire700 ?
                      $unsigned(reg730[(3'h4):(2'h2)]) : (~|(reg719 > (8'hba))))) ?
                  (|$unsigned(((wire3 >= (8'hba)) ?
                      $unsigned(reg711) : reg716[(4'h8):(3'h6)]))) : (reg715[(4'h9):(2'h3)] * wire703[(1'h0):(1'h0)]));
            end
          if ($signed($unsigned($unsigned(wire707[(4'h9):(3'h6)]))))
            begin
              reg736 = (8'ha5);
            end
          else
            begin
              reg737 <= (reg721 ?
                  $unsigned(reg735) : $unsigned((wire703 || $signed((^reg721)))));
              reg738 = ({wire702[(3'h5):(3'h4)]} ?
                  reg730 : (~($signed((reg729 && reg737)) ?
                      ($signed(wire4) & $signed(reg713)) : $unsigned($unsigned(reg732)))));
              reg739 <= reg730[(1'h0):(1'h0)];
            end
        end
      for (forvar740 = (1'h0); (forvar740 < (1'h0)); forvar740 = (forvar740 + (1'h1)))
        begin
          if ((^~$unsigned(({reg733} || reg721[(5'h10):(4'he)]))))
            begin
              reg741 <= wire704[(4'hc):(2'h3)];
              reg742 <= $unsigned($unsigned($unsigned(forvar718[(5'h11):(4'hb)])));
              reg743 = $signed($signed($unsigned(reg724[(2'h3):(2'h3)])));
            end
          else
            begin
              reg741 <= {reg733[(3'h7):(3'h4)], wire709[(4'ha):(2'h3)]};
              reg743 = ((wire704 ?
                  reg714[(4'h8):(3'h7)] : reg743) == wire707[(3'h7):(2'h2)]);
              reg744 <= {reg714};
              reg745 = ($signed(((8'hb3) ?
                  (((8'ha8) && (8'ha3)) ?
                      reg710[(2'h3):(1'h0)] : (~&wire702)) : $unsigned((reg721 ?
                      wire1 : (8'hb9))))) >= $unsigned((reg743[(2'h2):(1'h0)] ?
                  (+$unsigned((8'hb9))) : $unsigned((8'hb1)))));
            end
          for (forvar746 = (1'h0); (forvar746 < (3'h4)); forvar746 = (forvar746 + (1'h1)))
            begin
              reg747 <= {wire709[(3'h6):(3'h5)], reg732[(4'h8):(2'h2)]};
              reg748 <= ($signed(forvar710[(3'h6):(3'h5)]) - $unsigned($signed((|(&wire705)))));
              reg749 = ($signed((($signed(reg739) == ((8'h9d) | reg717)) ?
                  (((8'h9e) <<< reg715) - $unsigned(wire2)) : {(reg734 + (8'hb9)),
                      $signed(reg717)})) & reg748[(3'h4):(2'h3)]);
              reg750 <= ((~^{reg745[(4'ha):(3'h6)],
                  ((8'hac) ?
                      $unsigned((8'hb1)) : {reg710})}) && $signed(($unsigned({forvar718,
                  (8'hae)}) * ((reg744 ? wire4 : reg721) ?
                  $signed((8'ha8)) : (+wire0)))));
            end
          for (forvar751 = (1'h0); (forvar751 < (2'h2)); forvar751 = (forvar751 + (1'h1)))
            begin
              reg752 <= reg728;
              reg753 = ($signed((!(reg735 ?
                  (^wire4) : $unsigned((8'had))))) && forvar710);
              reg754 = ({{reg726, (&reg730[(3'h6):(1'h1)])},
                      $unsigned(wire709[(4'h8):(3'h4)])} ?
                  {((8'h9f) ?
                          $signed(reg714[(4'h9):(2'h3)]) : (reg734 ?
                              (wire702 != forvar710) : (reg738 ?
                                  reg735 : reg732)))} : (^~$signed((!reg745[(4'hf):(4'hb)]))));
              reg755 = (~(-(reg748 ? (~forvar751) : reg729[(1'h0):(1'h0)])));
              reg756 <= (^wire4);
            end
        end
      for (forvar757 = (1'h0); (forvar757 < (2'h3)); forvar757 = (forvar757 + (1'h1)))
        begin
          if ($signed(reg717))
            begin
              reg758 <= {(^reg733),
                  $signed($unsigned($unsigned((wire703 ?
                      reg745 : forvar751))))};
              reg759 <= wire700[(4'h8):(2'h2)];
            end
          else
            begin
              reg758 <= reg738[(4'ha):(3'h4)];
              reg760 = reg734;
              reg761 <= ((^~reg724) < $signed((((wire706 ?
                      (8'haa) : forvar710) ?
                  (|reg728) : (reg716 + reg728)) + $unsigned((reg743 < wire709)))));
              reg762 = (wire700[(5'h12):(4'hb)] ?
                  {$unsigned({reg724[(4'hf):(4'hc)]})} : forvar751);
            end
          reg763 = forvar710[(1'h1):(1'h0)];
        end
    end
  assign wire764 = ((wire707[(4'h8):(2'h2)] ?
                       reg734 : ({(~&wire4)} ?
                           (+(~&reg725)) : ($signed((8'hbc)) ?
                               reg714 : ((8'hbb) > reg711)))) || $unsigned(reg748[(3'h7):(3'h7)]));
  assign wire765 = reg735;
  assign wire766 = ($unsigned(($signed(reg719) ?
                           reg737[(2'h2):(2'h2)] : reg750)) ?
                       (~&reg734[(3'h4):(2'h2)]) : $signed(($signed($unsigned(wire703)) >= reg730)));
  assign wire767 = ($unsigned({{(^~reg722),
                           $signed((8'ha0))}}) | wire703[(4'h9):(1'h0)]);
  assign wire768 = (+(&{$signed((&reg726)),
                       {reg741[(3'h6):(2'h3)], reg719[(1'h0):(1'h0)]}}));
  assign wire769 = {reg752,
                       {$unsigned(reg744),
                           (^{wire765, ((7'h44) ? reg722 : wire3)})}};
  assign wire770 = reg742;
  assign wire771 = wire707[(4'ha):(3'h4)];
  assign wire772 = reg719[(1'h0):(1'h0)];
  assign wire773 = wire0;
  assign wire774 = $signed((reg730 << $signed($unsigned($signed(reg761)))));
  assign wire775 = ($unsigned((^($signed(wire769) < (wire709 >= reg756)))) ?
                       wire700[(4'hc):(4'h8)] : $signed({$signed({wire0})}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5  (y, clk, wire6, wire7, wire8, wire9);
  output wire [(32'h55a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire6;
  input wire signed [(4'hb):(1'h0)] wire7;
  input wire [(4'hb):(1'h0)] wire8;
  input wire signed [(4'ha):(1'h0)] wire9;
  wire [(5'h12):(1'h0)] wire557;
  wire [(4'he):(1'h0)] wire315;
  wire [(5'h11):(1'h0)] wire10;
  wire signed [(5'h10):(1'h0)] wire11;
  wire [(4'hc):(1'h0)] wire12;
  wire signed [(3'h7):(1'h0)] wire61;
  wire [(4'hc):(1'h0)] wire62;
  wire signed [(4'hd):(1'h0)] wire63;
  wire signed [(4'ha):(1'h0)] wire117;
  wire [(3'h7):(1'h0)] wire118;
  wire signed [(3'h7):(1'h0)] wire313;
  wire [(4'h9):(1'h0)] wire559;
  wire signed [(4'he):(1'h0)] wire698;
  reg signed [(5'h15):(1'h0)] reg116 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg115 = (1'h0);
  reg [(3'h6):(1'h0)] reg114 = (1'h0);
  reg [(2'h3):(1'h0)] reg112 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg111 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg108 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg103 = (1'h0);
  reg [(3'h5):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg96 = (1'h0);
  reg [(5'h15):(1'h0)] reg94 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg93 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg92 = (1'h0);
  reg [(3'h5):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg86 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg84 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg83 = (1'h0);
  reg [(4'hb):(1'h0)] reg82 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg79 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg78 = (1'h0);
  reg [(5'h15):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg73 = (1'h0);
  reg [(4'ha):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg68 = (1'h0);
  reg [(4'hc):(1'h0)] reg67 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg65 = (1'h0);
  reg [(5'h10):(1'h0)] reg60 = (1'h0);
  reg [(5'h13):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg54 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg50 = (1'h0);
  reg [(3'h7):(1'h0)] reg48 = (1'h0);
  reg [(4'h9):(1'h0)] reg47 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg45 = (1'h0);
  reg [(5'h14):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg43 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg40 = (1'h0);
  reg [(5'h12):(1'h0)] reg38 = (1'h0);
  reg [(5'h11):(1'h0)] reg37 = (1'h0);
  reg [(4'ha):(1'h0)] reg36 = (1'h0);
  reg [(4'he):(1'h0)] reg34 = (1'h0);
  reg [(3'h5):(1'h0)] reg33 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg30 = (1'h0);
  reg [(5'h13):(1'h0)] reg29 = (1'h0);
  reg [(4'hc):(1'h0)] reg28 = (1'h0);
  reg [(3'h5):(1'h0)] reg27 = (1'h0);
  reg [(4'he):(1'h0)] reg25 = (1'h0);
  reg [(5'h15):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg21 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg18 = (1'h0);
  reg [(3'h7):(1'h0)] reg17 = (1'h0);
  reg [(4'h8):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg15 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg113 = (1'h0);
  reg [(5'h13):(1'h0)] reg110 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg109 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg106 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar105 = (1'h0);
  reg [(4'hc):(1'h0)] reg104 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg102 = (1'h0);
  reg [(5'h12):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg100 = (1'h0);
  reg [(5'h14):(1'h0)] forvar98 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg97 = (1'h0);
  reg [(4'hf):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg91 = (1'h0);
  reg [(3'h6):(1'h0)] forvar90 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg88 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg87 = (1'h0);
  reg [(5'h10):(1'h0)] reg85 = (1'h0);
  reg [(4'hd):(1'h0)] reg80 = (1'h0);
  reg [(2'h2):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg76 = (1'h0);
  reg [(4'he):(1'h0)] reg75 = (1'h0);
  reg [(5'h15):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg70 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg69 = (1'h0);
  reg [(5'h14):(1'h0)] forvar66 = (1'h0);
  reg [(5'h15):(1'h0)] reg64 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar43 = (1'h0);
  reg [(5'h12):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar56 = (1'h0);
  reg [(3'h6):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg51 = (1'h0);
  reg [(4'ha):(1'h0)] reg49 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg46 = (1'h0);
  reg [(4'h8):(1'h0)] reg42 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg39 = (1'h0);
  reg [(5'h11):(1'h0)] reg35 = (1'h0);
  reg [(2'h3):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar32 = (1'h0);
  reg [(5'h11):(1'h0)] reg31 = (1'h0);
  reg [(4'h8):(1'h0)] reg26 = (1'h0);
  reg [(2'h2):(1'h0)] reg24 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg22 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg19 = (1'h0);
  reg [(4'hb):(1'h0)] reg14 = (1'h0);
  reg [(4'hf):(1'h0)] forvar13 = (1'h0);
  assign y = {wire557,
                 wire315,
                 wire10,
                 wire11,
                 wire12,
                 wire61,
                 wire62,
                 wire63,
                 wire117,
                 wire118,
                 wire313,
                 wire559,
                 wire698,
                 reg116,
                 reg115,
                 reg114,
                 reg112,
                 reg111,
                 reg108,
                 reg103,
                 reg99,
                 reg96,
                 reg94,
                 reg93,
                 reg92,
                 reg89,
                 reg86,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg79,
                 reg78,
                 reg74,
                 reg73,
                 reg72,
                 reg68,
                 reg67,
                 reg65,
                 reg60,
                 reg59,
                 reg58,
                 reg55,
                 reg54,
                 reg50,
                 reg48,
                 reg47,
                 reg45,
                 reg44,
                 reg43,
                 reg41,
                 reg40,
                 reg38,
                 reg37,
                 reg36,
                 reg34,
                 reg33,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg25,
                 reg23,
                 reg21,
                 reg20,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg113,
                 reg110,
                 reg109,
                 reg107,
                 reg106,
                 forvar105,
                 reg104,
                 reg102,
                 reg101,
                 reg100,
                 forvar98,
                 reg97,
                 reg95,
                 reg91,
                 forvar90,
                 reg88,
                 reg87,
                 reg85,
                 reg80,
                 reg77,
                 reg76,
                 reg75,
                 reg71,
                 reg70,
                 reg69,
                 forvar66,
                 reg64,
                 forvar43,
                 reg57,
                 forvar56,
                 reg53,
                 reg52,
                 reg51,
                 reg49,
                 reg46,
                 reg42,
                 reg39,
                 reg35,
                 reg32,
                 forvar32,
                 reg31,
                 reg26,
                 reg24,
                 reg22,
                 reg19,
                 reg14,
                 forvar13,
                 (1'h0)};
  assign wire10 = $signed(wire7[(2'h3):(2'h2)]);
  assign wire11 = (^wire9);
  assign wire12 = wire8;
  always
    @(posedge clk) begin
      for (forvar13 = (1'h0); (forvar13 < (2'h3)); forvar13 = (forvar13 + (1'h1)))
        begin
          reg14 = $unsigned($unsigned((8'hbd)));
          if ($signed(forvar13[(3'h7):(3'h5)]))
            begin
              reg15 <= forvar13;
              reg16 <= $signed({{$signed(reg14[(2'h2):(1'h1)]), reg14}});
              reg17 <= $unsigned(wire6[(1'h1):(1'h1)]);
              reg18 <= (({wire10[(1'h1):(1'h1)],
                      forvar13} | wire8[(4'ha):(3'h7)]) ?
                  $unsigned((~|wire7[(3'h4):(2'h2)])) : $unsigned($signed({(~^reg14),
                      $signed(wire8)})));
            end
          else
            begin
              reg15 <= wire12;
            end
          reg19 = ($signed((wire6 <<< reg16)) ? wire10 : reg16[(3'h5):(3'h4)]);
        end
      reg20 <= ((8'hbd) & ($signed(wire8) ^~ reg16[(3'h6):(3'h5)]));
      if ($unsigned(($unsigned((~|(8'hb7))) ?
          $signed(($unsigned(reg15) <= (reg18 > wire9))) : (reg17[(3'h7):(1'h1)] || (7'h41)))))
        begin
          if ((wire12[(1'h1):(1'h0)] ?
              ({wire7[(3'h5):(2'h3)]} ?
                  (^~(8'hae)) : (((wire6 * reg15) ?
                          (reg18 > reg20) : wire6[(2'h3):(2'h3)]) ?
                      $signed((wire12 ^ wire7)) : wire9)) : wire9[(2'h2):(1'h1)]))
            begin
              reg21 <= wire10;
              reg22 = ($signed((((7'h41) ?
                      ((8'hb7) ?
                          reg21 : (8'hac)) : $unsigned(reg20)) | $signed($unsigned(reg14)))) ?
                  $unsigned(({{(8'hb6), (8'hbd)}, $unsigned(wire10)} ?
                      $signed((reg16 ? reg21 : reg19)) : ($signed((8'hbd)) ?
                          $unsigned(reg19) : $signed(wire11)))) : reg17[(1'h1):(1'h1)]);
              reg23 <= ((({reg16} ?
                  ((reg19 ?
                      reg22 : (8'h9c)) >= (8'ha9)) : ((~&wire12) >>> (reg16 && reg16))) ^ {(~|(reg20 || wire11)),
                  reg19[(4'hb):(3'h7)]}) | $signed(reg21[(4'hf):(3'h5)]));
              reg24 = $signed((reg15 ~^ (+reg14)));
              reg25 <= ((^{(wire9 ? reg20[(1'h1):(1'h1)] : (^~reg23)),
                      wire11}) ?
                  (+reg20) : $unsigned(($unsigned((!(8'haa))) > $unsigned(wire11))));
            end
          else
            begin
              reg22 = $signed((($unsigned((~^wire6)) + ($signed(reg18) > (|(8'hb6)))) ^ $unsigned((wire6 < $unsigned(forvar13)))));
              reg23 <= (({($signed((8'ha1)) || $unsigned(reg17)),
                      (!reg22[(3'h4):(2'h2)])} ?
                  reg24[(1'h0):(1'h0)] : (~$unsigned(reg16))) >>> (!(|(wire11 < {wire9}))));
              reg24 = ((($signed(reg18[(3'h6):(2'h3)]) ?
                  {(reg17 >= reg23)} : (|forvar13[(4'hc):(4'h8)])) << {$signed($unsigned((8'hb3))),
                  $unsigned((8'hac))}) >>> ((^~$signed($signed(wire12))) << (wire7 + ($signed(reg25) ?
                  $signed(wire10) : $unsigned(wire11)))));
            end
          if ($unsigned((&(~|$signed((~&reg17))))))
            begin
              reg26 = (8'hb4);
              reg27 <= $signed((8'ha0));
              reg28 <= ((~^wire10) ?
                  reg19[(2'h2):(2'h2)] : ($signed(reg15) + ((-(~reg25)) ?
                      ((reg17 != reg24) ?
                          reg16[(1'h0):(1'h0)] : $unsigned(wire11)) : (((8'hb1) ?
                              reg21 : forvar13) ?
                          (reg24 ? reg21 : reg20) : (&(8'had))))));
              reg29 <= reg20[(1'h1):(1'h0)];
              reg30 <= (reg16 ?
                  wire12[(3'h4):(2'h3)] : (reg19 ?
                      $signed(((wire9 ?
                          wire10 : wire10) >= (reg17 & wire7))) : $signed(((reg22 <= wire12) ?
                          $signed(reg23) : $signed(reg29)))));
            end
          else
            begin
              reg27 <= {(reg19[(1'h0):(1'h0)] ?
                      reg23[(5'h11):(3'h6)] : ($unsigned((reg17 * wire12)) ?
                          {(wire10 - reg30)} : {reg25})),
                  {(~|$signed((reg18 >= wire11))),
                      ($unsigned(reg22) ? reg29 : (reg20 ? wire8 : reg15))}};
              reg31 = ((8'ha7) < {($unsigned($unsigned(reg22)) ?
                      reg16 : reg23[(2'h2):(1'h1)]),
                  (reg28[(3'h5):(1'h0)] && $unsigned((^reg25)))});
            end
          for (forvar32 = (1'h0); (forvar32 < (2'h2)); forvar32 = (forvar32 + (1'h1)))
            begin
              reg33 <= (!(^($signed(wire12) ?
                  $signed(reg21[(4'hf):(1'h0)]) : $signed(reg25[(4'hd):(4'h9)]))));
            end
        end
      else
        begin
          if ($signed($unsigned($signed($signed((wire12 ? (8'hbd) : wire7))))))
            begin
              reg21 <= (forvar32 <= (+(8'hb6)));
              reg23 <= ({$signed({$unsigned(wire8), (~reg21)}),
                  (+$signed($signed(reg24)))} < $signed(((~(reg18 ?
                      forvar13 : reg21)) ?
                  ($unsigned(reg27) ?
                      reg31 : (reg14 ?
                          reg16 : (8'hb3))) : reg14[(4'ha):(4'ha)])));
              reg24 = reg16;
            end
          else
            begin
              reg21 <= $unsigned(reg30[(2'h3):(1'h1)]);
            end
          reg26 = reg17[(3'h4):(1'h0)];
          if ($signed(($unsigned((8'hb7)) ?
              ($signed($signed(wire8)) ?
                  reg25[(4'h9):(2'h3)] : (reg28 ?
                      (8'ha6) : {reg17})) : $signed((+$signed(wire8))))))
            begin
              reg31 = $unsigned(wire6);
            end
          else
            begin
              reg31 = (~&wire9);
              reg32 = $signed((~^reg19));
              reg33 <= wire6;
              reg34 <= reg24;
            end
        end
      if (($signed(((~(~^forvar32)) ?
          ($unsigned(wire9) ~^ $unsigned(reg34)) : ((wire12 >> reg21) & {(8'hb1)}))) >>> $unsigned($unsigned(((reg19 << (7'h41)) > reg25)))))
        begin
          reg35 = wire12[(1'h0):(1'h0)];
        end
      else
        begin
          if ({$unsigned(($unsigned(reg20) ?
                  (reg34 ?
                      (wire12 == reg35) : $signed((8'hac))) : $unsigned($signed(forvar32)))),
              wire7})
            begin
              reg36 <= (~$signed($unsigned(reg20[(1'h1):(1'h1)])));
              reg37 <= wire11[(2'h3):(2'h2)];
            end
          else
            begin
              reg35 = {((-$unsigned(reg37)) ?
                      {$signed($unsigned((8'ha5)))} : (((reg14 ?
                                  (8'had) : reg33) ?
                              (reg33 ? (8'ha9) : wire7) : {wire11}) ?
                          ((~|reg15) ?
                              (~&wire11) : $unsigned((8'hbd))) : ((wire7 ?
                                  forvar13 : reg24) ?
                              (^(8'hae)) : $signed((8'ha2))))),
                  (+(($signed(reg30) ?
                      $signed((7'h40)) : (wire10 + reg19)) > (reg34[(1'h0):(1'h0)] != (reg23 ?
                      reg36 : (8'hbe)))))};
            end
          if ($unsigned($signed({$signed((reg18 ? (7'h44) : wire7)), reg17})))
            begin
              reg38 <= wire9[(1'h0):(1'h0)];
              reg39 = ($unsigned(((8'hb0) == $unsigned({reg31, wire12}))) ?
                  (($unsigned(reg28) > reg14) ^~ ((reg19[(4'h8):(2'h3)] ^~ (wire10 << wire7)) ?
                      $unsigned((reg23 ? reg35 : reg14)) : reg23)) : wire7);
              reg40 <= (8'h9e);
              reg41 <= (+($unsigned($unsigned(wire7)) ?
                  $unsigned((~|(reg35 <= reg17))) : (~^(-((8'hb4) ?
                      reg22 : wire8)))));
              reg42 = ((|((&(^~reg39)) ?
                      wire11 : $unsigned($unsigned(wire12)))) ?
                  $signed((wire8[(1'h1):(1'h1)] ?
                      (+{wire11,
                          reg20}) : (~|(wire11 & reg39)))) : ($unsigned({$signed((8'h9c)),
                      ((8'hac) * reg30)}) && $signed(({wire11} && (reg35 ?
                      reg28 : reg31)))));
            end
          else
            begin
              reg38 <= (~|$signed((wire8[(3'h7):(3'h5)] ?
                  ($unsigned(reg40) <= $signed(reg29)) : ({reg20,
                      reg41} | reg27))));
              reg39 = $signed((8'hb7));
            end
        end
      if ((({((^reg36) ?
              wire12[(1'h0):(1'h0)] : (reg26 ?
                  reg16 : wire10))} || ($unsigned(reg20) ?
          ((^~reg33) == ((8'hb9) <<< reg18)) : ($signed(reg20) != $unsigned(reg42)))) ^~ (-$signed(reg23))))
        begin
          if ($signed(($unsigned(($unsigned(wire10) ?
              (8'had) : (reg23 || wire9))) & reg19)))
            begin
              reg43 <= (reg41 & wire11[(3'h4):(2'h3)]);
            end
          else
            begin
              reg43 <= $unsigned($unsigned({$unsigned($unsigned((8'ha6))),
                  reg30[(1'h1):(1'h1)]}));
              reg44 <= $signed(reg35[(4'h8):(3'h6)]);
              reg45 <= reg39;
              reg46 = reg38[(4'hb):(4'ha)];
            end
          if ((wire8 << (reg41 + ((~(reg16 ? (8'haa) : reg37)) ?
              ((reg39 - reg18) >>> reg18[(4'h8):(3'h7)]) : wire10))))
            begin
              reg47 <= $signed((8'hb4));
            end
          else
            begin
              reg47 <= (($unsigned($unsigned((reg32 == reg20))) ?
                      {(reg34[(3'h5):(1'h0)] ?
                              reg30[(3'h6):(1'h1)] : $unsigned(forvar13)),
                          {$unsigned(reg18)}} : reg31[(1'h1):(1'h0)]) ?
                  reg25[(2'h2):(1'h1)] : $unsigned((^~((~|(8'hac)) ?
                      (wire11 == reg47) : $signed(reg35)))));
              reg48 <= $unsigned((~({{reg35}} ?
                  ((!reg30) ? (reg44 >> wire6) : (reg29 + reg17)) : ((-reg15) ?
                      $unsigned(wire12) : $unsigned(wire8)))));
              reg49 = reg30;
            end
          if ({((wire12[(4'h9):(3'h5)] ?
                  wire6[(4'hb):(4'hb)] : reg16[(2'h3):(1'h0)]) >= (forvar32 != reg16)),
              $signed((-(reg35 && reg44)))})
            begin
              reg50 <= ((!(8'hb9)) ? reg34[(4'hd):(3'h5)] : (8'hb3));
              reg51 = $unsigned(((~|($signed(reg29) - $unsigned(reg24))) ?
                  $unsigned(forvar13) : reg38));
              reg52 = reg36;
              reg53 = reg14;
              reg54 <= ($unsigned((~&(8'h9e))) ?
                  reg17 : $unsigned($unsigned(($unsigned(reg46) ^ (reg51 - reg17)))));
            end
          else
            begin
              reg51 = ($signed({(reg16 >= ((8'hbc) && (8'ha4))),
                  $unsigned(reg31)}) * reg31);
            end
          if ((($signed(($signed(reg52) + $signed(wire8))) <<< (8'h9f)) | ((!((reg41 ?
                  reg48 : (8'h9e)) ?
              (reg30 ? reg47 : reg49) : ((8'hb8) ?
                  (8'hbf) : reg44))) << $unsigned(reg33))))
            begin
              reg55 <= (reg53[(2'h2):(2'h2)] ?
                  {{reg36[(3'h4):(1'h0)]}} : ({$unsigned((~&wire7))} ?
                      $unsigned({(~&wire11)}) : {reg35[(4'hb):(4'hb)]}));
            end
          else
            begin
              reg55 <= ((reg26 <<< $unsigned((wire6[(2'h3):(1'h1)] >= (wire8 ?
                      reg33 : (8'hb6))))) ?
                  reg39[(4'h9):(1'h0)] : reg33[(3'h5):(3'h5)]);
            end
          for (forvar56 = (1'h0); (forvar56 < (2'h2)); forvar56 = (forvar56 + (1'h1)))
            begin
              reg57 = reg30[(1'h0):(1'h0)];
              reg58 <= reg44;
              reg59 <= (-$unsigned(reg37));
              reg60 <= (8'hb2);
            end
        end
      else
        begin
          for (forvar43 = (1'h0); (forvar43 < (2'h2)); forvar43 = (forvar43 + (1'h1)))
            begin
              reg46 = reg51[(4'h8):(4'h8)];
              reg47 <= (^~(($signed((reg41 >= forvar32)) < ($signed(forvar43) ?
                      reg50 : $unsigned(reg52))) ?
                  (~|(&$unsigned(reg52))) : ($unsigned((~^(8'hbe))) & (reg30[(4'h8):(2'h3)] || wire7[(4'hb):(4'h8)]))));
              reg49 = ($signed(($unsigned($signed(reg49)) ?
                  ((-reg37) >> {reg36}) : ((&reg46) <<< (reg30 <<< reg44)))) && wire11[(4'hd):(4'hc)]);
              reg51 = ($signed($unsigned({(reg52 ? (8'hb9) : reg46)})) ?
                  (forvar32 ?
                      (~reg36) : $signed(((reg46 ?
                          reg29 : reg40) <= $signed(reg53)))) : reg54[(4'h8):(1'h0)]);
            end
        end
    end
  assign wire61 = $signed((wire9 <<< $signed(reg58)));
  assign wire62 = $signed(reg43);
  assign wire63 = ($signed((reg25 ?
                      reg36 : $signed(reg18[(4'hb):(4'h8)]))) ^~ reg59[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg64 = reg20;
      reg65 <= (&$signed($signed($signed((reg20 ^~ reg44)))));
      for (forvar66 = (1'h0); (forvar66 < (3'h4)); forvar66 = (forvar66 + (1'h1)))
        begin
          if ($signed($signed(({wire7, $unsigned(reg18)} ?
              ($unsigned(reg16) < (^~reg60)) : reg43))))
            begin
              reg67 <= $unsigned($signed((((reg55 * reg29) | (reg45 ?
                  (8'ha1) : reg45)) < (reg17[(1'h1):(1'h1)] ?
                  (forvar66 ? wire61 : wire62) : (~|reg16)))));
              reg68 <= ($signed((~&reg41)) + reg27[(3'h5):(3'h4)]);
              reg69 = ($signed(reg33) & ((($unsigned(wire12) << reg64[(5'h13):(3'h6)]) >> {{reg47,
                      reg45}}) >> (reg18[(4'he):(2'h3)] ?
                  reg29[(2'h2):(2'h2)] : $unsigned($unsigned(reg18)))));
              reg70 = $signed(reg40);
              reg71 = (+($unsigned(reg48[(3'h4):(2'h3)]) >>> (~&({(8'hab)} ?
                  $unsigned(wire63) : reg38))));
            end
          else
            begin
              reg67 <= $unsigned($unsigned(reg60));
              reg69 = (+({($signed(wire7) - ((8'h9e) && reg47))} ?
                  $signed(((reg41 >> reg70) - (^(8'ha7)))) : (!(~|$unsigned(wire10)))));
            end
          if ($unsigned((reg23[(4'h9):(3'h5)] ? $unsigned(wire63) : reg37)))
            begin
              reg72 <= $signed((($unsigned(reg28) >= ((!wire8) ?
                      $unsigned(reg67) : (reg58 ~^ reg55))) ?
                  $unsigned($signed((forvar66 != reg45))) : reg33[(3'h5):(2'h2)]));
              reg73 <= wire61;
              reg74 <= ((^reg20[(1'h0):(1'h0)]) <= (+reg21[(4'hd):(3'h6)]));
              reg75 = (($unsigned(($unsigned(reg33) < $unsigned((8'hb4)))) || reg30[(3'h6):(3'h5)]) ?
                  $signed($unsigned($signed((&reg36)))) : $unsigned((~^reg34)));
              reg76 = ($signed({(forvar66[(3'h5):(2'h3)] - reg65)}) < wire12);
            end
          else
            begin
              reg75 = (8'hbd);
              reg76 = (~(reg45 ?
                  ((~&reg41[(1'h0):(1'h0)]) ?
                      reg73 : $unsigned(reg44)) : (((^reg59) ?
                      ((7'h41) + reg36) : (reg38 ^~ reg50)) >= (reg67[(2'h3):(1'h0)] ?
                      (!(8'hac)) : (~|reg71)))));
              reg77 = {{$unsigned((+wire11))}};
              reg78 <= $signed($signed((($unsigned(reg28) ?
                      (wire9 ? wire61 : reg40) : $signed((8'h9f))) ?
                  ((reg44 < reg74) ?
                      reg16[(1'h0):(1'h0)] : (&(8'ha4))) : $unsigned(((8'hab) ?
                      reg41 : reg71)))));
              reg79 <= $unsigned((reg72 ?
                  forvar66 : $unsigned((&((8'hbf) >> wire6)))));
            end
          reg80 = (((((wire61 ? wire63 : reg38) || reg43) ?
                  ((reg78 || reg43) < $unsigned(reg64)) : $unsigned(reg60[(4'hd):(4'hc)])) ?
              (reg70[(3'h6):(1'h0)] != (-(reg28 | reg59))) : reg50) ~^ $unsigned($signed({(reg72 ?
                  (8'hb8) : wire8)})));
          if (((7'h41) ^~ $unsigned(($unsigned($unsigned(wire10)) ?
              $signed(reg60) : $unsigned($unsigned(reg33))))))
            begin
              reg81 <= reg79[(3'h7):(3'h7)];
              reg82 <= reg80[(1'h0):(1'h0)];
              reg83 <= $unsigned(reg30);
              reg84 <= wire10[(4'hd):(2'h2)];
            end
          else
            begin
              reg81 <= $signed((&wire63));
              reg85 = ((8'ha1) ?
                  ($unsigned(($unsigned((8'haa)) ?
                          (!(8'ha6)) : $signed(reg23))) ?
                      ((|(~|reg81)) ?
                          ((reg67 >= reg15) ?
                              {reg33} : (reg84 != (8'haf))) : $signed((reg20 ?
                              (8'ha1) : (8'hab)))) : ({(reg73 >> reg70),
                              reg77} ?
                          reg68[(2'h2):(2'h2)] : (-(reg30 ^~ reg48)))) : {(~^$signed({reg16,
                          (8'hb9)})),
                      (wire12 ? (^~(reg73 << wire8)) : reg30)});
              reg86 <= $signed((^~(reg43 ?
                  {{(8'hbe), reg75},
                      reg70[(3'h6):(3'h5)]} : (((8'hbe) << reg20) * $signed(reg40)))));
              reg87 = $signed((+({$signed(reg70), (~&(8'hbc))} ?
                  $signed({reg15}) : wire9[(2'h2):(2'h2)])));
              reg88 = (8'ha4);
            end
          reg89 <= $signed(($signed(wire6) <= (8'hb1)));
        end
      for (forvar90 = (1'h0); (forvar90 < (1'h1)); forvar90 = (forvar90 + (1'h1)))
        begin
          if ((-(-(((8'ha4) == $signed(wire10)) ?
              reg34 : $signed((reg81 - reg80))))))
            begin
              reg91 = $signed($unsigned($unsigned(reg45)));
              reg92 <= (^~$unsigned($unsigned((|(wire8 == reg72)))));
              reg93 <= reg17[(3'h4):(2'h2)];
              reg94 <= $signed((8'h9e));
            end
          else
            begin
              reg92 <= $signed(($unsigned((~&$unsigned(reg58))) ?
                  (~|((~&wire61) ?
                      reg70[(3'h6):(2'h2)] : $signed(wire8))) : ($signed((~&(8'ha8))) ?
                      reg41 : (|$signed((8'hbc))))));
              reg93 <= $signed((reg44[(4'h9):(3'h7)] ?
                  wire7[(2'h2):(1'h1)] : {reg30}));
              reg95 = {(!$unsigned(reg92[(1'h0):(1'h0)]))};
              reg96 <= (^reg65);
              reg97 = $signed(reg34);
            end
          for (forvar98 = (1'h0); (forvar98 < (2'h2)); forvar98 = (forvar98 + (1'h1)))
            begin
              reg99 <= reg80;
              reg100 = (((~|reg20) ^ reg77[(1'h0):(1'h0)]) ~^ (~|$unsigned((reg92[(1'h0):(1'h0)] ?
                  ((8'ha6) || reg95) : $unsigned(reg55)))));
              reg101 = {reg71, reg74};
            end
          reg102 = (!((&(((8'hb1) ? reg88 : reg77) ?
                  $signed(wire12) : ((8'hb9) || wire9))) ?
              reg67 : $signed(($signed(reg45) ^ (&(8'hb7))))));
          reg103 <= ((8'ha4) ?
              reg41 : (($unsigned(reg21) ?
                  {(reg102 ? reg60 : reg94),
                      $unsigned(reg82)} : $signed(reg68)) + ($unsigned(reg87[(2'h3):(2'h2)]) ?
                  reg37[(3'h6):(2'h3)] : (reg44[(2'h2):(1'h0)] <<< reg44))));
        end
    end
  always
    @(posedge clk) begin
      reg104 = $signed($signed(reg92));
      for (forvar105 = (1'h0); (forvar105 < (1'h1)); forvar105 = (forvar105 + (1'h1)))
        begin
          reg106 = $unsigned({wire61[(3'h5):(3'h5)]});
        end
      if ((~|((7'h42) | $unsigned($signed($signed(reg86))))))
        begin
          reg107 = (reg45[(4'h9):(3'h4)] ~^ (reg45 ?
              ($signed($unsigned(reg48)) ?
                  {$signed(reg44)} : ((8'hba) ?
                      reg58[(5'h11):(4'hc)] : $unsigned((7'h44)))) : {{(wire8 * reg43),
                      $signed(reg21)}}));
        end
      else
        begin
          if ($unsigned($unsigned(reg94)))
            begin
              reg108 <= wire12;
              reg109 = ($unsigned((|$signed($signed((8'hbe))))) <= (~(($unsigned(wire8) > reg34[(2'h3):(2'h3)]) + reg89[(2'h3):(2'h3)])));
              reg110 = $signed(reg82[(1'h0):(1'h0)]);
            end
          else
            begin
              reg108 <= (^$signed($unsigned((|(reg55 ? (8'hb3) : reg104)))));
              reg111 <= (8'hb4);
            end
          if ($unsigned(reg83[(3'h7):(3'h6)]))
            begin
              reg112 <= (reg50[(3'h5):(2'h2)] ?
                  reg103[(4'hc):(1'h0)] : reg27[(1'h0):(1'h0)]);
              reg113 = (-reg50[(4'h8):(2'h3)]);
            end
          else
            begin
              reg113 = (reg108 ?
                  (reg23[(5'h13):(4'hb)] ?
                      (reg79 >= $unsigned((+reg34))) : ($signed({reg17}) ?
                          $signed($unsigned(reg23)) : wire62)) : {(!$signed(((8'hab) ?
                          reg111 : reg93))),
                      $unsigned($signed((reg45 ? reg15 : reg21)))});
              reg114 <= $unsigned(reg79);
              reg115 <= $unsigned($unsigned(reg55[(1'h0):(1'h0)]));
              reg116 <= $unsigned((((8'hba) < {$unsigned(reg21)}) <<< $signed(reg113[(2'h3):(2'h2)])));
            end
        end
    end
  assign wire117 = $unsigned(reg37);
  assign wire118 = (~^reg17[(3'h6):(2'h3)]);
  module119 #() modinst314 (wire313, clk, wire9, reg116, wire10, wire8, reg73);
  assign wire315 = reg73[(3'h4):(1'h1)];
  module316 #() modinst558 (wire557, clk, wire8, reg72, reg74, reg73);
  assign wire559 = (!({reg50[(2'h2):(1'h0)], $signed((+reg116))} ?
                       $unsigned({wire8[(4'h9):(3'h5)],
                           (8'h9c)}) : $signed($unsigned({wire313, reg73}))));
  module560 #() modinst699 (.wire561(reg68), .wire564(reg41), .y(wire698), .clk(clk), .wire563(reg18), .wire562(wire6));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module560
#(parameter param696 = ((({(^~(8'hac))} ? (~|((8'ha0) - (7'h44))) : {((8'ha9) ? (8'hb1) : (8'ha3))}) <= ((((8'hbc) ? (8'hb0) : (8'hb6)) ? (^~(8'h9f)) : (~|(8'ha2))) ? ((8'hbf) ? {(8'hbf)} : ((8'hba) ? (8'ha9) : (8'hb0))) : (~&{(8'hbd)}))) ? ((((^~(8'ha0)) - ((8'ha1) ? (8'hb7) : (8'hba))) * (((8'hb6) ? (8'hb5) : (8'ha4)) ? ((8'ha2) ? (8'ha2) : (8'ha4)) : ((8'hbe) == (8'ha6)))) ? (((^(7'h40)) ? ((8'hb1) ? (8'h9e) : (8'ha0)) : (8'hb4)) ^~ (((8'hbf) << (8'hbe)) == (^~(8'hb3)))) : (+((~&(8'hab)) ? (~^(8'hb1)) : (8'hb0)))) : (((~&((7'h43) * (8'hac))) && {(-(8'ha2)), {(7'h40)}}) == (&(8'hb3)))), 
parameter param697 = (~^((^(~{(8'hb0)})) ? ((param696 ? {param696, param696} : (8'ha3)) ? {(|(8'ha0)), param696} : param696) : param696)))
(y, clk, wire564, wire563, wire562, wire561);
  output wire [(32'h647):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire564;
  input wire signed [(4'h9):(1'h0)] wire563;
  input wire signed [(5'h10):(1'h0)] wire562;
  input wire signed [(3'h4):(1'h0)] wire561;
  wire signed [(4'h9):(1'h0)] wire674;
  wire signed [(4'h8):(1'h0)] wire673;
  wire [(5'h15):(1'h0)] wire672;
  wire signed [(4'h8):(1'h0)] wire572;
  wire [(3'h4):(1'h0)] wire571;
  wire signed [(5'h12):(1'h0)] wire570;
  wire signed [(2'h2):(1'h0)] wire569;
  wire signed [(4'h8):(1'h0)] wire568;
  wire signed [(5'h13):(1'h0)] wire567;
  wire signed [(5'h15):(1'h0)] wire566;
  wire signed [(4'he):(1'h0)] wire565;
  reg signed [(2'h3):(1'h0)] reg694 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg692 = (1'h0);
  reg [(4'hb):(1'h0)] reg690 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg689 = (1'h0);
  reg [(4'hb):(1'h0)] reg676 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg688 = (1'h0);
  reg [(3'h7):(1'h0)] reg686 = (1'h0);
  reg [(4'h9):(1'h0)] reg684 = (1'h0);
  reg [(4'h9):(1'h0)] reg683 = (1'h0);
  reg [(4'hd):(1'h0)] reg681 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg680 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg679 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg677 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg675 = (1'h0);
  reg [(4'hd):(1'h0)] reg671 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg669 = (1'h0);
  reg [(4'he):(1'h0)] reg668 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg666 = (1'h0);
  reg [(3'h4):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg660 = (1'h0);
  reg [(4'hf):(1'h0)] reg658 = (1'h0);
  reg [(4'h8):(1'h0)] reg657 = (1'h0);
  reg signed [(4'he):(1'h0)] reg655 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg652 = (1'h0);
  reg [(2'h3):(1'h0)] reg651 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg650 = (1'h0);
  reg signed [(4'he):(1'h0)] reg649 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg648 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg647 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg645 = (1'h0);
  reg signed [(4'he):(1'h0)] reg644 = (1'h0);
  reg [(3'h7):(1'h0)] reg642 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg643 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg635 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg634 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg633 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg631 = (1'h0);
  reg [(3'h6):(1'h0)] reg630 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg626 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg625 = (1'h0);
  reg [(5'h15):(1'h0)] reg624 = (1'h0);
  reg [(4'hf):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg622 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg621 = (1'h0);
  reg [(5'h11):(1'h0)] reg620 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg618 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg617 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg611 = (1'h0);
  reg [(4'ha):(1'h0)] reg608 = (1'h0);
  reg [(4'h9):(1'h0)] reg607 = (1'h0);
  reg [(4'h8):(1'h0)] reg606 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg605 = (1'h0);
  reg [(5'h11):(1'h0)] reg604 = (1'h0);
  reg [(3'h6):(1'h0)] reg603 = (1'h0);
  reg [(4'h9):(1'h0)] reg599 = (1'h0);
  reg [(3'h7):(1'h0)] reg597 = (1'h0);
  reg [(4'h9):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg593 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg590 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg589 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg588 = (1'h0);
  reg [(3'h6):(1'h0)] reg587 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg585 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg584 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg582 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg581 = (1'h0);
  reg [(4'he):(1'h0)] reg580 = (1'h0);
  reg [(4'hb):(1'h0)] reg578 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg577 = (1'h0);
  reg [(4'h9):(1'h0)] reg575 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg695 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg693 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar691 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar684 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg687 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg685 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg682 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg678 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar676 = (1'h0);
  reg [(4'hf):(1'h0)] reg670 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg663 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg662 = (1'h0);
  reg [(5'h14):(1'h0)] forvar659 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar653 = (1'h0);
  reg [(3'h6):(1'h0)] reg656 = (1'h0);
  reg [(2'h2):(1'h0)] reg654 = (1'h0);
  reg [(4'hc):(1'h0)] reg653 = (1'h0);
  reg [(5'h11):(1'h0)] reg646 = (1'h0);
  reg [(4'hc):(1'h0)] forvar642 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg641 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg640 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg639 = (1'h0);
  reg [(4'h8):(1'h0)] reg638 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg637 = (1'h0);
  reg [(2'h2):(1'h0)] reg636 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg629 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar622 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg627 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg619 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg616 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg615 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar614 = (1'h0);
  reg [(3'h4):(1'h0)] reg613 = (1'h0);
  reg [(4'hc):(1'h0)] reg610 = (1'h0);
  reg [(5'h14):(1'h0)] reg609 = (1'h0);
  reg [(5'h13):(1'h0)] reg602 = (1'h0);
  reg [(4'ha):(1'h0)] reg601 = (1'h0);
  reg [(4'hc):(1'h0)] reg600 = (1'h0);
  reg [(5'h15):(1'h0)] reg598 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg594 = (1'h0);
  reg [(5'h15):(1'h0)] reg592 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg591 = (1'h0);
  reg [(3'h6):(1'h0)] reg586 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg583 = (1'h0);
  reg [(4'h8):(1'h0)] reg579 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg576 = (1'h0);
  reg [(5'h11):(1'h0)] forvar573 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar576 = (1'h0);
  reg [(3'h7):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg573 = (1'h0);
  assign y = {wire674,
                 wire673,
                 wire672,
                 wire572,
                 wire571,
                 wire570,
                 wire569,
                 wire568,
                 wire567,
                 wire566,
                 wire565,
                 reg694,
                 reg692,
                 reg690,
                 reg689,
                 reg676,
                 reg688,
                 reg686,
                 reg684,
                 reg683,
                 reg681,
                 reg680,
                 reg679,
                 reg677,
                 reg675,
                 reg671,
                 reg669,
                 reg668,
                 reg666,
                 reg665,
                 reg664,
                 reg661,
                 reg660,
                 reg658,
                 reg657,
                 reg655,
                 reg652,
                 reg651,
                 reg650,
                 reg649,
                 reg648,
                 reg647,
                 reg645,
                 reg644,
                 reg642,
                 reg643,
                 reg635,
                 reg634,
                 reg633,
                 reg631,
                 reg630,
                 reg628,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 reg618,
                 reg617,
                 reg612,
                 reg611,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg599,
                 reg597,
                 reg596,
                 reg595,
                 reg593,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg585,
                 reg584,
                 reg582,
                 reg581,
                 reg580,
                 reg578,
                 reg577,
                 reg575,
                 reg695,
                 reg693,
                 forvar691,
                 forvar684,
                 reg687,
                 reg685,
                 reg682,
                 reg678,
                 forvar676,
                 reg670,
                 reg667,
                 reg663,
                 reg662,
                 forvar659,
                 forvar653,
                 reg656,
                 reg654,
                 reg653,
                 reg646,
                 forvar642,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 reg632,
                 reg629,
                 forvar622,
                 reg627,
                 reg619,
                 reg616,
                 reg615,
                 forvar614,
                 reg613,
                 reg610,
                 reg609,
                 reg602,
                 reg601,
                 reg600,
                 reg598,
                 reg594,
                 reg592,
                 reg591,
                 reg586,
                 reg583,
                 reg579,
                 reg576,
                 forvar573,
                 forvar576,
                 reg574,
                 reg573,
                 (1'h0)};
  assign wire565 = (&(((~&(wire564 ? wire563 : wire561)) && $unsigned((wire564 ?
                       wire564 : wire564))) != wire564[(2'h3):(1'h1)]));
  assign wire566 = {wire565};
  assign wire567 = (-wire562);
  assign wire568 = {$signed(($signed($unsigned(wire562)) ?
                           (~&(&wire561)) : $signed($unsigned(wire565))))};
  assign wire569 = wire561[(2'h3):(2'h2)];
  assign wire570 = $signed((&($unsigned($signed(wire568)) ?
                       ((^wire561) ~^ (wire562 ~^ wire567)) : (^$signed((8'hab))))));
  assign wire571 = $signed(wire564[(4'h9):(3'h4)]);
  assign wire572 = {{(-(^$signed(wire563)))},
                       ((({wire567} ? (~|wire566) : (8'hb2)) && wire564) ?
                           (-$signed((wire571 ?
                               wire568 : wire568))) : $signed($unsigned((~wire562))))};
  always
    @(posedge clk) begin
      if (({$signed((wire565[(3'h4):(1'h0)] ?
                  $unsigned(wire570) : (^~wire571)))} ?
          (-wire572[(3'h6):(3'h4)]) : (7'h42)))
        begin
          if (wire572)
            begin
              reg573 = (|(((wire566 ?
                      ((8'hbd) ?
                          wire568 : wire570) : wire565) ^ (~(wire561 == wire561))) ?
                  ($signed(wire566[(4'he):(1'h0)]) + $signed((wire564 ?
                      wire568 : wire567))) : (($unsigned((8'ha2)) ?
                          wire569[(1'h1):(1'h0)] : $signed((8'ha3))) ?
                      wire570 : wire566)));
              reg574 = ((+$unsigned(((wire568 >= (8'ha4)) + $signed((7'h41))))) <= wire562[(4'h8):(3'h4)]);
            end
          else
            begin
              reg573 = ((~wire569) ^~ (~wire569[(1'h1):(1'h0)]));
              reg575 <= ((((+(wire570 * wire572)) ?
                  (+$signed(wire571)) : ((reg573 ?
                      wire562 : wire570) >>> wire561)) != $signed(((wire563 ?
                      (7'h44) : wire571) ?
                  wire563 : $unsigned(wire569)))) >>> ($unsigned((+wire565[(4'h9):(3'h7)])) ?
                  wire563[(4'h9):(1'h1)] : wire565));
            end
          for (forvar576 = (1'h0); (forvar576 < (2'h3)); forvar576 = (forvar576 + (1'h1)))
            begin
              reg577 <= (~|((-$signed((wire561 << wire570))) >>> $signed(wire563)));
            end
        end
      else
        begin
          for (forvar573 = (1'h0); (forvar573 < (2'h3)); forvar573 = (forvar573 + (1'h1)))
            begin
              reg575 <= $signed({(~^reg574)});
              reg576 = forvar576[(1'h1):(1'h0)];
              reg577 <= $unsigned(((!wire564[(1'h0):(1'h0)]) ^~ ((forvar573 ?
                  {wire564} : ((8'ha9) >= wire561)) >> (!{wire570, wire570}))));
              reg578 <= $signed(wire564[(3'h5):(1'h0)]);
            end
          if ((!(((^~{reg576, reg574}) ?
              $unsigned((!(8'ha1))) : {wire562,
                  $signed(wire572)}) << ($unsigned(wire569) & ($unsigned(wire561) ^~ $unsigned(wire572))))))
            begin
              reg579 = $signed(($signed($signed(wire567[(1'h1):(1'h1)])) ?
                  ((~^forvar573[(1'h0):(1'h0)]) - wire561[(2'h3):(1'h0)]) : (((wire570 ?
                      forvar576 : reg574) <= reg575) || $signed($signed(wire561)))));
              reg580 <= $unsigned(reg577);
              reg581 <= (((~&$signed($signed((7'h44)))) ?
                  (reg578[(3'h6):(3'h6)] ?
                      $unsigned((~^wire570)) : {(8'hb7),
                          $signed(wire564)}) : (wire565[(3'h6):(1'h0)] ^~ ($unsigned(forvar576) >= $signed(wire561)))) == (reg574[(3'h4):(2'h2)] ?
                  ($unsigned({wire568}) ?
                      ((|wire563) ?
                          $unsigned(reg573) : (reg577 >>> reg576)) : $signed($signed(wire569))) : ((|(wire561 ~^ (8'hb7))) || (^~(reg580 ?
                      (8'ha1) : reg580)))));
            end
          else
            begin
              reg580 <= $unsigned((|(&$signed(forvar576[(2'h3):(1'h0)]))));
              reg581 <= {($signed(reg576[(4'hc):(4'hb)]) ^ ($signed((wire563 * wire562)) << reg576))};
              reg582 <= (!(($unsigned(wire567[(4'hd):(2'h2)]) + {reg580,
                      (forvar573 ? wire565 : (8'ha8))}) ?
                  $unsigned({$unsigned(wire565),
                      (forvar576 >= wire565)}) : reg581));
              reg583 = (&($unsigned(($unsigned((7'h44)) == (wire567 ?
                  wire565 : (7'h42)))) > {(8'hbb), {(^wire566)}}));
              reg584 <= {$unsigned(reg576), wire570};
            end
          if ($unsigned((8'hbc)))
            begin
              reg585 <= $unsigned($signed($unsigned(wire569[(1'h1):(1'h0)])));
              reg586 = wire562;
              reg587 <= (~|(reg586 == (~|(reg577 ?
                  $signed(reg579) : wire569[(2'h2):(2'h2)]))));
              reg588 <= $unsigned((($unsigned(reg575) >>> reg584) ?
                  $unsigned(reg580[(4'h8):(4'h8)]) : reg585[(1'h0):(1'h0)]));
            end
          else
            begin
              reg586 = (({wire565[(3'h5):(1'h0)]} ?
                  reg581[(3'h6):(3'h5)] : (^(((8'h9c) || reg580) - reg580[(4'hd):(4'ha)]))) << (^~wire566[(1'h1):(1'h1)]));
              reg587 <= $unsigned((wire564 <<< (&(~|$signed(reg588)))));
              reg588 <= reg584;
              reg589 <= wire572[(3'h6):(1'h1)];
              reg590 <= $signed(wire572);
            end
        end
      if ($signed((-(~|wire565))))
        begin
          reg591 = (|(!reg578[(4'h8):(2'h2)]));
          if (reg581)
            begin
              reg592 = wire568;
            end
          else
            begin
              reg592 = $unsigned($signed({wire564[(2'h3):(2'h2)]}));
              reg593 <= $unsigned(reg580);
              reg594 = {$unsigned(wire570),
                  (($unsigned((reg585 ? wire563 : reg575)) >>> {(reg578 ?
                          wire572 : wire571),
                      (&wire563)}) ~^ ((^$signed(reg588)) ?
                      (!(wire572 - reg580)) : (~&reg589)))};
              reg595 <= reg588[(3'h4):(3'h4)];
              reg596 <= reg589[(4'h8):(3'h7)];
            end
          if (reg583[(4'hc):(3'h5)])
            begin
              reg597 <= reg587[(3'h5):(1'h1)];
              reg598 = $unsigned($signed(({$unsigned(reg576)} > (~(reg580 ?
                  reg576 : reg578)))));
              reg599 <= $signed(reg580);
            end
          else
            begin
              reg597 <= reg584[(3'h6):(3'h4)];
              reg599 <= reg597[(3'h6):(3'h6)];
              reg600 = {wire564};
            end
          if ($unsigned($unsigned((~&wire568))))
            begin
              reg601 = {wire566[(2'h2):(1'h1)],
                  $signed({wire569,
                      ($signed(reg595) ?
                          wire572[(1'h1):(1'h0)] : ((8'haf) ?
                              reg582 : reg597))})};
              reg602 = ($signed(reg584) << ((reg578[(2'h3):(1'h1)] ?
                      reg577[(1'h0):(1'h0)] : (8'hab)) ?
                  ($signed($signed(reg598)) ?
                      $unsigned((reg586 << wire570)) : (&(wire564 ?
                          reg579 : reg589))) : reg588[(3'h4):(1'h1)]));
            end
          else
            begin
              reg603 <= wire570;
              reg604 <= (reg601[(3'h6):(2'h2)] < (~|$signed(($signed(reg577) ?
                  (^~reg585) : $signed(reg590)))));
              reg605 <= $signed($unsigned(reg592[(2'h2):(1'h1)]));
              reg606 <= reg583;
            end
          if ((~|(wire563[(4'h9):(3'h6)] ^ $signed($unsigned((~|reg577))))))
            begin
              reg607 <= $signed((reg582 ?
                  {(~(~|reg573)),
                      ({reg583} ?
                          reg593[(1'h0):(1'h0)] : wire568[(1'h1):(1'h0)])} : reg579));
              reg608 <= (-$unsigned(forvar576[(1'h0):(1'h0)]));
            end
          else
            begin
              reg609 = (reg579[(1'h1):(1'h0)] ^~ reg585);
              reg610 = (((~&$signed({reg601})) >>> $signed($unsigned((&reg579)))) == (~^reg574));
              reg611 <= reg580[(3'h6):(3'h4)];
              reg612 <= ((reg607[(3'h4):(3'h4)] + (~&$signed((reg585 << reg611)))) ?
                  wire561[(2'h3):(1'h0)] : {$signed(reg600[(1'h0):(1'h0)])});
            end
        end
      else
        begin
          reg593 <= (-{(reg608[(3'h4):(1'h0)] <<< $signed(reg607[(4'h9):(2'h3)])),
              $unsigned((reg601 || ((8'ha8) ? wire563 : forvar576)))});
          if ((~&$signed(reg585[(1'h0):(1'h0)])))
            begin
              reg594 = $unsigned(($signed(reg592[(4'ha):(4'h9)]) ?
                  wire565 : $unsigned((-(-reg589)))));
              reg595 <= ((+reg576) ?
                  reg580[(4'hd):(1'h0)] : $unsigned(({$signed(wire564)} ?
                      (~wire569) : {(~^reg592), (+wire564)})));
            end
          else
            begin
              reg594 = (reg585 >> (((~reg607) || ((reg575 ? reg610 : reg593) ?
                  $signed(reg596) : $signed(reg579))) && ((reg610[(3'h5):(1'h1)] ?
                  (wire569 <= reg607) : $unsigned(wire571)) << {(reg599 ?
                      reg597 : reg593),
                  reg603})));
              reg598 = reg585[(1'h1):(1'h1)];
              reg600 = reg580[(2'h3):(2'h2)];
              reg603 <= $signed($unsigned((!$unsigned((reg596 ?
                  (8'hb2) : wire566)))));
              reg604 <= (~&$unsigned($signed(reg601)));
            end
          if ((8'hb8))
            begin
              reg605 <= $unsigned($unsigned(reg592));
              reg609 = $signed((8'hbd));
              reg611 <= ((((~^(+reg601)) != ($signed(reg598) != (wire566 ^ forvar573))) ?
                      $signed((^$signed(reg612))) : reg586[(3'h6):(3'h4)]) ?
                  reg574[(2'h3):(1'h1)] : $unsigned(reg586[(3'h5):(1'h1)]));
            end
          else
            begin
              reg609 = wire570[(4'hc):(3'h5)];
              reg611 <= wire563[(3'h7):(1'h0)];
              reg613 = reg610;
            end
          for (forvar614 = (1'h0); (forvar614 < (2'h2)); forvar614 = (forvar614 + (1'h1)))
            begin
              reg615 = reg589;
              reg616 = wire562[(2'h3):(2'h2)];
            end
        end
      if ((~|reg573[(3'h6):(3'h4)]))
        begin
          if (($unsigned(wire563) ?
              $unsigned((reg592 + {reg608[(1'h0):(1'h0)]})) : $signed((8'h9d))))
            begin
              reg617 <= $signed(((-(~reg584)) ?
                  $signed($signed(reg598)) : reg585[(2'h2):(1'h0)]));
              reg618 <= (8'hbc);
            end
          else
            begin
              reg617 <= (~reg609);
              reg619 = $signed(wire572[(3'h7):(2'h3)]);
            end
          reg620 <= forvar576;
          reg621 <= (-(reg601 >= (8'ha5)));
          if ($signed(reg598[(1'h1):(1'h1)]))
            begin
              reg622 <= (reg584 <<< reg608);
              reg623 <= ((reg596[(4'h8):(1'h1)] << reg585[(1'h1):(1'h0)]) ?
                  reg598 : (wire571 ? $signed((|$signed(wire567))) : reg587));
              reg624 <= $unsigned($signed((reg597 <= (((7'h43) ~^ (8'ha1)) ?
                  $signed((7'h43)) : (reg596 ? (8'hbc) : reg605)))));
              reg625 <= $signed((|$unsigned({(wire567 ^~ wire569)})));
              reg626 <= reg603[(3'h5):(3'h4)];
            end
          else
            begin
              reg622 <= $unsigned(reg624[(5'h14):(4'h9)]);
              reg623 <= reg600;
            end
          if ($unsigned((^~reg612[(4'h9):(3'h5)])))
            begin
              reg627 = reg584;
            end
          else
            begin
              reg628 <= ((~&(~^forvar573[(2'h3):(2'h2)])) ?
                  (^~{$unsigned($unsigned((8'had))),
                      (~reg594[(4'ha):(3'h7)])}) : (!reg589));
            end
        end
      else
        begin
          reg619 = ((~&wire564[(2'h2):(1'h0)]) < $signed($unsigned((-(reg574 == (8'hbb))))));
          if ($unsigned(((~^$unsigned((reg577 ^~ (8'hbc)))) ?
              {{(|(8'ha7))}, (~(8'hb6))} : (reg577 << ($unsigned(reg575) ?
                  (wire569 * reg586) : {reg591})))))
            begin
              reg620 <= ((({(wire568 ? wire567 : (7'h44)),
                      ((8'hb5) ~^ reg607)} != (wire565 ?
                      reg582[(4'hc):(3'h4)] : (8'ha4))) ?
                  reg621 : (&(~reg580[(1'h0):(1'h0)]))) << (~^((8'ha4) >> {((8'h9d) ?
                      wire567 : reg602)})));
              reg621 <= $signed((reg577[(1'h1):(1'h1)] ?
                  (^~$signed((reg591 - reg589))) : $unsigned($unsigned($unsigned(wire562)))));
            end
          else
            begin
              reg620 <= {$signed(reg587),
                  (reg611[(4'hb):(4'h9)] ?
                      ({(|reg617),
                          {reg602,
                              reg579}} >>> (reg622 != reg591[(4'ha):(4'ha)])) : wire572)};
            end
          for (forvar622 = (1'h0); (forvar622 < (2'h3)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 <= (&($unsigned(reg596[(4'h8):(3'h7)]) ?
                  (reg580[(1'h0):(1'h0)] >>> (reg599[(1'h1):(1'h0)] ?
                      {(7'h43), reg573} : (forvar573 ?
                          (8'had) : reg608))) : (8'ha7)));
              reg627 = (reg587[(3'h4):(1'h0)] >= reg588[(2'h3):(2'h2)]);
              reg628 <= $signed(wire562[(4'hd):(2'h3)]);
              reg629 = ((reg576 && $unsigned((wire572[(2'h3):(2'h2)] >= {wire569,
                      forvar576}))) ?
                  {($signed(reg599) ?
                          ((~reg623) ?
                              $unsigned(reg608) : reg580[(4'ha):(4'ha)]) : (8'h9f)),
                      (^$signed($signed(reg603)))} : (reg599 ?
                      reg583 : $signed((~|reg608[(2'h2):(1'h0)]))));
            end
          if (reg624)
            begin
              reg630 <= (^~$signed(reg619[(3'h5):(1'h1)]));
            end
          else
            begin
              reg630 <= $signed($signed(wire562));
              reg631 <= $unsigned(reg630);
              reg632 = $signed(wire562);
              reg633 <= reg592;
            end
          if (((reg576 || {$signed(reg575[(3'h6):(1'h1)])}) ?
              (8'hba) : ((+$unsigned((reg592 & reg582))) ?
                  ((reg579 <<< (^~reg609)) ?
                      reg627 : $signed($signed(reg581))) : $signed(((wire570 ?
                          reg602 : wire564) ?
                      (reg618 ? reg575 : reg581) : (|(8'ha9)))))))
            begin
              reg634 <= (wire563 ?
                  reg609[(4'ha):(3'h5)] : (-wire564[(1'h1):(1'h0)]));
              reg635 <= $signed((~^(&reg611[(3'h7):(1'h1)])));
            end
          else
            begin
              reg636 = {reg617,
                  (|{((8'hb3) > reg623[(4'he):(4'hd)]),
                      reg613[(2'h3):(1'h0)]})};
              reg637 = $unsigned(reg623[(3'h5):(2'h3)]);
              reg638 = (&(reg631[(4'h8):(2'h2)] ?
                  {((^reg587) >> (|reg633))} : reg588));
              reg639 = {$unsigned($signed((reg618[(1'h1):(1'h1)] <= forvar576))),
                  $signed(forvar573)};
              reg640 = ($unsigned((reg603 >= {$unsigned((7'h41))})) | ((((-reg622) ?
                          (reg586 ? (8'hbe) : reg631) : {reg599, forvar622}) ?
                      $unsigned(reg580) : ($unsigned(reg616) ?
                          $unsigned(reg575) : forvar576[(1'h0):(1'h0)])) ?
                  {reg607, reg586} : reg597[(2'h2):(1'h0)]));
            end
        end
      if (({$signed(wire569),
          (8'ha5)} & ($unsigned(reg621[(3'h6):(2'h2)]) ^~ ($signed($signed(wire561)) ?
          $signed(reg621) : reg606))))
        begin
          reg641 = reg626;
          for (forvar642 = (1'h0); (forvar642 < (1'h0)); forvar642 = (forvar642 + (1'h1)))
            begin
              reg643 <= reg619;
            end
        end
      else
        begin
          if ((((({forvar642} ?
                      {(8'hb0),
                          reg611} : $signed(reg625)) && (reg609[(4'ha):(3'h6)] ?
                      (reg610 + (8'hb9)) : reg591)) ?
                  (7'h43) : reg596) ?
              ($unsigned($unsigned($unsigned(reg602))) ?
                  (!{$unsigned(wire570),
                      reg626[(3'h4):(2'h3)]}) : $signed((8'hbd))) : $signed(($signed(reg579) ?
                  reg632[(3'h7):(1'h1)] : ((&reg605) << reg627[(1'h1):(1'h0)])))))
            begin
              reg642 <= (($signed({reg584[(1'h1):(1'h0)],
                  (reg582 ? reg574 : reg594)}) >> (~{(reg623 ?
                      reg610 : reg580)})) & reg573);
              reg643 <= reg633[(4'h8):(2'h3)];
              reg644 <= reg582[(3'h5):(3'h4)];
              reg645 <= ((~^$signed($unsigned((reg640 ? reg618 : reg581)))) ?
                  (8'hbd) : ($unsigned(($unsigned(reg577) ?
                      (wire571 ?
                          reg586 : (8'ha4)) : (-wire561))) >= (((reg632 - reg596) ?
                          (-reg587) : (reg594 ^ reg623)) ?
                      reg604 : $signed(reg584))));
            end
          else
            begin
              reg642 <= $signed(((reg591[(3'h5):(1'h1)] ?
                      ($unsigned(reg620) ?
                          $unsigned((8'h9d)) : ((8'hba) ?
                              reg637 : reg576)) : reg581) ?
                  (^~reg645) : reg634));
            end
          if ((^~$signed(forvar622[(5'h11):(3'h7)])))
            begin
              reg646 = {(|$unsigned($signed($signed(reg616)))),
                  reg640[(3'h6):(1'h0)]};
              reg647 <= (~&(8'h9e));
              reg648 <= (~^($unsigned($unsigned($unsigned(reg647))) ?
                  forvar642[(3'h7):(3'h4)] : $signed(({reg630, reg622} ?
                      (reg627 ? reg628 : reg611) : ((8'hbe) ?
                          reg620 : reg591)))));
              reg649 <= reg602[(1'h0):(1'h0)];
            end
          else
            begin
              reg647 <= (((-(forvar614 ? reg633 : reg619)) ?
                  $signed(({reg588,
                      wire568} ^~ reg617)) : $unsigned(($signed(reg592) ^~ (reg594 ?
                      (8'h9e) : reg610)))) && (~^reg630));
              reg648 <= reg638;
              reg649 <= (($unsigned((~^$unsigned((8'hb4)))) | {(~|{reg604})}) ?
                  $unsigned((((reg646 ?
                      wire568 : reg580) << $unsigned(reg613)) > (wire572[(1'h1):(1'h1)] ?
                      {reg603} : ((8'ha5) ?
                          reg581 : reg576)))) : $unsigned(((8'hb1) || reg607[(3'h4):(3'h4)])));
              reg650 <= $signed($signed($signed(((reg637 ? reg645 : wire561) ?
                  (reg646 ? reg633 : (7'h41)) : (reg617 ? reg616 : wire564)))));
              reg651 <= (^reg621);
            end
        end
      if (((7'h40) ? {reg642} : reg622[(4'hf):(4'hc)]))
        begin
          if (reg599[(1'h0):(1'h0)])
            begin
              reg652 <= $unsigned(reg615[(3'h5):(1'h0)]);
            end
          else
            begin
              reg653 = (wire571 != $signed(($signed($signed(wire568)) >>> ($signed(reg613) - (reg573 & (7'h42))))));
              reg654 = (((reg577[(1'h0):(1'h0)] >>> reg619) << reg609[(4'hf):(2'h3)]) ^~ (reg609[(3'h5):(1'h0)] ?
                  {wire562} : (!$signed(forvar576))));
              reg655 <= $signed((~&{(&reg631[(1'h1):(1'h1)])}));
              reg656 = $unsigned(({reg632, reg579[(3'h5):(3'h4)]} && reg648));
            end
        end
      else
        begin
          reg652 <= reg616;
          for (forvar653 = (1'h0); (forvar653 < (2'h3)); forvar653 = (forvar653 + (1'h1)))
            begin
              reg655 <= ((^(((|reg609) ?
                          reg647[(2'h2):(1'h1)] : ((8'ha7) ? reg634 : reg641)) ?
                      $signed($signed((8'hbd))) : {(~&reg638), (~|wire568)})) ?
                  (!(((wire569 ?
                      reg618 : reg585) >>> ((8'hb1) || reg648)) - (~(reg653 ?
                      wire570 : reg643)))) : ($signed($unsigned($unsigned(forvar614))) ?
                      $signed((^~(~&reg588))) : ((~^(~^reg597)) ?
                          ((reg592 ?
                              reg602 : reg633) | $unsigned(reg644)) : $signed((forvar622 ?
                              reg590 : reg587)))));
              reg656 = (~&reg607[(1'h0):(1'h0)]);
              reg657 <= (-(($signed(reg601) ?
                  {(reg643 ? reg640 : wire561),
                      $signed(wire569)} : $signed((reg574 | reg652))) <<< reg617));
              reg658 <= (((-reg636) == (forvar614 ~^ $signed((|reg585)))) ?
                  reg598 : {reg573, forvar653[(1'h1):(1'h1)]});
            end
          for (forvar659 = (1'h0); (forvar659 < (2'h2)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 <= (~^$unsigned(reg579[(3'h4):(3'h4)]));
              reg661 <= $signed((reg645 ?
                  wire564 : (!(reg598[(4'hd):(3'h6)] ?
                      $signed(reg608) : reg631))));
              reg662 = reg651;
              reg663 = (reg604 ? (8'hb0) : $unsigned((8'ha2)));
              reg664 <= {$signed(((&reg575) ? reg630 : reg585[(1'h1):(1'h1)]))};
            end
          if ((^~{(8'hbe), (|reg603[(1'h1):(1'h0)])}))
            begin
              reg665 <= $signed(((reg589[(2'h3):(2'h3)] > ((reg630 <= reg637) >> (reg646 + reg609))) - $unsigned((^~reg588[(3'h4):(2'h2)]))));
              reg666 <= reg610[(2'h3):(2'h2)];
              reg667 = ((+(~&(!(~&reg607)))) >= $signed($unsigned(reg606)));
            end
          else
            begin
              reg665 <= reg621[(1'h0):(1'h0)];
              reg666 <= forvar576;
              reg668 <= reg658;
              reg669 <= reg646[(2'h3):(1'h1)];
              reg670 = ($unsigned({{$signed(forvar576)},
                  {$unsigned((8'had))}}) < ($unsigned((~^reg641)) >> reg620[(4'hd):(1'h1)]));
            end
          reg671 <= $unsigned((~|reg645[(3'h7):(1'h0)]));
        end
    end
  assign wire672 = $signed(((reg648 ? reg664[(4'hc):(4'hc)] : reg625) ?
                       ($unsigned($unsigned(reg647)) >>> wire568[(2'h3):(1'h1)]) : reg584[(1'h1):(1'h1)]));
  assign wire673 = $unsigned($signed(($unsigned($unsigned((8'ha6))) > reg617[(3'h5):(2'h3)])));
  assign wire674 = (reg621 >>> (($signed((reg657 || reg578)) ?
                           ((reg630 ? reg644 : reg644) ?
                               $unsigned(reg618) : reg580) : reg634[(4'ha):(1'h0)]) ?
                       ($signed($signed(reg620)) != $unsigned((reg669 || reg647))) : ($unsigned($signed(wire569)) ?
                           wire562 : $unsigned(wire563[(3'h7):(3'h6)]))));
  always
    @(posedge clk) begin
      reg675 <= reg642[(3'h4):(1'h0)];
      if ($signed((&(((+(8'hab)) ?
          reg608 : $signed((8'hba))) >= $signed(reg608[(4'h9):(2'h3)])))))
        begin
          for (forvar676 = (1'h0); (forvar676 < (2'h2)); forvar676 = (forvar676 + (1'h1)))
            begin
              reg677 <= {(~reg644[(4'h9):(4'h9)])};
            end
          if (reg628[(5'h12):(5'h10)])
            begin
              reg678 = (^~(7'h40));
              reg679 <= ((~^$unsigned((^{(8'hb0)}))) >> (($unsigned(reg677[(4'h9):(1'h0)]) <= ((reg665 >>> reg590) ?
                      $unsigned(reg648) : {reg596})) ?
                  (&forvar676) : $signed({(reg631 ^ reg612),
                      (reg675 && reg608)})));
              reg680 <= $signed(wire563);
              reg681 <= (((wire564[(3'h7):(3'h6)] | ({wire672, reg669} ?
                          wire674[(3'h5):(1'h0)] : (|(8'ha8)))) ?
                      (!reg651) : $signed((+(7'h44)))) ?
                  $signed(reg635[(2'h2):(2'h2)]) : reg645[(4'h8):(4'h8)]);
              reg682 = (reg585[(1'h0):(1'h0)] > ($signed({(~|reg635),
                      (reg668 ? reg623 : reg634)}) ?
                  (reg630[(1'h1):(1'h0)] ?
                      {reg668,
                          (reg596 ?
                              reg603 : wire673)} : ($signed(reg611) >> ((8'hac) ~^ wire674))) : $unsigned({(wire566 ?
                          reg604 : reg624)})));
            end
          else
            begin
              reg678 = reg642[(3'h4):(1'h0)];
              reg679 <= ((((~$unsigned(reg666)) <= {(!reg644)}) ?
                      wire674[(1'h0):(1'h0)] : $unsigned($unsigned(wire673[(2'h2):(1'h1)]))) ?
                  (~&$signed((|(wire566 == reg666)))) : (wire563 <= (~^(~&reg665[(3'h4):(3'h4)]))));
              reg682 = (reg604[(1'h0):(1'h0)] ?
                  reg634[(4'he):(3'h5)] : (&({{wire564},
                      (~&reg631)} >> reg669[(3'h5):(2'h2)])));
            end
          if ($unsigned(($signed({reg599[(1'h1):(1'h0)], $signed(reg608)}) ?
              $signed({reg606}) : (($signed(reg605) & (~&reg580)) ?
                  ((reg635 < reg660) <= reg599) : $signed(reg652[(2'h2):(2'h2)])))))
            begin
              reg683 <= reg597[(2'h2):(1'h0)];
              reg684 <= reg634;
              reg685 = $unsigned($unsigned(((&$unsigned(reg630)) && ($unsigned(reg680) ?
                  (reg578 ? reg625 : reg589) : $unsigned(reg599)))));
              reg686 <= $unsigned(reg626);
              reg687 = (|$signed(reg630[(1'h0):(1'h0)]));
            end
          else
            begin
              reg683 <= ($unsigned(($signed($unsigned(wire567)) ?
                      (~(reg608 && reg635)) : ($signed(reg685) ?
                          reg630[(3'h4):(1'h1)] : (reg611 + reg647)))) ?
                  {reg658, (8'ha3)} : reg666);
              reg684 <= (|($signed(reg578) ?
                  $unsigned({(+reg633)}) : wire672[(5'h13):(3'h5)]));
              reg686 <= (~^reg625);
              reg688 <= reg635[(2'h2):(2'h2)];
            end
        end
      else
        begin
          if ($signed($unsigned(((reg628 <<< (^(8'haa))) ~^ $unsigned((wire566 ?
              (8'ha2) : reg681))))))
            begin
              reg676 <= $unsigned(((reg645 || $unsigned($signed(wire570))) ?
                  reg593[(5'h10):(4'h9)] : (-reg677)));
              reg677 <= reg657[(1'h0):(1'h0)];
              reg679 <= $unsigned((^~$unsigned(({(8'hb5), reg676} ?
                  {reg658} : $unsigned(reg607)))));
              reg680 <= reg588[(1'h1):(1'h0)];
            end
          else
            begin
              reg678 = reg666[(3'h4):(2'h2)];
              reg682 = $signed((7'h43));
              reg683 <= $signed((reg643 ?
                  $unsigned($signed($unsigned(reg617))) : reg608));
            end
          for (forvar684 = (1'h0); (forvar684 < (3'h4)); forvar684 = (forvar684 + (1'h1)))
            begin
              reg686 <= (^(~^((8'had) & reg575[(3'h4):(3'h4)])));
              reg688 <= wire564;
              reg689 <= (^(^~$unsigned(((reg634 ? reg671 : reg650) ^~ {wire572,
                  (7'h41)}))));
              reg690 <= $signed($signed($signed($signed(reg577))));
            end
          for (forvar691 = (1'h0); (forvar691 < (3'h4)); forvar691 = (forvar691 + (1'h1)))
            begin
              reg692 <= (|reg682);
              reg693 = (|(~|$unsigned(reg676)));
              reg694 <= $signed($unsigned(reg658));
              reg695 = $unsigned(((^reg676) < (+reg595)));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module316
#(parameter param556 = ((8'ha4) >= ((~&(^~{(8'h9c)})) ? ((((8'had) == (8'ha9)) ? (&(8'hb8)) : (^(8'hb5))) == (((8'hb3) ? (7'h41) : (8'hb5)) <= ((8'hbb) ? (7'h40) : (8'ha6)))) : ((((8'ha5) ? (7'h40) : (8'hbb)) ? (-(7'h41)) : ((8'haa) ? (8'hbb) : (8'ha9))) ? (|(7'h44)) : (8'hb2)))))
(y, clk, wire320, wire319, wire318, wire317);
  output wire [(32'haff):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire320;
  input wire [(4'ha):(1'h0)] wire319;
  input wire signed [(5'h15):(1'h0)] wire318;
  input wire signed [(2'h3):(1'h0)] wire317;
  wire signed [(4'hd):(1'h0)] wire555;
  wire signed [(3'h5):(1'h0)] wire481;
  wire [(5'h11):(1'h0)] wire480;
  wire signed [(4'hc):(1'h0)] wire389;
  wire signed [(4'hb):(1'h0)] wire388;
  wire [(4'hb):(1'h0)] wire387;
  wire signed [(4'h9):(1'h0)] wire386;
  wire [(5'h15):(1'h0)] wire385;
  wire [(3'h7):(1'h0)] wire321;
  reg [(4'h9):(1'h0)] reg554 = (1'h0);
  reg [(2'h3):(1'h0)] reg553 = (1'h0);
  reg [(5'h10):(1'h0)] reg551 = (1'h0);
  reg [(5'h10):(1'h0)] reg550 = (1'h0);
  reg [(3'h5):(1'h0)] reg549 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg548 = (1'h0);
  reg [(2'h3):(1'h0)] reg544 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg543 = (1'h0);
  reg [(4'he):(1'h0)] reg541 = (1'h0);
  reg [(5'h10):(1'h0)] reg538 = (1'h0);
  reg [(4'h8):(1'h0)] reg537 = (1'h0);
  reg [(5'h14):(1'h0)] reg532 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg531 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg530 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg526 = (1'h0);
  reg [(4'he):(1'h0)] reg524 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg523 = (1'h0);
  reg [(4'hf):(1'h0)] reg519 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg518 = (1'h0);
  reg [(5'h12):(1'h0)] reg517 = (1'h0);
  reg [(5'h12):(1'h0)] reg513 = (1'h0);
  reg [(2'h3):(1'h0)] reg512 = (1'h0);
  reg [(4'hd):(1'h0)] reg511 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg509 = (1'h0);
  reg [(4'hc):(1'h0)] reg507 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg506 = (1'h0);
  reg [(4'hb):(1'h0)] reg504 = (1'h0);
  reg signed [(4'he):(1'h0)] reg502 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg499 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg497 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg494 = (1'h0);
  reg [(3'h6):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg491 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg488 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg487 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg486 = (1'h0);
  reg [(3'h4):(1'h0)] reg485 = (1'h0);
  reg signed [(4'he):(1'h0)] reg483 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg479 = (1'h0);
  reg [(4'hb):(1'h0)] reg477 = (1'h0);
  reg [(5'h14):(1'h0)] reg473 = (1'h0);
  reg [(5'h14):(1'h0)] reg472 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg470 = (1'h0);
  reg [(4'h8):(1'h0)] reg468 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg467 = (1'h0);
  reg [(4'he):(1'h0)] reg465 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg464 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg463 = (1'h0);
  reg [(3'h5):(1'h0)] reg462 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg457 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg456 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg453 = (1'h0);
  reg [(4'h8):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg446 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg441 = (1'h0);
  reg [(5'h10):(1'h0)] reg440 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg439 = (1'h0);
  reg [(5'h15):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg436 = (1'h0);
  reg [(5'h14):(1'h0)] reg434 = (1'h0);
  reg [(4'hb):(1'h0)] reg431 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg430 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg417 = (1'h0);
  reg [(5'h14):(1'h0)] reg428 = (1'h0);
  reg [(5'h10):(1'h0)] reg425 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg422 = (1'h0);
  reg [(4'hb):(1'h0)] reg419 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg414 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg413 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg412 = (1'h0);
  reg [(3'h7):(1'h0)] reg410 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg409 = (1'h0);
  reg [(5'h15):(1'h0)] reg403 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg402 = (1'h0);
  reg [(2'h3):(1'h0)] reg401 = (1'h0);
  reg [(4'he):(1'h0)] reg399 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg397 = (1'h0);
  reg signed [(4'he):(1'h0)] reg396 = (1'h0);
  reg [(4'ha):(1'h0)] reg394 = (1'h0);
  reg [(4'hb):(1'h0)] reg393 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg380 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg379 = (1'h0);
  reg [(5'h13):(1'h0)] reg376 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg375 = (1'h0);
  reg [(5'h15):(1'h0)] reg374 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg368 = (1'h0);
  reg [(2'h3):(1'h0)] reg366 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg361 = (1'h0);
  reg [(5'h14):(1'h0)] reg360 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg359 = (1'h0);
  reg [(5'h10):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg356 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg355 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg353 = (1'h0);
  reg [(2'h3):(1'h0)] reg350 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg351 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg349 = (1'h0);
  reg [(3'h7):(1'h0)] reg345 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg344 = (1'h0);
  reg [(5'h12):(1'h0)] reg343 = (1'h0);
  reg [(3'h7):(1'h0)] reg340 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg337 = (1'h0);
  reg [(3'h5):(1'h0)] reg336 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg335 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg333 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg330 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg329 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg328 = (1'h0);
  reg [(5'h13):(1'h0)] reg326 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg325 = (1'h0);
  reg [(5'h12):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar552 = (1'h0);
  reg [(4'hb):(1'h0)] reg547 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg546 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar545 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar542 = (1'h0);
  reg [(5'h14):(1'h0)] reg525 = (1'h0);
  reg [(2'h2):(1'h0)] forvar540 = (1'h0);
  reg [(4'ha):(1'h0)] reg539 = (1'h0);
  reg [(4'h8):(1'h0)] reg536 = (1'h0);
  reg [(3'h7):(1'h0)] reg535 = (1'h0);
  reg [(3'h7):(1'h0)] reg534 = (1'h0);
  reg [(4'hb):(1'h0)] reg533 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg527 = (1'h0);
  reg [(5'h14):(1'h0)] forvar525 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg522 = (1'h0);
  reg signed [(4'he):(1'h0)] reg521 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg520 = (1'h0);
  reg [(5'h10):(1'h0)] reg516 = (1'h0);
  reg [(3'h4):(1'h0)] forvar515 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg514 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg508 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg503 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg501 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar500 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg498 = (1'h0);
  reg [(5'h10):(1'h0)] reg496 = (1'h0);
  reg [(5'h12):(1'h0)] reg495 = (1'h0);
  reg [(5'h15):(1'h0)] reg493 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg490 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg489 = (1'h0);
  reg [(4'hf):(1'h0)] reg484 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg482 = (1'h0);
  reg [(4'hb):(1'h0)] reg478 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg476 = (1'h0);
  reg [(4'hb):(1'h0)] reg475 = (1'h0);
  reg [(5'h12):(1'h0)] forvar474 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar471 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg469 = (1'h0);
  reg [(4'h8):(1'h0)] reg466 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg461 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg460 = (1'h0);
  reg [(2'h3):(1'h0)] reg459 = (1'h0);
  reg [(4'h9):(1'h0)] forvar455 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg454 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg452 = (1'h0);
  reg [(4'he):(1'h0)] reg451 = (1'h0);
  reg [(4'h9):(1'h0)] reg450 = (1'h0);
  reg [(4'h8):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg447 = (1'h0);
  reg [(4'hd):(1'h0)] reg445 = (1'h0);
  reg [(4'ha):(1'h0)] reg444 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg443 = (1'h0);
  reg [(5'h12):(1'h0)] reg442 = (1'h0);
  reg [(4'hd):(1'h0)] reg435 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar433 = (1'h0);
  reg [(4'hb):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar429 = (1'h0);
  reg [(4'hf):(1'h0)] forvar421 = (1'h0);
  reg [(2'h2):(1'h0)] reg427 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg426 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg424 = (1'h0);
  reg [(4'hb):(1'h0)] reg423 = (1'h0);
  reg [(5'h10):(1'h0)] reg421 = (1'h0);
  reg [(3'h7):(1'h0)] reg420 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar417 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg415 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg411 = (1'h0);
  reg [(4'h9):(1'h0)] reg408 = (1'h0);
  reg [(4'hf):(1'h0)] forvar407 = (1'h0);
  reg [(5'h10):(1'h0)] reg406 = (1'h0);
  reg [(4'ha):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar400 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg400 = (1'h0);
  reg [(3'h7):(1'h0)] reg398 = (1'h0);
  reg signed [(4'he):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg392 = (1'h0);
  reg [(4'hd):(1'h0)] forvar390 = (1'h0);
  reg [(4'hf):(1'h0)] reg384 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg381 = (1'h0);
  reg [(3'h7):(1'h0)] forvar378 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg377 = (1'h0);
  reg [(5'h10):(1'h0)] forvar373 = (1'h0);
  reg [(5'h10):(1'h0)] forvar372 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg371 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar370 = (1'h0);
  reg signed [(4'he):(1'h0)] reg369 = (1'h0);
  reg [(2'h3):(1'h0)] reg367 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg365 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg363 = (1'h0);
  reg [(5'h12):(1'h0)] reg362 = (1'h0);
  reg [(4'h8):(1'h0)] reg358 = (1'h0);
  reg [(4'hb):(1'h0)] reg354 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg352 = (1'h0);
  reg [(5'h15):(1'h0)] forvar350 = (1'h0);
  reg [(5'h13):(1'h0)] reg348 = (1'h0);
  reg [(5'h15):(1'h0)] reg347 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg346 = (1'h0);
  reg [(4'h8):(1'h0)] reg342 = (1'h0);
  reg [(5'h10):(1'h0)] forvar341 = (1'h0);
  reg [(4'hf):(1'h0)] reg339 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg338 = (1'h0);
  reg [(4'hf):(1'h0)] forvar329 = (1'h0);
  reg [(5'h14):(1'h0)] reg334 = (1'h0);
  reg [(4'hb):(1'h0)] reg332 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg331 = (1'h0);
  reg [(2'h3):(1'h0)] reg327 = (1'h0);
  reg [(4'hd):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg322 = (1'h0);
  assign y = {wire555,
                 wire481,
                 wire480,
                 wire389,
                 wire388,
                 wire387,
                 wire386,
                 wire385,
                 wire321,
                 reg554,
                 reg553,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg544,
                 reg543,
                 reg541,
                 reg538,
                 reg537,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg526,
                 reg524,
                 reg523,
                 reg519,
                 reg518,
                 reg517,
                 reg513,
                 reg512,
                 reg511,
                 reg509,
                 reg507,
                 reg506,
                 reg504,
                 reg502,
                 reg499,
                 reg497,
                 reg494,
                 reg492,
                 reg491,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg483,
                 reg479,
                 reg477,
                 reg473,
                 reg472,
                 reg470,
                 reg468,
                 reg467,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg458,
                 reg457,
                 reg456,
                 reg453,
                 reg448,
                 reg446,
                 reg433,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg434,
                 reg431,
                 reg430,
                 reg417,
                 reg428,
                 reg425,
                 reg422,
                 reg419,
                 reg418,
                 reg416,
                 reg414,
                 reg413,
                 reg412,
                 reg410,
                 reg409,
                 reg403,
                 reg402,
                 reg401,
                 reg399,
                 reg397,
                 reg396,
                 reg394,
                 reg393,
                 reg391,
                 reg383,
                 reg382,
                 reg380,
                 reg379,
                 reg376,
                 reg375,
                 reg374,
                 reg368,
                 reg366,
                 reg364,
                 reg361,
                 reg360,
                 reg359,
                 reg357,
                 reg356,
                 reg355,
                 reg353,
                 reg350,
                 reg351,
                 reg349,
                 reg345,
                 reg344,
                 reg343,
                 reg340,
                 reg337,
                 reg336,
                 reg335,
                 reg333,
                 reg330,
                 reg329,
                 reg328,
                 reg326,
                 reg325,
                 reg324,
                 forvar552,
                 reg547,
                 reg546,
                 forvar545,
                 forvar542,
                 reg525,
                 forvar540,
                 reg539,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 reg527,
                 forvar525,
                 reg522,
                 reg521,
                 reg520,
                 reg516,
                 forvar515,
                 reg514,
                 reg510,
                 reg508,
                 reg505,
                 reg503,
                 reg501,
                 forvar500,
                 reg498,
                 reg496,
                 reg495,
                 reg493,
                 reg490,
                 reg489,
                 reg484,
                 reg482,
                 reg478,
                 reg476,
                 reg475,
                 forvar474,
                 forvar471,
                 reg469,
                 reg466,
                 reg461,
                 reg460,
                 reg459,
                 forvar455,
                 reg454,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg447,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg435,
                 forvar433,
                 reg432,
                 forvar429,
                 forvar421,
                 reg427,
                 reg426,
                 reg424,
                 reg423,
                 reg421,
                 reg420,
                 forvar417,
                 reg415,
                 reg411,
                 reg408,
                 forvar407,
                 reg406,
                 reg405,
                 reg404,
                 forvar400,
                 reg400,
                 reg398,
                 reg395,
                 reg392,
                 forvar390,
                 reg384,
                 reg381,
                 forvar378,
                 reg377,
                 forvar373,
                 forvar372,
                 reg371,
                 forvar370,
                 reg369,
                 reg367,
                 reg365,
                 reg363,
                 reg362,
                 reg358,
                 reg354,
                 reg352,
                 forvar350,
                 reg348,
                 reg347,
                 reg346,
                 reg342,
                 forvar341,
                 reg339,
                 reg338,
                 forvar329,
                 reg334,
                 reg332,
                 reg331,
                 reg327,
                 reg323,
                 reg322,
                 (1'h0)};
  assign wire321 = $unsigned(($unsigned({$unsigned((8'hb5)),
                       (wire320 ?
                           wire317 : wire319)}) ^ (((wire320 && wire320) ?
                           wire319[(3'h5):(1'h0)] : (8'ha7)) ?
                       (&(wire320 > wire320)) : $signed(((8'hac) ?
                           wire317 : wire317)))));
  always
    @(posedge clk) begin
      if (((^~$unsigned(wire317[(1'h1):(1'h0)])) ?
          wire321 : (~^wire318[(2'h2):(1'h0)])))
        begin
          if ($signed((|$unsigned($unsigned((wire320 <= wire317))))))
            begin
              reg322 = $signed(wire317);
              reg323 = ($signed($signed((&(-reg322)))) <= $unsigned(((!$unsigned(wire318)) ?
                  (8'hbb) : $unsigned($unsigned(wire320)))));
              reg324 <= ((wire320[(1'h0):(1'h0)] >>> reg323) ?
                  wire319[(2'h3):(2'h2)] : (-$signed(($unsigned(wire318) ?
                      (wire317 ? wire321 : reg322) : (reg322 ?
                          (8'hb1) : wire319)))));
              reg325 <= {(~^$signed(({reg322, wire318} ?
                      (reg323 ? wire320 : wire318) : (reg324 >= wire318))))};
              reg326 <= reg323;
            end
          else
            begin
              reg324 <= (wire319 && (({(reg322 ? reg326 : wire317),
                  (|wire318)} >> (wire318 ?
                  $signed(reg322) : reg325)) + wire319));
              reg325 <= $unsigned($unsigned($unsigned((&wire320[(2'h2):(1'h0)]))));
            end
          reg327 = $unsigned(wire321);
          if (((&$signed(($unsigned(reg322) ?
              (wire317 ?
                  wire317 : reg322) : ((8'ha3) | wire317)))) >>> ($signed({reg324[(3'h6):(2'h2)]}) ?
              reg325 : ((^(-reg327)) ?
                  (^~((8'hbd) != wire320)) : reg322[(5'h14):(4'h8)]))))
            begin
              reg328 <= wire320;
              reg329 <= (^$signed(reg324));
              reg330 <= ({({(8'ha1)} != {$unsigned(reg322),
                      (wire319 > reg322)}),
                  ($unsigned((reg326 ?
                      reg326 : reg327)) == (!$signed(reg322)))} && reg328[(2'h2):(2'h2)]);
            end
          else
            begin
              reg331 = ({wire317[(2'h3):(2'h2)],
                  $signed(reg327[(1'h1):(1'h1)])} >= (reg330 ?
                  (reg329 <<< reg326[(3'h4):(3'h4)]) : ($unsigned({reg327,
                          reg327}) ?
                      (!{reg329}) : (&(reg322 ? reg322 : (8'h9c))))));
              reg332 = (^~$unsigned($unsigned($signed($signed(reg323)))));
              reg333 <= $signed($signed($unsigned((~|(~^wire321)))));
              reg334 = ($unsigned((reg329[(3'h4):(3'h4)] ?
                  reg324 : $unsigned($unsigned(reg322)))) ~^ $unsigned(((&{(8'hb4),
                  reg330}) | wire321[(2'h3):(2'h3)])));
            end
        end
      else
        begin
          if (wire320)
            begin
              reg322 = {reg330};
              reg324 <= {(+$signed((^(reg332 <= reg326))))};
              reg327 = $unsigned(((^~(~|$unsigned(reg325))) || reg326));
            end
          else
            begin
              reg324 <= $signed({(((&(7'h42)) ?
                          (reg322 ? reg333 : reg331) : (|wire321)) ?
                      $signed((8'hbb)) : (reg332 == (reg330 ?
                          reg331 : reg333)))});
              reg325 <= wire317[(2'h3):(2'h3)];
              reg326 <= $unsigned($signed(((-$signed(wire317)) ^ $unsigned(reg330))));
              reg328 <= {(|$unsigned(wire320[(1'h1):(1'h1)])),
                  ((+((~^reg330) ?
                      reg328 : $signed(reg327))) != (~^$unsigned((reg334 < reg326))))};
            end
          for (forvar329 = (1'h0); (forvar329 < (2'h2)); forvar329 = (forvar329 + (1'h1)))
            begin
              reg330 <= (~&(((8'h9f) || (reg323[(2'h3):(1'h1)] ^ (reg323 ?
                      reg329 : wire320))) ?
                  ($signed((!wire317)) + wire320) : ((reg322[(2'h3):(2'h2)] ?
                          $signed((8'ha1)) : $signed(wire318)) ?
                      reg331 : ((^~reg332) >> (reg327 ? reg333 : reg328)))));
              reg331 = $signed($signed((8'ha9)));
              reg333 <= (reg323 && reg330[(2'h2):(2'h2)]);
              reg335 <= wire321[(3'h5):(1'h1)];
              reg336 <= forvar329;
            end
          if (({$signed(reg331)} <= $unsigned($unsigned(($signed(reg322) ?
              $unsigned(wire320) : (reg327 ? wire319 : reg332))))))
            begin
              reg337 <= $signed($unsigned(((wire320 << reg329[(3'h5):(2'h2)]) ?
                  {(reg328 ? (8'ha4) : reg326)} : (^$unsigned(reg333)))));
              reg338 = ((($signed($unsigned(reg331)) >> wire321) ^~ {$signed(reg336),
                  (~{reg328, reg325})}) < $unsigned(reg336));
              reg339 = reg330[(2'h2):(1'h1)];
              reg340 <= reg329[(1'h1):(1'h0)];
            end
          else
            begin
              reg337 <= (!(reg327[(2'h3):(1'h1)] ?
                  {((reg323 - reg326) <<< reg340[(3'h5):(2'h3)]),
                      (wire319 ?
                          ((8'hbb) ? wire318 : wire318) : (wire321 ?
                              reg327 : wire320))} : $signed((reg325[(1'h1):(1'h1)] || reg329[(2'h2):(2'h2)]))));
            end
          for (forvar341 = (1'h0); (forvar341 < (2'h2)); forvar341 = (forvar341 + (1'h1)))
            begin
              reg342 = wire318[(3'h7):(3'h5)];
              reg343 <= ($signed($signed(reg326)) > reg333);
            end
          if (($signed(wire320[(2'h2):(1'h1)]) ?
              (~^$unsigned(({reg327, reg338} ?
                  ((8'hb5) ?
                      wire319 : wire319) : reg340[(3'h5):(3'h4)]))) : $unsigned(($unsigned($signed(reg337)) ?
                  ($unsigned((7'h41)) ?
                      (reg333 >= reg323) : $signed(reg322)) : (wire318[(5'h12):(4'hb)] ?
                      (forvar341 || (8'ha2)) : (reg332 ? wire317 : reg333))))))
            begin
              reg344 <= $unsigned({reg342[(1'h0):(1'h0)],
                  $signed((~&(reg324 ? forvar341 : reg335)))});
              reg345 <= (reg344[(3'h7):(2'h2)] & $signed(wire319));
            end
          else
            begin
              reg346 = (forvar329 && $signed($unsigned(wire319[(3'h7):(1'h1)])));
              reg347 = (reg339[(3'h7):(3'h6)] ^~ reg333[(1'h0):(1'h0)]);
              reg348 = reg326;
              reg349 <= (-$unsigned({reg342}));
            end
        end
      if (($signed(reg338) || $unsigned((8'hae))))
        begin
          for (forvar350 = (1'h0); (forvar350 < (2'h2)); forvar350 = (forvar350 + (1'h1)))
            begin
              reg351 <= {reg344, reg349};
              reg352 = ($signed($unsigned((reg335 <= wire319[(1'h1):(1'h0)]))) ?
                  reg343[(4'h8):(3'h6)] : (-$signed($signed($signed(reg335)))));
            end
        end
      else
        begin
          if ((^~$unsigned({(reg336 ? $signed((7'h40)) : $signed(reg345)),
              (reg345[(3'h5):(2'h3)] ? $unsigned(reg338) : reg332)})))
            begin
              reg350 <= $unsigned($unsigned($unsigned((~|reg344))));
            end
          else
            begin
              reg352 = reg350[(1'h0):(1'h0)];
              reg353 <= reg340;
            end
          reg354 = $signed(({(&$signed((7'h40)))} ?
              (8'hb4) : reg322[(4'hb):(4'h9)]));
          if (wire317)
            begin
              reg355 <= wire320;
              reg356 <= (8'hb6);
              reg357 <= $signed($signed(($unsigned($signed(wire318)) ?
                  $signed(wire319[(3'h4):(1'h1)]) : $unsigned(wire320))));
            end
          else
            begin
              reg355 <= (~^$signed(({reg345} >= ($signed(reg332) ?
                  (~&reg355) : reg345))));
              reg356 <= (|reg350);
            end
        end
      if ((reg345[(2'h2):(2'h2)] ^~ $unsigned(($unsigned({reg328}) <= (8'hba)))))
        begin
          if ({((-$signed(((8'ha5) << reg355))) ?
                  {(~&$unsigned((8'ha0))),
                      $unsigned((!reg325))} : (&(~$signed(reg348)))),
              $signed(reg350[(1'h1):(1'h0)])})
            begin
              reg358 = {($unsigned({$signed(reg340), wire320[(2'h2):(1'h0)]}) ?
                      (+reg355) : reg322[(3'h6):(1'h0)])};
            end
          else
            begin
              reg359 <= $unsigned(reg351[(4'h8):(3'h4)]);
              reg360 <= {$unsigned(reg331[(2'h3):(2'h2)]),
                  (reg323[(4'hc):(4'hb)] >>> reg357[(3'h6):(1'h1)])};
              reg361 <= reg348[(4'hb):(4'h8)];
              reg362 = ((reg343 ?
                  (reg351 >> ((~|reg342) << $signed(forvar350))) : (8'h9e)) != (($signed((reg342 > reg344)) ?
                      reg326[(5'h10):(4'hd)] : reg346[(1'h0):(1'h0)]) ?
                  forvar329 : (+(-reg342[(2'h3):(1'h0)]))));
            end
          if ((^($signed($unsigned(((8'hbb) <= (8'hb7)))) ?
              $unsigned(((reg332 ?
                  (8'ha2) : (7'h44)) - (wire317 || wire317))) : (~&(^reg329)))))
            begin
              reg363 = reg357[(1'h1):(1'h0)];
              reg364 <= (^(forvar329 ?
                  $unsigned(((reg330 ?
                      reg350 : (8'hb9)) >>> (reg337 & reg356))) : wire320));
              reg365 = (8'hbc);
              reg366 <= ((^~reg358) ?
                  {(((reg362 ? (8'h9d) : reg327) ?
                          (reg350 + reg326) : $unsigned(reg344)) >>> $unsigned(wire320[(1'h1):(1'h0)]))} : $signed($signed(reg339)));
            end
          else
            begin
              reg364 <= reg337[(1'h0):(1'h0)];
              reg366 <= (~$signed($unsigned(((reg335 ~^ reg324) != reg345[(3'h4):(2'h2)]))));
              reg367 = reg323;
            end
        end
      else
        begin
          if ({$signed((^((wire318 >= (8'h9d)) ? {reg338, reg324} : (8'hac)))),
              $unsigned($signed((^(-(8'hab)))))})
            begin
              reg358 = (|$signed(($signed(reg328[(4'ha):(3'h7)]) ?
                  (reg367 & (reg328 >= (8'haf))) : ((wire317 || forvar341) ?
                      {reg325, (8'hbb)} : (-(8'hb7))))));
              reg362 = $signed(forvar341[(4'he):(3'h6)]);
              reg363 = reg361[(1'h1):(1'h1)];
              reg364 <= reg355;
              reg366 <= (((~({(8'hb9), reg349} == (8'ha5))) ?
                  (((~reg361) ? $unsigned(reg367) : reg329) ?
                      $signed((reg338 ? reg337 : reg330)) : {(reg355 || reg324),
                          reg364}) : reg322[(5'h11):(3'h4)]) && reg327);
            end
          else
            begin
              reg358 = (~{((reg340[(3'h4):(1'h1)] ?
                          (|reg350) : $signed(reg365)) ?
                      (~|(reg335 ? (8'h9c) : reg339)) : (^~$signed((8'hbf)))),
                  ((forvar350 ? forvar329[(3'h7):(3'h4)] : $signed(reg353)) ?
                      $signed(reg326) : reg363)});
              reg359 <= reg343;
            end
          if (reg346)
            begin
              reg367 = $unsigned((((reg347[(5'h13):(3'h4)] > (|reg344)) < $signed($unsigned(reg344))) ^ wire321[(3'h5):(3'h5)]));
            end
          else
            begin
              reg367 = (&{$signed({{reg322}}),
                  ($signed(reg363[(4'ha):(1'h0)]) ?
                      $signed(reg348[(3'h4):(1'h0)]) : ((forvar329 ?
                          wire318 : (7'h44)) + (~&reg358)))});
              reg368 <= $unsigned(($signed($signed($unsigned(reg351))) && reg331));
              reg369 = {reg347[(5'h12):(4'h8)],
                  $unsigned(({(~^reg331), (reg335 >> (8'ha6))} ?
                      reg353[(3'h4):(2'h2)] : forvar350[(4'hb):(4'h9)]))};
            end
          for (forvar370 = (1'h0); (forvar370 < (2'h3)); forvar370 = (forvar370 + (1'h1)))
            begin
              reg371 = reg337[(1'h1):(1'h0)];
            end
        end
      for (forvar372 = (1'h0); (forvar372 < (3'h4)); forvar372 = (forvar372 + (1'h1)))
        begin
          for (forvar373 = (1'h0); (forvar373 < (1'h0)); forvar373 = (forvar373 + (1'h1)))
            begin
              reg374 <= ($unsigned((wire321[(2'h2):(1'h0)] ?
                  $signed((reg369 != reg346)) : reg361)) >= {(~^(+$unsigned((8'ha6))))});
              reg375 <= (reg371[(4'hd):(4'hb)] ?
                  ($unsigned(({(8'h9e), reg332} <= $unsigned(reg358))) ?
                      (reg345 ?
                          $signed(((8'haa) ? reg364 : (8'hba))) : (reg354 ?
                              $unsigned(wire320) : wire317)) : {(wire318[(1'h0):(1'h0)] ?
                              $signed((8'h9c)) : $unsigned(reg333))}) : ((!$signed(forvar350)) ?
                      (reg365 >= (|wire317)) : reg328[(4'hf):(4'ha)]));
              reg376 <= (~^$unsigned(reg367[(1'h1):(1'h1)]));
              reg377 = $unsigned((+{(reg343[(4'h9):(2'h2)] != (8'ha0))}));
            end
          for (forvar378 = (1'h0); (forvar378 < (1'h1)); forvar378 = (forvar378 + (1'h1)))
            begin
              reg379 <= $unsigned(($unsigned(((forvar341 >> reg352) & reg329)) << $signed((8'hba))));
              reg380 <= reg339[(3'h7):(2'h3)];
              reg381 = (((8'ha6) ?
                  (reg375[(2'h3):(1'h1)] < $signed((forvar341 ?
                      reg339 : reg353))) : forvar373[(4'hd):(3'h7)]) <<< forvar373[(4'hc):(2'h3)]);
              reg382 <= reg361[(3'h5):(3'h5)];
              reg383 <= (((((forvar341 > reg334) ? reg326 : (-(8'hb0))) ?
                      (reg375 ?
                          (reg330 >= reg349) : (~|forvar329)) : reg333[(2'h2):(1'h1)]) || reg323[(4'hb):(4'ha)]) ?
                  $unsigned(reg371[(4'h9):(3'h4)]) : ((wire317[(1'h0):(1'h0)] >> reg330[(2'h3):(2'h3)]) ?
                      (&{(|(8'ha1)), $unsigned(reg349)}) : (reg352 ?
                          (reg362 ?
                              (~|reg336) : $signed(reg366)) : $signed((reg366 ?
                              reg322 : reg328)))));
            end
        end
      reg384 = reg350[(1'h1):(1'h1)];
    end
  assign wire385 = ($signed($unsigned((~^(reg353 ? wire321 : reg353)))) ?
                       $signed((^((reg324 | reg361) >> $signed(reg375)))) : ((-(reg336 ?
                           (reg344 << reg382) : (reg382 ?
                               reg343 : reg324))) ^ ((^~reg345[(3'h6):(3'h4)]) ?
                           (+(&reg335)) : ($unsigned(reg364) | reg330[(2'h3):(1'h1)]))));
  assign wire386 = reg357;
  assign wire387 = $unsigned(wire318);
  assign wire388 = $unsigned($signed({((reg364 >> (8'hb6)) << $signed((8'ha7))),
                       (-reg345)}));
  assign wire389 = {$unsigned($unsigned(reg344[(1'h1):(1'h0)])),
                       ($signed(((8'hb7) || wire320[(2'h2):(2'h2)])) ?
                           (^(reg382 ?
                               $unsigned((8'hb8)) : (+reg380))) : $unsigned(reg333))};
  always
    @(posedge clk) begin
      for (forvar390 = (1'h0); (forvar390 < (1'h0)); forvar390 = (forvar390 + (1'h1)))
        begin
          if (reg376[(5'h10):(4'hd)])
            begin
              reg391 <= $unsigned((-$signed(((+reg330) ?
                  $signed(reg361) : $unsigned((8'ha9))))));
            end
          else
            begin
              reg392 = reg359;
            end
          if ((($signed((~(reg340 >> (8'ha8)))) ?
              forvar390 : wire317) || (~|forvar390[(2'h2):(1'h0)])))
            begin
              reg393 <= (!reg383);
              reg394 <= reg324[(5'h12):(3'h7)];
              reg395 = $unsigned({(-((~&wire321) != $signed(reg333))),
                  (wire320[(2'h2):(2'h2)] ^~ ({reg366} - reg364[(1'h0):(1'h0)]))});
            end
          else
            begin
              reg395 = reg383;
              reg396 <= (~|$unsigned(($unsigned((reg380 && reg343)) ?
                  $unsigned(reg336) : reg345[(3'h6):(3'h4)])));
            end
          if ((($unsigned(wire317) <<< (8'ha8)) >= (^~wire386)))
            begin
              reg397 <= ({$signed((^~(&reg345)))} ?
                  reg355 : ($signed($signed($signed(reg343))) ?
                      ({$signed(reg356),
                          (reg360 ?
                              reg356 : wire388)} != {$unsigned(wire319)}) : ($unsigned((wire318 ?
                          reg356 : reg336)) & (8'hae))));
              reg398 = $unsigned(reg328);
              reg399 <= reg356;
            end
          else
            begin
              reg397 <= (~$signed(($unsigned(reg399) >>> {(reg330 ~^ reg380),
                  reg395[(4'hb):(2'h3)]})));
              reg399 <= reg345[(1'h1):(1'h0)];
            end
        end
      if ($signed(reg329))
        begin
          reg400 = reg376;
        end
      else
        begin
          for (forvar400 = (1'h0); (forvar400 < (2'h3)); forvar400 = (forvar400 + (1'h1)))
            begin
              reg401 <= $signed($unsigned(reg392[(4'ha):(1'h1)]));
              reg402 <= ({reg374, $signed({(+wire321), $unsigned(reg360)})} ?
                  reg380[(1'h1):(1'h0)] : (+{$signed($unsigned((8'hbd)))}));
              reg403 <= (reg368 ?
                  wire389 : ($unsigned(($signed(reg357) ?
                          (8'hb5) : (reg326 ? reg379 : wire318))) ?
                      reg397 : $unsigned(reg379)));
            end
          if (({$unsigned($unsigned({reg368, reg376}))} ?
              (($unsigned({wire388, reg345}) <<< wire318) ?
                  $signed($unsigned(((8'hae) ?
                      reg357 : (8'ha1)))) : (^~wire318[(3'h5):(3'h5)])) : (($unsigned((reg382 ?
                      wire320 : reg345)) && reg343[(5'h12):(4'hc)]) ?
                  $signed(((reg361 & reg382) ?
                      reg383[(3'h5):(1'h1)] : $signed((8'ha9)))) : (reg393 >> $signed((reg392 + reg344))))))
            begin
              reg404 = ($unsigned({((^~reg380) ? reg379 : {reg403, reg382}),
                      {$signed(reg374), (8'ha5)}}) ?
                  (7'h42) : {(8'ha2)});
              reg405 = (!(8'hb9));
              reg406 = (|reg391[(4'hb):(3'h5)]);
            end
          else
            begin
              reg404 = (8'hb9);
            end
          for (forvar407 = (1'h0); (forvar407 < (3'h4)); forvar407 = (forvar407 + (1'h1)))
            begin
              reg408 = $signed((~|({(!reg344)} >> (!{reg406}))));
              reg409 <= {(|(8'h9f)), (reg326 | $signed(reg404))};
              reg410 <= $unsigned(reg401);
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg357[(1'h0):(1'h0)])
        begin
          if (wire386[(3'h7):(1'h1)])
            begin
              reg411 = $unsigned({reg359[(2'h3):(1'h0)],
                  {reg394[(4'h9):(3'h4)]}});
              reg412 <= (&(^~($unsigned(reg335[(1'h1):(1'h0)]) ?
                  {(8'hb8)} : $unsigned((reg353 ^~ (8'ha2))))));
              reg413 <= $unsigned((~$signed(reg401[(1'h1):(1'h1)])));
              reg414 <= (^(8'h9f));
              reg415 = (($unsigned($signed(wire320[(1'h0):(1'h0)])) + (wire385[(3'h6):(3'h4)] - ((reg343 ?
                  (8'h9c) : reg364) & (reg412 & reg391)))) && {(reg350[(2'h3):(1'h0)] ?
                      $signed($unsigned(reg360)) : reg412[(3'h4):(2'h3)]),
                  $signed($unsigned((reg361 ? reg361 : wire389)))});
            end
          else
            begin
              reg412 <= {reg366,
                  $unsigned(($signed((reg414 + reg359)) - reg380))};
              reg413 <= (!$unsigned($unsigned({$signed(wire321), {(8'ha6)}})));
              reg414 <= (7'h43);
              reg416 <= reg414;
            end
          for (forvar417 = (1'h0); (forvar417 < (2'h2)); forvar417 = (forvar417 + (1'h1)))
            begin
              reg418 <= ((((~|$signed(reg329)) >> (8'hb9)) || $unsigned(($signed((7'h40)) ?
                  reg357[(1'h1):(1'h0)] : (8'hba)))) * (reg349[(1'h1):(1'h1)] ?
                  reg359 : reg335[(4'ha):(4'h9)]));
              reg419 <= reg336[(2'h3):(2'h3)];
              reg420 = reg335;
            end
          if ((^~$signed(({reg420[(1'h1):(1'h0)]} << (reg343[(4'hb):(4'h8)] << $signed(reg376))))))
            begin
              reg421 = $unsigned(reg340[(3'h6):(1'h0)]);
              reg422 <= reg391;
              reg423 = $unsigned(reg402[(1'h1):(1'h0)]);
              reg424 = (~|(reg375[(1'h1):(1'h0)] ?
                  $unsigned((reg351[(4'h8):(3'h7)] ?
                      {reg420} : (reg396 ?
                          wire319 : (8'hb9)))) : reg330[(3'h6):(3'h5)]));
              reg425 <= (&({reg420[(2'h2):(1'h1)]} && ($unsigned(reg401) ?
                  ((~&(7'h43)) ?
                      reg351 : (reg422 ? reg333 : reg376)) : reg399)));
            end
          else
            begin
              reg422 <= $unsigned(reg425);
              reg423 = (!(reg396[(4'hb):(4'h9)] ?
                  (reg376[(1'h0):(1'h0)] & reg329) : $unsigned((wire389 ?
                      $unsigned(reg335) : $unsigned((8'hba))))));
            end
          if (reg393)
            begin
              reg426 = reg394;
              reg427 = reg413;
              reg428 <= reg361;
            end
          else
            begin
              reg428 <= reg366[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg412 <= reg330;
          if ({((((reg411 ?
                      reg428 : reg411) == $unsigned(reg416)) & $signed({(8'hab),
                      reg324})) ?
                  $signed(wire317[(2'h2):(2'h2)]) : $signed($signed($unsigned(reg382)))),
              $unsigned((reg337 ? reg345[(3'h4):(2'h3)] : (8'hb5)))})
            begin
              reg413 <= ($unsigned(((reg382[(3'h5):(1'h1)] ?
                  (reg412 ?
                      reg410 : reg402) : $signed(reg343)) && (~(reg382 <= (8'hbe))))) >>> ($signed(((reg340 ?
                  wire385 : reg391) | (~&reg328))) & wire318[(3'h4):(2'h2)]));
              reg414 <= {($unsigned($unsigned((-reg326))) ?
                      (($signed(wire320) ?
                          (reg374 ?
                              reg423 : reg402) : reg335[(3'h6):(3'h4)]) << $unsigned((~(8'hbd)))) : (^~$signed((reg393 ?
                          reg425 : reg361)))),
                  $signed((reg324[(5'h12):(3'h5)] ?
                      (|reg414) : (reg411 ?
                          $signed(reg333) : ((8'ha5) ? reg343 : wire385))))};
              reg416 <= ((~$signed({((8'ha5) ?
                      (8'had) : reg328)})) == $unsigned((~^(-$signed(reg329)))));
            end
          else
            begin
              reg413 <= $unsigned(({$signed($signed((8'hb6)))} - reg330[(3'h6):(3'h6)]));
              reg414 <= ($signed(reg382) ?
                  $signed(reg415) : $unsigned((((~reg359) ?
                          $unsigned(wire321) : $signed(reg409)) ?
                      (reg350[(1'h1):(1'h1)] ?
                          $signed(reg423) : (forvar417 >> wire317)) : {$unsigned(reg325)})));
              reg416 <= ($signed(forvar417[(4'hb):(3'h5)]) ?
                  reg421[(4'h8):(3'h4)] : reg336[(3'h4):(1'h1)]);
              reg417 <= ((&($signed(wire386[(1'h1):(1'h1)]) ?
                  {reg374[(2'h3):(1'h1)]} : {$unsigned((8'hac))})) - reg423);
              reg420 = (($signed((-(reg343 >>> reg382))) ?
                  {$signed(reg426[(1'h0):(1'h0)])} : $signed((wire385[(5'h10):(3'h4)] == (~|reg344)))) <<< $signed($unsigned(($unsigned(reg428) ?
                  wire321[(3'h7):(1'h1)] : (reg403 ? reg351 : reg425)))));
            end
          for (forvar421 = (1'h0); (forvar421 < (1'h1)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg422 <= {(reg421[(3'h7):(1'h0)] + reg344[(1'h1):(1'h1)])};
              reg425 <= ({$signed($signed((reg374 ~^ (7'h40)))),
                  (~^$unsigned(reg340))} ^~ reg364[(2'h2):(1'h0)]);
            end
          if ($unsigned($signed(reg394)))
            begin
              reg426 = {{$unsigned(((reg360 <<< reg410) & (reg399 ?
                          reg403 : (7'h40))))},
                  (^$unsigned((~&(^reg375))))};
            end
          else
            begin
              reg428 <= $signed($signed((reg417 ?
                  (+(reg396 ~^ reg409)) : $signed((wire385 ?
                      reg375 : (8'ha9))))));
            end
          for (forvar429 = (1'h0); (forvar429 < (1'h1)); forvar429 = (forvar429 + (1'h1)))
            begin
              reg430 <= (~|(~($signed((reg421 ?
                  wire385 : (8'hb0))) | $unsigned(reg359))));
              reg431 <= (wire388 <= reg357);
              reg432 = $unsigned($signed(((~&$signed(reg355)) ?
                  (~^$unsigned(reg391)) : (~&{reg344, reg401}))));
            end
        end
      if ($unsigned((!(8'ha8))))
        begin
          for (forvar433 = (1'h0); (forvar433 < (1'h1)); forvar433 = (forvar433 + (1'h1)))
            begin
              reg434 <= ($signed(reg410[(3'h4):(1'h0)]) ^ ((wire389[(3'h7):(1'h0)] ?
                  ({reg431, forvar421} ?
                      reg402 : (8'ha7)) : $signed($unsigned(reg324))) ^ $signed(((reg355 ?
                      reg432 : wire320) ?
                  reg425 : (8'hb5)))));
              reg435 = (($unsigned($unsigned(reg403[(5'h15):(4'hb)])) | reg368[(3'h7):(2'h3)]) != (8'hbc));
              reg436 <= reg351;
              reg437 <= $unsigned(reg436);
            end
          if (reg416[(4'h9):(3'h5)])
            begin
              reg438 <= (((reg326 | $signed(reg415)) | (^~$signed((reg420 || (8'hb0))))) ?
                  reg419 : $unsigned($unsigned($unsigned({reg393}))));
              reg439 <= {(($unsigned($unsigned(reg391)) && reg420[(3'h6):(1'h0)]) < $unsigned(wire385[(4'h8):(1'h0)]))};
              reg440 <= $unsigned(($signed(reg419) & reg436[(1'h0):(1'h0)]));
              reg441 <= $unsigned($signed(reg418));
              reg442 = ($signed(reg428[(4'hb):(4'h8)]) & (|($unsigned(reg361) ?
                  $signed(wire385[(4'he):(3'h5)]) : ((7'h40) ?
                      $signed(reg344) : wire319))));
            end
          else
            begin
              reg442 = $unsigned(reg418[(3'h5):(1'h1)]);
              reg443 = (reg396[(3'h4):(3'h4)] + {$unsigned(($unsigned((8'h9f)) ?
                      reg356 : (reg353 ? (8'hbe) : reg421)))});
            end
        end
      else
        begin
          reg433 <= reg329[(3'h7):(1'h0)];
        end
      reg444 = reg401[(2'h2):(1'h0)];
      if (((!($signed(reg333) <<< $signed($unsigned((8'ha2))))) ?
          forvar429 : (8'ha9)))
        begin
          if ($signed($unsigned((~^$signed(reg399)))))
            begin
              reg445 = (8'hb1);
              reg446 <= reg410[(3'h7):(1'h1)];
              reg447 = (($unsigned(({reg360, reg396} ?
                  $unsigned(reg416) : wire318)) > (wire389[(4'h8):(2'h2)] ?
                  ((wire387 - (7'h43)) ?
                      (8'ha2) : (reg402 ?
                          reg350 : reg366)) : $signed(reg345[(3'h4):(3'h4)]))) >>> $unsigned($unsigned({(reg397 || reg391)})));
              reg448 <= (~^reg444[(4'h9):(2'h3)]);
            end
          else
            begin
              reg446 <= ((reg391 ?
                  ((-(~&reg353)) != $signed(((8'hb8) ?
                      reg441 : reg361))) : $signed({$signed(reg426)})) ~^ ((((reg421 ?
                      reg441 : reg396) == (^~reg336)) ?
                  $signed((8'hb8)) : (~|wire321)) && ({(reg437 <= reg399)} > $unsigned({reg351}))));
              reg448 <= reg432;
            end
          if (reg351[(1'h1):(1'h1)])
            begin
              reg449 = $signed((|$unsigned(wire388[(1'h0):(1'h0)])));
              reg450 = ($unsigned((8'h9c)) ?
                  $unsigned({(&reg380[(2'h3):(2'h2)]),
                      wire321[(1'h1):(1'h1)]}) : (($unsigned($unsigned(reg423)) ?
                      (&((8'hb3) == reg411)) : (+(^~reg391))) == {{$unsigned((8'hb2)),
                          (^reg443)}}));
              reg451 = $signed((~^$unsigned((-(forvar433 ?
                  wire387 : reg382)))));
              reg452 = ((($signed($unsigned((7'h44))) & (^((8'ha4) ?
                      (8'hae) : reg432))) ?
                  wire317[(1'h0):(1'h0)] : reg412) >= $signed((($unsigned(reg344) * (8'hae)) ?
                  reg447 : (^~(^reg375)))));
            end
          else
            begin
              reg453 <= (~^reg333);
              reg454 = $unsigned(reg330[(1'h0):(1'h0)]);
            end
        end
      else
        begin
          reg446 <= reg450;
        end
      for (forvar455 = (1'h0); (forvar455 < (1'h1)); forvar455 = (forvar455 + (1'h1)))
        begin
          if ($unsigned((reg357 ?
              reg359[(3'h5):(3'h5)] : $signed($signed(((8'ha3) ?
                  (7'h40) : reg326))))))
            begin
              reg456 <= (($signed(((reg413 < (8'hb9)) ?
                      (~^reg420) : forvar417)) ?
                  (8'ha4) : $signed($signed(reg454[(3'h6):(1'h1)]))) >= reg412);
              reg457 <= $unsigned(reg442[(2'h3):(2'h3)]);
              reg458 <= (((^~({reg448, wire385} ?
                      $unsigned(wire318) : (reg450 ~^ reg421))) ?
                  (((reg350 ? wire389 : reg432) ?
                      $unsigned(reg433) : (^reg422)) ^ reg443) : $unsigned($signed((wire387 - reg329)))) < (((^reg412[(2'h2):(1'h0)]) << forvar429[(4'h9):(4'h9)]) <<< (reg434 ?
                  forvar429 : $unsigned({(8'ha9), reg415}))));
            end
          else
            begin
              reg456 <= (~|{$unsigned($unsigned(reg433)),
                  reg325[(2'h3):(1'h0)]});
              reg457 <= reg393;
              reg459 = ($unsigned(reg417) ?
                  $signed(((|{reg383}) > $unsigned($signed(wire388)))) : reg427[(2'h2):(1'h0)]);
              reg460 = $unsigned(($unsigned((~&(|reg430))) ?
                  (reg396[(1'h0):(1'h0)] << ((wire385 ?
                      (8'hb1) : reg452) + (reg324 + reg333))) : reg452[(1'h1):(1'h0)]));
            end
          if ($signed(((&reg441) ?
              $signed(reg359[(4'hb):(3'h6)]) : $unsigned($signed($signed(reg349))))))
            begin
              reg461 = reg409;
            end
          else
            begin
              reg462 <= reg349;
              reg463 <= wire389[(4'hc):(1'h0)];
              reg464 <= (~^{(reg326 ? (reg445 & $signed(reg418)) : (-reg462)),
                  ($unsigned(reg344[(3'h5):(3'h5)]) && (&(reg422 ?
                      reg364 : reg411)))});
            end
          if ((^~{(~|(reg419 > reg379))}))
            begin
              reg465 <= wire385[(4'ha):(4'h8)];
              reg466 = {reg449[(3'h6):(2'h3)],
                  (!{{reg335[(4'ha):(1'h1)], (^~reg330)},
                      $signed((reg412 >> reg419))})};
            end
          else
            begin
              reg465 <= {$unsigned((-reg374))};
              reg467 <= ($signed((8'ha3)) ?
                  ((($unsigned((8'ha3)) ^ (reg439 * reg328)) ?
                      $unsigned($unsigned(reg350)) : (&$signed((8'ha0)))) ^ $signed(((reg402 >= wire386) ?
                      {reg423,
                          reg463} : (reg423 ^~ reg456)))) : (wire387[(3'h5):(1'h1)] || (&({reg325,
                          reg375} ?
                      (reg356 ? reg335 : reg416) : $signed(reg459)))));
              reg468 <= reg463[(2'h3):(2'h3)];
              reg469 = ((~reg441[(3'h4):(2'h2)]) ?
                  (&{(-reg456[(5'h12):(5'h11)])}) : reg402[(3'h6):(3'h6)]);
              reg470 <= reg379[(1'h0):(1'h0)];
            end
          for (forvar471 = (1'h0); (forvar471 < (2'h3)); forvar471 = (forvar471 + (1'h1)))
            begin
              reg472 <= (~&(($signed(reg452) != $unsigned((reg416 ?
                      reg444 : reg414))) ?
                  {(&$signed(reg426)),
                      reg359} : $unsigned((^(reg335 >> reg380)))));
              reg473 <= (wire387[(2'h2):(1'h0)] - ($signed({(8'ha0)}) ?
                  (8'ha7) : reg324));
            end
          for (forvar474 = (1'h0); (forvar474 < (2'h2)); forvar474 = (forvar474 + (1'h1)))
            begin
              reg475 = reg364;
              reg476 = {$signed($signed(((!reg438) == $signed(reg366)))),
                  reg430};
              reg477 <= ($signed((reg351 ?
                  $signed(reg351) : $unsigned((wire318 && (8'hba))))) || (!(((reg431 ?
                  reg433 : reg456) | reg403) >>> ((forvar471 ~^ reg426) <<< (wire318 >= reg364)))));
              reg478 = (-(|$signed((^(reg439 << reg432)))));
              reg479 <= reg434[(2'h2):(2'h2)];
            end
        end
    end
  assign wire480 = reg396[(2'h2):(2'h2)];
  assign wire481 = (reg368[(3'h5):(3'h5)] >> {reg422[(1'h0):(1'h0)]});
  always
    @(posedge clk) begin
      if ($unsigned(reg337))
        begin
          reg482 = (~&reg328[(4'hf):(4'hf)]);
          reg483 <= $signed({reg439});
        end
      else
        begin
          if ($unsigned(reg355))
            begin
              reg482 = $unsigned($unsigned(((!(reg467 <= reg403)) - ($unsigned(reg456) <<< reg397[(2'h2):(2'h2)]))));
              reg484 = (reg402 >> wire318[(4'ha):(3'h4)]);
              reg485 <= $signed($unsigned(reg473));
              reg486 <= wire480;
              reg487 <= $unsigned($unsigned({(^~reg477[(4'h8):(1'h0)])}));
            end
          else
            begin
              reg482 = $signed(((~(~|(reg357 && reg446))) >= $unsigned(reg439[(4'hf):(2'h2)])));
              reg483 <= ($unsigned($signed((+{reg356,
                  reg364}))) - $signed($signed((reg336 ?
                  reg394[(1'h1):(1'h0)] : (reg468 ^ reg431)))));
              reg485 <= reg359;
              reg486 <= (reg463 > $unsigned((!(+$signed(reg462)))));
            end
          reg488 <= (($signed($unsigned(wire389[(4'ha):(2'h3)])) != reg353[(1'h0):(1'h0)]) ?
              reg359[(3'h6):(3'h4)] : {reg438});
          if ((($unsigned(((^~(7'h41)) == reg351[(2'h3):(1'h1)])) ?
                  ((8'hb6) == ((reg401 ^ reg417) ?
                      reg484[(4'hc):(2'h2)] : reg416[(3'h5):(1'h0)])) : (&reg453[(1'h0):(1'h0)])) ?
              (~^((reg441[(3'h6):(2'h2)] ?
                  reg419 : {reg428}) >= reg357[(4'hc):(3'h4)])) : reg488))
            begin
              reg489 = reg418;
              reg490 = {((reg366[(2'h3):(2'h3)] ?
                      {(8'ha8),
                          (~|(8'hab))} : reg402[(3'h7):(3'h4)]) < $signed($unsigned(reg376)))};
            end
          else
            begin
              reg489 = (($unsigned($unsigned((wire319 * reg418))) ?
                  $unsigned({reg479[(1'h1):(1'h1)],
                      wire387}) : ((wire318 >> reg439) < ((reg462 ?
                      wire317 : (7'h44)) ^~ (~|reg484)))) >>> (reg473 ?
                  ((reg462[(3'h4):(2'h3)] ? (8'hbd) : $unsigned(reg470)) ?
                      (reg353 ^ $signed(reg376)) : wire318) : (~^$unsigned($signed(reg463)))));
              reg491 <= ($signed((((~reg402) ?
                      $unsigned(reg422) : $signed(reg374)) ?
                  reg356 : (+(^reg345)))) | {reg472[(3'h5):(1'h0)]});
            end
        end
      if ((((($signed(reg374) ^ $signed(reg413)) - (^~((7'h43) ?
              reg457 : reg326))) ?
          ($unsigned(reg472) ?
              (&(^reg413)) : $unsigned($unsigned((8'hbd)))) : reg353) << reg434[(4'hc):(3'h7)]))
        begin
          if ((|$unsigned({$signed(reg482[(4'h8):(2'h2)])})))
            begin
              reg492 <= $signed(reg490[(5'h11):(4'ha)]);
              reg493 = ($signed($unsigned($unsigned($unsigned((8'h9d))))) ~^ (~^(~&((reg439 ?
                  reg467 : (7'h41)) <= (~reg482)))));
              reg494 <= ((8'hb1) ?
                  {reg486[(2'h3):(2'h2)]} : (($unsigned({reg376, reg374}) ?
                      reg403 : reg489[(4'ha):(3'h4)]) < $unsigned({(reg351 < reg380)})));
              reg495 = $unsigned($signed($signed($unsigned($signed((8'hb5))))));
              reg496 = ($unsigned($unsigned((!(8'hbd)))) > (8'ha5));
            end
          else
            begin
              reg492 <= ($unsigned($signed(reg431)) ?
                  reg393[(3'h7):(1'h1)] : reg422[(2'h2):(2'h2)]);
            end
        end
      else
        begin
          reg493 = $unsigned((7'h41));
          if ($unsigned(wire387))
            begin
              reg494 <= (~|$signed(reg462[(1'h1):(1'h0)]));
              reg495 = reg337[(1'h1):(1'h1)];
              reg497 <= reg495[(4'h8):(1'h1)];
              reg498 = ({reg401[(2'h3):(1'h0)],
                      ((-$unsigned(reg410)) & {(^~reg351)})} ?
                  reg453[(2'h2):(2'h2)] : (reg456 ?
                      ((~^reg493[(1'h1):(1'h1)]) ?
                          ($signed((7'h40)) * reg491) : reg487[(2'h3):(2'h3)]) : $signed($unsigned((8'ha7)))));
              reg499 <= (+{(8'hb8), reg391[(1'h1):(1'h0)]});
            end
          else
            begin
              reg494 <= ($signed((~(^~(+reg391)))) ?
                  reg403[(5'h15):(4'hf)] : ($unsigned(reg493[(3'h6):(3'h4)]) ?
                      reg410[(1'h1):(1'h1)] : ((~^wire481) ?
                          ($unsigned(reg376) ?
                              reg485[(2'h2):(2'h2)] : (wire318 & (8'hb3))) : (wire321[(3'h5):(3'h4)] ?
                              ((8'hae) ?
                                  reg380 : wire389) : $unsigned(reg465)))));
              reg497 <= reg394;
              reg498 = reg391[(2'h2):(1'h1)];
              reg499 <= ((-(reg340 + reg493[(5'h11):(4'hb)])) ?
                  (8'ha9) : $unsigned(reg488));
            end
          for (forvar500 = (1'h0); (forvar500 < (2'h3)); forvar500 = (forvar500 + (1'h1)))
            begin
              reg501 = ((reg419 && $signed($unsigned((reg464 ?
                  reg351 : reg477)))) <= $signed($signed(reg416[(4'ha):(1'h1)])));
              reg502 <= reg366[(2'h2):(1'h1)];
              reg503 = ((|reg437[(2'h2):(1'h1)]) < $signed(reg410[(2'h3):(1'h0)]));
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed($unsigned($unsigned((reg497 ? (~&reg397) : (7'h41))))))
        begin
          if ((reg464 ? reg396[(1'h1):(1'h0)] : reg333[(1'h1):(1'h0)]))
            begin
              reg504 <= reg394[(3'h7):(3'h7)];
              reg505 = (reg325 ~^ $signed({$signed($signed(wire388)),
                  ((reg446 ~^ (8'hb7)) ? reg417[(3'h5):(1'h1)] : wire387)}));
              reg506 <= (^~(^($unsigned(reg353) ?
                  (^reg410[(2'h3):(1'h1)]) : ((reg457 ?
                      reg401 : reg344) ^~ reg344[(2'h3):(2'h3)]))));
            end
          else
            begin
              reg504 <= $signed((7'h40));
            end
          reg507 <= (+{$signed(((~|reg403) ? (&wire388) : reg344))});
        end
      else
        begin
          reg505 = $unsigned(wire386[(3'h5):(3'h5)]);
          if ((($unsigned((+((8'hab) ?
                  reg402 : reg468))) > $signed(reg343[(5'h10):(4'h8)])) ?
              ((({reg419, reg473} ?
                  {reg366} : (reg438 ? reg492 : reg430)) ^ ($unsigned(wire388) ?
                  (reg391 ?
                      reg418 : reg440) : reg494[(3'h5):(1'h1)])) - (((8'ha9) ?
                      $signed(reg499) : reg355) ?
                  ($signed(reg353) | $signed(reg343)) : $unsigned(reg507[(3'h4):(2'h3)]))) : wire385[(1'h0):(1'h0)]))
            begin
              reg506 <= reg473;
              reg508 = (((-({(8'hbf),
                      (8'h9c)} == $signed(reg413))) & $signed(reg507)) ?
                  (+$signed(reg462[(1'h0):(1'h0)])) : wire389);
              reg509 <= (~&$signed(reg356));
            end
          else
            begin
              reg508 = $signed(reg359);
            end
          if ($unsigned((~(reg416[(4'hb):(1'h1)] < ((reg468 ?
                  wire480 : (7'h42)) ?
              reg458 : {reg467})))))
            begin
              reg510 = $unsigned(reg336);
              reg511 <= ((&$unsigned($unsigned($signed((8'ha8))))) ?
                  $unsigned((8'hb4)) : (~|($signed($unsigned(reg374)) != reg494[(1'h0):(1'h0)])));
              reg512 <= ($unsigned(((((8'hb6) ?
                      reg368 : (7'h41)) ^~ reg401) << ((reg409 <= reg473) ?
                      (~reg397) : (reg479 ~^ reg453)))) ?
                  {reg374[(5'h11):(3'h5)],
                      $unsigned(reg337)} : $unsigned($unsigned($signed(wire320))));
            end
          else
            begin
              reg511 <= $unsigned({((^(~(8'hbe))) * reg437)});
              reg512 <= (wire321 ?
                  $signed($unsigned($signed(reg417))) : ((7'h40) ?
                      $unsigned((8'h9e)) : $signed($unsigned($signed(reg463)))));
              reg513 <= ((-reg437) > wire385);
              reg514 = ((((((8'hb6) ? reg437 : wire320) ?
                      ((8'haa) ? reg458 : (8'hb4)) : (reg344 ?
                          reg479 : reg402)) >> reg464) ?
                  {($signed(reg491) & {(8'hbb)})} : reg380) != $signed($signed(({reg437} || $signed(reg366)))));
            end
          for (forvar515 = (1'h0); (forvar515 < (3'h4)); forvar515 = (forvar515 + (1'h1)))
            begin
              reg516 = reg383;
            end
          if ($signed($unsigned($unsigned(reg336[(3'h5):(3'h5)]))))
            begin
              reg517 <= $signed((reg360 ?
                  (^~(reg361[(4'h9):(1'h0)] ?
                      (reg364 ?
                          reg479 : reg336) : reg345)) : $unsigned($unsigned((reg439 ?
                      reg509 : wire480)))));
              reg518 <= wire319;
              reg519 <= $signed(((reg337 && ((8'ha0) ?
                  reg506 : reg393[(1'h0):(1'h0)])) >= reg412));
            end
          else
            begin
              reg520 = reg399;
            end
        end
      if (reg456[(4'hd):(4'hd)])
        begin
          if (((7'h43) ?
              (((reg514[(4'ha):(4'h9)] ?
                      wire320 : $signed(reg330)) >>> (reg417[(3'h5):(3'h5)] + (reg360 ?
                      reg368 : reg510))) ?
                  ($unsigned((8'hb0)) ? {(~|reg391)} : {{reg505}}) : (-(reg349 ?
                      {reg375} : $signed(reg438)))) : $signed((~|wire321))))
            begin
              reg521 = $signed((reg417 ?
                  reg434[(4'hb):(4'h8)] : wire321[(2'h3):(2'h2)]));
              reg522 = reg499;
            end
          else
            begin
              reg521 = (reg418[(1'h1):(1'h1)] ? reg333 : (~^wire320));
              reg523 <= (((+(((8'hb5) ? reg399 : reg470) ?
                      (reg456 && reg368) : (reg393 || (8'ha2)))) ?
                  reg383[(3'h5):(2'h3)] : reg329[(2'h2):(2'h2)]) + $signed($unsigned($signed({reg324,
                  wire480}))));
              reg524 <= wire480[(3'h7):(3'h7)];
            end
          for (forvar525 = (1'h0); (forvar525 < (2'h3)); forvar525 = (forvar525 + (1'h1)))
            begin
              reg526 <= $unsigned($signed({$unsigned(reg439[(4'he):(4'hc)]),
                  ($signed(wire321) & (reg382 || reg522))}));
              reg527 = (($unsigned($unsigned((reg433 >> reg349))) <= {{(&reg376)},
                      reg446}) ?
                  (reg472 ?
                      reg409[(3'h7):(2'h3)] : $unsigned(((reg486 < reg523) * reg399))) : $unsigned($signed(reg353[(2'h3):(2'h2)])));
              reg528 <= (reg368[(2'h2):(1'h1)] ?
                  (^$unsigned((((8'haa) > wire481) ?
                      (~|reg517) : (reg417 ?
                          (8'ha6) : reg397)))) : $signed(($signed((reg463 ?
                          (8'hbf) : wire385)) ?
                      reg353 : $signed(reg512[(1'h0):(1'h0)]))));
              reg529 <= (8'hb8);
            end
          if ((reg436[(4'h8):(4'h8)] ?
              (reg439[(3'h6):(3'h4)] && $signed($unsigned((reg397 < forvar525)))) : $unsigned($signed(($unsigned(reg376) * $unsigned(reg462))))))
            begin
              reg530 <= ((^~$signed(wire319[(4'h8):(1'h1)])) ?
                  (~&$unsigned((reg440 ?
                      reg519[(3'h5):(1'h0)] : ((7'h44) > reg436)))) : reg360);
              reg531 <= reg379;
              reg532 <= $unsigned((8'hb9));
              reg533 = ($unsigned(reg456[(1'h1):(1'h1)]) ?
                  $unsigned(($unsigned({reg431,
                      reg355}) >>> (wire388[(1'h1):(1'h0)] ?
                      reg505[(4'hd):(2'h2)] : (8'ha4)))) : ($signed(reg441) ?
                      wire318 : reg446));
              reg534 = (reg532 ?
                  (reg527 <= reg522[(4'h8):(3'h5)]) : (reg510 == wire319[(4'ha):(3'h5)]));
            end
          else
            begin
              reg533 = $signed(wire321[(2'h2):(1'h1)]);
              reg534 = ($signed($unsigned(reg412[(2'h2):(1'h0)])) ?
                  $unsigned((8'hbe)) : $unsigned(reg413));
            end
          if ($signed(reg417[(1'h1):(1'h0)]))
            begin
              reg535 = $unsigned($unsigned((((&reg416) ?
                  (&reg512) : (!reg366)) ~^ ((reg479 ?
                  wire385 : reg477) | $signed(reg472)))));
              reg536 = ((reg430[(2'h2):(1'h1)] == reg437) >= (+($unsigned((reg446 <= reg505)) * ({reg330} << (reg505 >>> reg521)))));
            end
          else
            begin
              reg535 = $unsigned(reg356);
              reg537 <= (~&(~&$unsigned(((|reg513) + {reg393}))));
              reg538 <= reg326;
              reg539 = $signed((((reg380[(3'h4):(1'h0)] == {(8'h9d), reg467}) ?
                      reg465[(4'hc):(4'ha)] : (8'hb4)) ?
                  (&reg344) : reg413[(2'h3):(1'h0)]));
            end
          for (forvar540 = (1'h0); (forvar540 < (3'h4)); forvar540 = (forvar540 + (1'h1)))
            begin
              reg541 <= $signed((^~(|reg537[(3'h6):(1'h1)])));
            end
        end
      else
        begin
          if (($unsigned(((reg379[(4'h8):(3'h4)] && $signed(reg417)) ?
              reg456 : {$unsigned(reg412)})) && $unsigned(reg529)))
            begin
              reg523 <= (((~^reg375[(1'h1):(1'h0)]) ?
                      ({(^reg487), (reg518 > reg337)} ?
                          $signed(reg529[(3'h5):(2'h3)]) : reg497) : (+(^(~^reg414)))) ?
                  $unsigned((&{reg433,
                      $unsigned(reg533)})) : ({reg463[(1'h1):(1'h1)],
                      wire320[(2'h2):(1'h1)]} ^~ (($unsigned(reg439) == $signed((8'hb4))) ?
                      $unsigned({reg494, reg485}) : {((8'hbe) == reg328)})));
              reg525 = {(8'ha1), $unsigned(reg325[(2'h2):(2'h2)])};
            end
          else
            begin
              reg521 = ((reg337[(3'h5):(1'h0)] != $signed(reg430[(2'h2):(1'h1)])) - $unsigned($signed($signed($signed(forvar540)))));
              reg523 <= $unsigned(((reg465 <= (~^((8'hae) ?
                  wire320 : reg446))) ~^ {$unsigned({reg351, reg468})}));
            end
          if (((^($signed($unsigned(reg491)) != ((reg351 ?
                  (8'h9e) : (8'ha8)) != reg529))) ?
              $unsigned({reg324[(5'h11):(5'h11)],
                  ((reg492 && reg368) < $signed(reg494))}) : reg541))
            begin
              reg526 <= $signed($unsigned(reg528[(3'h7):(3'h6)]));
              reg527 = ((|reg328[(3'h5):(1'h1)]) != (8'hb8));
              reg528 <= $unsigned((-reg416));
              reg533 = reg436;
            end
          else
            begin
              reg526 <= (reg505[(4'he):(1'h0)] && reg457[(4'ha):(2'h3)]);
              reg528 <= (8'ha7);
              reg529 <= {({reg526} == reg440)};
              reg530 <= reg349;
            end
        end
      for (forvar542 = (1'h0); (forvar542 < (2'h3)); forvar542 = (forvar542 + (1'h1)))
        begin
          if (reg467)
            begin
              reg543 <= {(~^reg351[(3'h5):(3'h4)]),
                  ($unsigned(($unsigned(wire321) ?
                      reg530 : reg511)) || reg328)};
              reg544 <= {(!(~^$signed($unsigned(reg506))))};
            end
          else
            begin
              reg543 <= reg520[(1'h1):(1'h1)];
            end
          for (forvar545 = (1'h0); (forvar545 < (1'h0)); forvar545 = (forvar545 + (1'h1)))
            begin
              reg546 = ($signed((reg487 ?
                      {(reg470 ? reg491 : forvar542), (-reg541)} : ({(8'hbb),
                          reg533} - {reg462}))) ?
                  ((((reg465 ? (8'hb0) : reg488) ?
                          $signed(reg497) : (~|wire317)) ?
                      $unsigned(reg520) : reg399[(3'h7):(1'h1)]) >>> (&$signed(reg374))) : ((~^reg530[(3'h4):(3'h4)]) | (8'ha5)));
              reg547 = reg431[(4'hb):(4'h9)];
              reg548 <= (~^reg364[(1'h0):(1'h0)]);
              reg549 <= (&$signed((reg414 ?
                  ($signed(reg497) ^~ reg543[(1'h0):(1'h0)]) : reg328[(4'hb):(4'h8)])));
            end
          if (reg350[(2'h2):(1'h1)])
            begin
              reg550 <= reg546[(1'h0):(1'h0)];
              reg551 <= reg512[(2'h3):(1'h0)];
            end
          else
            begin
              reg550 <= ((~&$unsigned(($signed((8'hbd)) != reg403))) & {($signed({reg543}) ?
                      $unsigned(reg440) : (^(reg379 * reg462)))});
            end
          for (forvar552 = (1'h0); (forvar552 < (2'h3)); forvar552 = (forvar552 + (1'h1)))
            begin
              reg553 <= ((~|($signed($signed(reg350)) <= forvar542[(2'h2):(1'h1)])) ?
                  (^reg441[(4'hc):(3'h6)]) : wire480[(4'hb):(3'h6)]);
              reg554 <= reg412;
            end
        end
    end
  assign wire555 = ((reg488[(1'h1):(1'h1)] ?
                           (8'hbb) : $unsigned($signed((^~reg402)))) ?
                       ((reg437 ?
                           (+reg376[(1'h1):(1'h1)]) : wire389[(4'ha):(4'ha)]) || $unsigned((~|(wire318 ?
                           reg401 : reg343)))) : ($signed($signed({(8'h9f),
                           reg393})) ^~ (((reg528 * reg453) << (!(8'ha1))) ?
                           reg497[(1'h1):(1'h1)] : $unsigned($signed((8'ha9))))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module119  (y, clk, wire124, wire123, wire122, wire121, wire120);
  output wire [(32'h91a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire124;
  input wire signed [(5'h15):(1'h0)] wire123;
  input wire signed [(4'he):(1'h0)] wire122;
  input wire signed [(4'hb):(1'h0)] wire121;
  input wire [(5'h13):(1'h0)] wire120;
  wire [(5'h10):(1'h0)] wire248;
  wire signed [(4'h8):(1'h0)] wire247;
  wire [(5'h10):(1'h0)] wire246;
  wire signed [(2'h2):(1'h0)] wire245;
  wire signed [(5'h10):(1'h0)] wire207;
  wire signed [(3'h6):(1'h0)] wire206;
  wire [(5'h15):(1'h0)] wire205;
  wire signed [(3'h5):(1'h0)] wire204;
  wire signed [(4'ha):(1'h0)] wire127;
  wire signed [(4'he):(1'h0)] wire126;
  wire [(5'h13):(1'h0)] wire125;
  reg signed [(4'he):(1'h0)] reg312 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg310 = (1'h0);
  reg [(5'h10):(1'h0)] reg308 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg306 = (1'h0);
  reg signed [(4'he):(1'h0)] reg305 = (1'h0);
  reg [(4'hb):(1'h0)] reg303 = (1'h0);
  reg [(4'h8):(1'h0)] reg298 = (1'h0);
  reg signed [(4'he):(1'h0)] reg295 = (1'h0);
  reg [(3'h7):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg291 = (1'h0);
  reg [(2'h2):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg287 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg286 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg283 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg282 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg275 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg274 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg272 = (1'h0);
  reg [(3'h6):(1'h0)] reg269 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg268 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg264 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg260 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg259 = (1'h0);
  reg [(5'h10):(1'h0)] reg256 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg255 = (1'h0);
  reg [(5'h12):(1'h0)] reg254 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg244 = (1'h0);
  reg [(2'h2):(1'h0)] reg243 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg241 = (1'h0);
  reg [(3'h7):(1'h0)] reg240 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg239 = (1'h0);
  reg [(4'hf):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg235 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg231 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg225 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg224 = (1'h0);
  reg [(4'hc):(1'h0)] reg223 = (1'h0);
  reg [(3'h4):(1'h0)] reg222 = (1'h0);
  reg [(4'h9):(1'h0)] reg220 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg217 = (1'h0);
  reg [(4'h9):(1'h0)] reg213 = (1'h0);
  reg [(4'ha):(1'h0)] reg212 = (1'h0);
  reg [(5'h11):(1'h0)] reg210 = (1'h0);
  reg [(4'h8):(1'h0)] reg209 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg202 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg201 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg199 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg198 = (1'h0);
  reg [(5'h10):(1'h0)] reg197 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg195 = (1'h0);
  reg [(5'h14):(1'h0)] reg187 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg186 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg183 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg182 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg179 = (1'h0);
  reg [(3'h4):(1'h0)] reg157 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg175 = (1'h0);
  reg [(3'h6):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg167 = (1'h0);
  reg [(5'h11):(1'h0)] reg163 = (1'h0);
  reg [(2'h3):(1'h0)] reg162 = (1'h0);
  reg [(5'h12):(1'h0)] reg161 = (1'h0);
  reg [(2'h3):(1'h0)] reg160 = (1'h0);
  reg [(4'hb):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg158 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg155 = (1'h0);
  reg [(5'h14):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg141 = (1'h0);
  reg [(4'hf):(1'h0)] reg140 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg138 = (1'h0);
  reg [(4'hb):(1'h0)] reg137 = (1'h0);
  reg [(3'h6):(1'h0)] reg136 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg131 = (1'h0);
  reg [(5'h14):(1'h0)] reg129 = (1'h0);
  reg [(5'h13):(1'h0)] reg311 = (1'h0);
  reg [(2'h3):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg304 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg302 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg300 = (1'h0);
  reg [(4'h8):(1'h0)] reg299 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg297 = (1'h0);
  reg [(2'h2):(1'h0)] reg296 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg293 = (1'h0);
  reg [(4'hf):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg284 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg281 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg280 = (1'h0);
  reg [(5'h10):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar278 = (1'h0);
  reg [(4'hd):(1'h0)] reg277 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg276 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg271 = (1'h0);
  reg [(5'h14):(1'h0)] reg270 = (1'h0);
  reg [(3'h6):(1'h0)] reg267 = (1'h0);
  reg signed [(4'he):(1'h0)] reg265 = (1'h0);
  reg [(4'he):(1'h0)] reg263 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar258 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg [(5'h11):(1'h0)] forvar253 = (1'h0);
  reg [(5'h10):(1'h0)] reg252 = (1'h0);
  reg [(2'h2):(1'h0)] forvar251 = (1'h0);
  reg [(4'ha):(1'h0)] forvar249 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar239 = (1'h0);
  reg [(4'hd):(1'h0)] forvar242 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg237 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg236 = (1'h0);
  reg [(4'hd):(1'h0)] reg234 = (1'h0);
  reg [(3'h4):(1'h0)] reg233 = (1'h0);
  reg [(5'h11):(1'h0)] reg232 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg229 = (1'h0);
  reg signed [(4'he):(1'h0)] reg228 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg227 = (1'h0);
  reg [(4'hd):(1'h0)] reg226 = (1'h0);
  reg [(2'h2):(1'h0)] reg221 = (1'h0);
  reg [(3'h6):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg218 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg216 = (1'h0);
  reg [(4'hf):(1'h0)] reg215 = (1'h0);
  reg [(3'h5):(1'h0)] forvar214 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg211 = (1'h0);
  reg [(4'ha):(1'h0)] forvar208 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg203 = (1'h0);
  reg [(5'h11):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar196 = (1'h0);
  reg [(5'h12):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg193 = (1'h0);
  reg signed [(4'he):(1'h0)] reg192 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg191 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar190 = (1'h0);
  reg [(5'h10):(1'h0)] reg189 = (1'h0);
  reg [(4'hb):(1'h0)] reg188 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar185 = (1'h0);
  reg [(4'ha):(1'h0)] forvar184 = (1'h0);
  reg [(4'hf):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg180 = (1'h0);
  reg [(5'h13):(1'h0)] reg178 = (1'h0);
  reg [(4'h8):(1'h0)] forvar177 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg174 = (1'h0);
  reg [(4'hf):(1'h0)] reg173 = (1'h0);
  reg [(5'h14):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg170 = (1'h0);
  reg [(2'h3):(1'h0)] reg169 = (1'h0);
  reg [(5'h11):(1'h0)] reg166 = (1'h0);
  reg [(4'hf):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg164 = (1'h0);
  reg [(4'hf):(1'h0)] forvar157 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg156 = (1'h0);
  reg [(5'h13):(1'h0)] reg154 = (1'h0);
  reg [(5'h11):(1'h0)] reg152 = (1'h0);
  reg [(4'hd):(1'h0)] reg151 = (1'h0);
  reg [(4'ha):(1'h0)] reg150 = (1'h0);
  reg [(4'h9):(1'h0)] reg147 = (1'h0);
  reg [(4'hc):(1'h0)] reg146 = (1'h0);
  reg [(5'h11):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar143 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg142 = (1'h0);
  reg [(5'h14):(1'h0)] forvar135 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg139 = (1'h0);
  reg [(5'h14):(1'h0)] reg135 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg128 = (1'h0);
  assign y = {wire248,
                 wire247,
                 wire246,
                 wire245,
                 wire207,
                 wire206,
                 wire205,
                 wire204,
                 wire127,
                 wire126,
                 wire125,
                 reg312,
                 reg310,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg303,
                 reg298,
                 reg295,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg287,
                 reg286,
                 reg285,
                 reg283,
                 reg282,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg269,
                 reg268,
                 reg266,
                 reg264,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg256,
                 reg255,
                 reg254,
                 reg250,
                 reg244,
                 reg243,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg235,
                 reg231,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg220,
                 reg217,
                 reg213,
                 reg212,
                 reg210,
                 reg209,
                 reg202,
                 reg201,
                 reg199,
                 reg198,
                 reg197,
                 reg195,
                 reg187,
                 reg186,
                 reg183,
                 reg182,
                 reg179,
                 reg157,
                 reg176,
                 reg175,
                 reg171,
                 reg168,
                 reg167,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg155,
                 reg153,
                 reg149,
                 reg148,
                 reg141,
                 reg140,
                 reg138,
                 reg137,
                 reg136,
                 reg134,
                 reg133,
                 reg131,
                 reg129,
                 reg311,
                 reg309,
                 reg304,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg297,
                 reg296,
                 reg294,
                 reg293,
                 reg288,
                 reg284,
                 reg281,
                 reg280,
                 reg279,
                 forvar278,
                 reg277,
                 reg276,
                 reg271,
                 reg270,
                 reg267,
                 reg265,
                 reg263,
                 forvar258,
                 reg257,
                 forvar253,
                 reg252,
                 forvar251,
                 forvar249,
                 reg242,
                 forvar239,
                 forvar242,
                 reg237,
                 reg236,
                 reg234,
                 reg233,
                 reg232,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg221,
                 reg219,
                 reg218,
                 reg216,
                 reg215,
                 forvar214,
                 reg211,
                 forvar208,
                 reg203,
                 reg200,
                 forvar196,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 forvar190,
                 reg189,
                 reg188,
                 forvar185,
                 forvar184,
                 reg181,
                 reg180,
                 reg178,
                 forvar177,
                 reg174,
                 reg173,
                 reg172,
                 reg170,
                 reg169,
                 reg166,
                 reg165,
                 reg164,
                 forvar157,
                 reg156,
                 reg154,
                 reg152,
                 reg151,
                 reg150,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 forvar143,
                 reg142,
                 forvar135,
                 reg139,
                 reg135,
                 reg132,
                 reg130,
                 reg128,
                 (1'h0)};
  assign wire125 = $unsigned($signed(($signed(wire120[(5'h12):(3'h7)]) - $unsigned((wire124 ?
                       wire121 : wire123)))));
  assign wire126 = (wire123[(5'h11):(3'h7)] << (~|(!(|{wire123, wire122}))));
  assign wire127 = $signed((wire126 ^~ ((wire120 ?
                       {wire122} : wire124) + ((wire121 ? wire126 : wire123) ?
                       (wire122 != (8'hb3)) : wire123[(4'h9):(3'h4)]))));
  always
    @(posedge clk) begin
      if ((wire121[(4'h8):(3'h6)] == wire121))
        begin
          if ((((8'ha6) > wire122) || wire120[(4'he):(4'hb)]))
            begin
              reg128 = wire122;
              reg129 <= ($signed(wire124) ?
                  $signed($unsigned((~&(wire120 ^ wire123)))) : (($signed(wire120[(3'h6):(1'h1)]) ?
                      wire124[(3'h4):(2'h2)] : (wire123 != wire121[(4'ha):(4'ha)])) - $unsigned($unsigned(wire122[(2'h2):(2'h2)]))));
              reg130 = {(^((^~(~wire127)) & {$unsigned((8'hb6)),
                      $signed(reg128)})),
                  reg129[(4'ha):(1'h0)]};
              reg131 <= $signed($unsigned((&$unsigned((^wire124)))));
            end
          else
            begin
              reg129 <= $unsigned($signed($signed($unsigned(reg131))));
              reg131 <= ((~^$unsigned(($signed(wire121) <<< $signed(wire125)))) ?
                  ($signed(wire126) ?
                      (!((wire122 - (8'ha3)) ?
                          $unsigned(wire123) : (~&reg128))) : ((8'hba) ?
                          $unsigned(reg129[(4'h8):(1'h1)]) : (^(wire125 ?
                              reg131 : wire123)))) : ($signed(($unsigned((8'hb6)) >= $signed(wire120))) ?
                      ($signed((wire121 ? wire124 : reg131)) ?
                          $unsigned($signed(reg129)) : {$unsigned((8'ha8))}) : $unsigned(($unsigned(wire120) ?
                          $unsigned((8'ha8)) : $unsigned((7'h42))))));
              reg132 = ($unsigned(wire124[(3'h6):(1'h0)]) ?
                  ((-{(8'hb1)}) ^ (wire127[(4'h8):(2'h2)] <= (reg130 ?
                      (wire120 ? reg130 : wire124) : (wire122 ?
                          reg129 : reg130)))) : (wire125[(4'h9):(3'h7)] <<< ($signed((8'hba)) ?
                      wire121[(2'h2):(1'h1)] : $unsigned((8'haa)))));
              reg133 <= wire126;
              reg134 <= ((&$unsigned($signed(wire121))) ?
                  wire121[(4'hb):(2'h3)] : wire122[(4'hd):(4'h8)]);
            end
          if ($signed($signed(reg134)))
            begin
              reg135 = ($signed((~&$unsigned($unsigned(reg132)))) ?
                  $unsigned($unsigned(reg129)) : (^$signed(((reg131 ?
                          wire120 : reg134) ?
                      {(7'h40), wire120} : $signed(reg134)))));
              reg136 <= reg132[(3'h6):(1'h0)];
              reg137 <= {reg131[(5'h14):(4'hd)]};
              reg138 <= (8'ha4);
            end
          else
            begin
              reg136 <= ((reg129[(1'h0):(1'h0)] ?
                      wire125[(4'hd):(4'ha)] : $signed(wire127)) ?
                  (8'ha2) : (~reg134));
              reg137 <= reg132;
              reg139 = reg138[(4'hd):(4'ha)];
              reg140 <= reg128;
              reg141 <= $signed($signed((($signed(reg133) & (reg128 ?
                      reg134 : wire127)) ?
                  ((wire123 > reg131) <<< (~^wire121)) : reg134)));
            end
        end
      else
        begin
          if (reg130[(4'hf):(1'h1)])
            begin
              reg128 = reg140;
              reg130 = reg133[(2'h2):(1'h0)];
              reg132 = (wire120 ?
                  $signed($unsigned((8'h9c))) : $unsigned($signed($signed(reg131))));
            end
          else
            begin
              reg128 = (($signed((reg132[(1'h1):(1'h0)] ?
                      (reg140 > reg141) : {(7'h43)})) + (^($unsigned(reg133) ?
                      $signed(wire121) : (&wire121)))) ?
                  (^$signed($signed(wire122[(4'h9):(4'h8)]))) : ($signed(({reg134,
                              reg134} ?
                          $unsigned(reg134) : (reg130 ^ reg139))) ?
                      $unsigned(reg133[(1'h0):(1'h0)]) : ((((8'ha9) ?
                                  reg140 : (8'haf)) ?
                              {reg136} : $unsigned(wire122)) ?
                          $unsigned((reg128 ^ reg138)) : reg132[(1'h0):(1'h0)])));
              reg129 <= {(|({wire122} * ({reg128,
                      reg128} > $signed(wire121))))};
              reg130 = ($unsigned((+reg135)) ?
                  (($unsigned($signed(wire124)) <= $unsigned((reg136 ?
                      reg130 : wire124))) == wire122) : reg128);
              reg131 <= $unsigned($signed($signed((reg141[(5'h14):(5'h13)] < (reg134 ?
                  wire126 : reg134)))));
              reg133 <= reg130[(1'h0):(1'h0)];
            end
          reg134 <= reg133[(3'h4):(1'h0)];
          for (forvar135 = (1'h0); (forvar135 < (2'h3)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= wire126;
            end
          if (reg131[(5'h14):(2'h2)])
            begin
              reg137 <= ($unsigned(($unsigned(((8'h9d) >= wire120)) - (&$unsigned(reg140)))) ?
                  (reg132 >> reg132[(3'h4):(2'h2)]) : $unsigned(reg137[(4'h9):(3'h5)]));
            end
          else
            begin
              reg137 <= (8'hb9);
              reg138 <= $signed($unsigned((~^(8'ha4))));
            end
          if ($signed($unsigned({$unsigned((reg136 ? wire125 : wire120))})))
            begin
              reg139 = (-reg141);
              reg140 <= forvar135;
              reg142 = {reg131};
            end
          else
            begin
              reg139 = (~|$signed(reg141));
            end
        end
      if ($unsigned(reg137))
        begin
          for (forvar143 = (1'h0); (forvar143 < (1'h1)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg144 = (7'h40);
              reg145 = {(^~reg130),
                  $signed(($unsigned({wire127, reg128}) ?
                      ((8'hb3) <= $signed((8'ha7))) : reg140[(2'h2):(1'h0)]))};
              reg146 = ((!$unsigned($unsigned($unsigned(reg137)))) != $signed(forvar135));
              reg147 = forvar135[(5'h11):(3'h6)];
              reg148 <= $unsigned(((!$signed(reg147[(3'h5):(1'h0)])) ?
                  (~&(~|(~^(8'hb0)))) : ((~^$signed(reg133)) ^~ $signed($signed(reg137)))));
            end
        end
      else
        begin
          for (forvar143 = (1'h0); (forvar143 < (2'h3)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg144 = reg142[(4'hb):(2'h3)];
              reg148 <= ($signed(reg147[(1'h0):(1'h0)]) != reg146);
              reg149 <= reg146;
              reg150 = reg132;
              reg151 = ({(!((wire121 << reg150) ?
                          (^forvar143) : reg133[(2'h2):(2'h2)])),
                      $signed($unsigned((reg148 ? (8'hae) : (7'h42))))} ?
                  {(((reg148 ?
                          forvar135 : reg149) ^~ reg129[(3'h5):(3'h4)]) <<< reg137[(2'h3):(2'h3)])} : forvar143);
            end
          if (({$unsigned($unsigned(wire125[(2'h3):(1'h0)])),
                  (forvar143 == ($signed(reg149) ?
                      {reg136} : reg139[(1'h0):(1'h0)]))} ?
              ($unsigned((wire127[(3'h6):(2'h3)] ?
                      ((8'ha9) <<< (8'hac)) : (reg137 - reg136))) ?
                  (|$unsigned({wire122, reg145})) : reg138) : (~&reg131)))
            begin
              reg152 = reg135[(3'h7):(3'h7)];
              reg153 <= $signed(($signed(reg128) + (reg142[(4'hb):(1'h1)] == ((~|wire125) ?
                  wire125[(5'h13):(3'h5)] : $unsigned(reg132)))));
            end
          else
            begin
              reg153 <= (reg134 ?
                  (reg141[(3'h4):(1'h1)] ?
                      reg130[(3'h7):(3'h5)] : reg136[(2'h3):(1'h1)]) : reg147);
              reg154 = reg135[(3'h7):(3'h4)];
              reg155 <= {{(~&$unsigned(wire124[(4'h8):(3'h4)])),
                      $signed($unsigned(reg140))},
                  $signed((reg150 ^~ wire127))};
            end
        end
      if (((~^($signed((reg145 ? wire120 : reg139)) ?
              reg144 : reg131[(4'ha):(3'h4)])) ?
          (~|($signed($signed(reg144)) ?
              (((8'hbb) ?
                  wire121 : wire122) < {reg147}) : (~&((8'hb2) >= wire120)))) : {forvar143[(4'hf):(4'h9)]}))
        begin
          reg156 = ($signed({reg136}) ?
              (~|reg139[(2'h2):(1'h1)]) : (reg129 == (8'ha2)));
          for (forvar157 = (1'h0); (forvar157 < (3'h4)); forvar157 = (forvar157 + (1'h1)))
            begin
              reg158 <= ($unsigned(reg155) ?
                  $unsigned(((reg135 && {reg134}) ?
                      reg142 : wire123)) : (wire126 ?
                      $signed((((8'hb8) ? wire123 : (8'ha6)) ?
                          reg136 : $signed(forvar157))) : {reg145[(4'h8):(2'h3)]}));
            end
          if ($unsigned(($signed(((wire123 ? reg145 : reg142) ?
              $signed(wire122) : $unsigned(wire123))) * reg131[(4'h8):(2'h2)])))
            begin
              reg159 <= {reg135,
                  {wire123[(4'he):(3'h4)],
                      ((8'h9f) ? reg139 : {reg134[(3'h4):(1'h0)], reg158})}};
              reg160 <= $signed({reg141});
              reg161 <= (reg146 >>> (8'hbd));
              reg162 <= forvar135;
              reg163 <= reg155[(1'h0):(1'h0)];
            end
          else
            begin
              reg164 = (!(^~$signed(((reg163 >= reg155) ?
                  $unsigned(reg137) : {wire120}))));
              reg165 = $unsigned(wire122);
            end
          if (((8'hb2) << wire120[(5'h11):(4'hc)]))
            begin
              reg166 = $signed(((($unsigned(reg158) << $unsigned((8'hb3))) || reg138[(4'hb):(4'h9)]) ?
                  ($unsigned(reg158[(4'hb):(3'h5)]) <= wire120) : wire127));
              reg167 <= (~|(!((8'hbb) ^~ $signed($signed((8'hb2))))));
              reg168 <= (reg158[(1'h0):(1'h0)] << ((+$unsigned($unsigned(reg156))) ?
                  $signed((^~(reg151 ^~ reg130))) : $unsigned(reg152)));
              reg169 = ((~reg156[(2'h2):(1'h0)]) ?
                  wire127[(3'h4):(3'h4)] : reg167);
              reg170 = reg154[(4'hd):(4'ha)];
            end
          else
            begin
              reg167 <= $unsigned(({($signed(reg128) ~^ (~reg147))} >>> $unsigned(reg155[(2'h2):(1'h1)])));
              reg168 <= ((wire120 > ($signed((!reg146)) << $signed((reg155 > reg139)))) ?
                  (&{(^((8'hb9) >>> reg155))}) : {$unsigned($unsigned($unsigned(reg164)))});
              reg169 = (+forvar135);
              reg171 <= {($unsigned((reg130[(5'h11):(3'h4)] >>> $signed(wire126))) <= reg153)};
            end
          if (($unsigned(forvar143[(4'ha):(2'h3)]) >> $signed(reg149[(1'h0):(1'h0)])))
            begin
              reg172 = $unsigned(reg155);
              reg173 = reg137;
              reg174 = $signed((~&(8'ha3)));
            end
          else
            begin
              reg172 = {$signed($signed((^(^reg171)))),
                  (($signed({reg160}) ?
                          wire121 : $unsigned(reg130[(3'h7):(3'h4)])) ?
                      ((reg136 - ((8'ha9) ^ reg169)) >>> (+$unsigned(reg139))) : reg155)};
              reg175 <= (($unsigned((((8'hb8) ^~ (8'ha9)) ?
                          (^(8'hb9)) : reg158[(5'h12):(4'ha)])) ?
                      reg128 : $unsigned(reg162[(2'h3):(2'h2)])) ?
                  $signed(reg139[(4'ha):(1'h1)]) : (^~(8'hb6)));
              reg176 <= (^$signed({reg164, $unsigned((wire127 <<< reg146))}));
            end
        end
      else
        begin
          if ((8'ha3))
            begin
              reg157 <= {((&$signed((forvar157 ? wire120 : reg165))) ?
                      reg152 : (($signed(reg144) ?
                          {reg140,
                              reg136} : wire122[(4'ha):(3'h7)]) || ({reg139} ?
                          (reg142 ? reg132 : reg154) : $unsigned(reg164)))),
                  (wire125[(4'hc):(3'h7)] ?
                      ((-reg152) != ((+(8'hbb)) ?
                          $unsigned(wire127) : (reg133 || reg161))) : {(+{reg131,
                              reg152}),
                          $unsigned((^~reg145))})};
              reg158 <= (((reg159 * (reg141 ?
                      $unsigned((8'hab)) : wire120)) + $signed(reg134)) ?
                  ($signed($signed((~(8'ha2)))) < (^((reg144 ^ reg164) || (reg142 ?
                      reg132 : reg171)))) : reg150[(4'h8):(3'h5)]);
              reg159 <= ((wire121[(3'h4):(1'h1)] * ({$unsigned(reg129)} ?
                  (~^$signed(reg165)) : (wire123 || (~|(8'hac))))) * (((~|(reg145 >= reg167)) ?
                  $signed((reg169 - reg167)) : wire125) && reg133));
              reg164 = reg172;
              reg167 <= $signed((&(wire121[(1'h0):(1'h0)] ?
                  (forvar143 != (~reg138)) : reg140[(4'he):(2'h2)])));
            end
          else
            begin
              reg156 = ((~^(reg164 ?
                  reg133 : {reg150[(4'h8):(3'h6)]})) | (reg129[(3'h4):(2'h3)] ?
                  $unsigned($signed((reg153 ?
                      reg167 : reg174))) : wire122[(2'h3):(2'h3)]));
            end
          if ((~{(reg135[(4'h8):(2'h2)] & (~{forvar135}))}))
            begin
              reg169 = (({((!forvar143) == wire125[(1'h1):(1'h0)])} && ($signed((+reg176)) * $signed((reg149 != reg154)))) << (wire120[(5'h10):(3'h4)] >= {($signed(reg162) <<< (wire124 && wire124))}));
              reg170 = (({forvar143[(4'ha):(4'ha)]} + (^((reg137 ?
                          (8'hb8) : wire123) ?
                      (reg160 < reg162) : $unsigned(reg147)))) ?
                  $unsigned(forvar135) : $signed(reg172[(3'h4):(2'h2)]));
              reg172 = $signed($signed($signed($signed((~|wire123)))));
              reg175 <= $unsigned(reg158[(4'hd):(3'h4)]);
              reg176 <= (reg144[(4'hd):(4'h8)] ?
                  reg129 : ((wire121[(4'h8):(2'h2)] * $signed((reg150 + reg173))) ?
                      $unsigned((reg139[(4'hc):(1'h1)] ^~ (~&(8'ha6)))) : (reg166[(4'ha):(2'h3)] >>> ({reg166} ?
                          reg137[(4'hb):(4'h8)] : (reg148 ?
                              reg156 : reg158)))));
            end
          else
            begin
              reg169 = (~&($signed({reg152[(4'hf):(3'h6)],
                      reg164[(4'hf):(3'h5)]}) ?
                  (^reg130[(4'hb):(4'ha)]) : reg159[(4'hb):(3'h6)]));
              reg171 <= $signed((reg137[(4'h9):(4'h9)] >>> {(reg150[(4'ha):(2'h3)] ~^ $signed(reg140)),
                  $signed(reg141[(1'h1):(1'h0)])}));
              reg175 <= wire121;
            end
          for (forvar177 = (1'h0); (forvar177 < (2'h3)); forvar177 = (forvar177 + (1'h1)))
            begin
              reg178 = (reg148 ^ ($signed((^reg149[(2'h3):(1'h1)])) ?
                  ((~(reg132 ? forvar135 : reg161)) ?
                      (((8'hb4) != (8'ha9)) ?
                          reg153[(4'ha):(4'ha)] : {reg133}) : ((reg174 >> forvar135) ^ (~|reg149))) : {$signed({forvar143,
                          reg161})}));
              reg179 <= (((^(forvar143[(3'h6):(2'h2)] ?
                      $signed(reg158) : $signed(reg154))) ?
                  $unsigned($unsigned(((8'ha4) ? reg133 : reg152))) : {({reg132,
                              reg151} ?
                          $unsigned(reg131) : $signed(reg163)),
                      (+{wire122})}) != {reg156, (&reg162)});
              reg180 = ($unsigned((~&($unsigned(reg139) ?
                  $signed(reg137) : ((8'ha0) ? reg167 : (8'ha9))))) || reg155);
            end
          if ((&reg141))
            begin
              reg181 = forvar157[(4'ha):(3'h6)];
            end
          else
            begin
              reg182 <= (&$unsigned(((8'hb1) != ((reg139 | reg162) ?
                  (~&reg164) : $signed(wire126)))));
              reg183 <= $unsigned((^wire123[(4'h8):(1'h0)]));
            end
        end
      for (forvar184 = (1'h0); (forvar184 < (3'h4)); forvar184 = (forvar184 + (1'h1)))
        begin
          for (forvar185 = (1'h0); (forvar185 < (2'h3)); forvar185 = (forvar185 + (1'h1)))
            begin
              reg186 <= $unsigned($unsigned(wire125[(2'h2):(1'h0)]));
              reg187 <= $signed(reg168[(4'h8):(1'h0)]);
              reg188 = wire122[(4'hb):(2'h3)];
              reg189 = reg146[(4'hb):(3'h4)];
            end
        end
      for (forvar190 = (1'h0); (forvar190 < (2'h2)); forvar190 = (forvar190 + (1'h1)))
        begin
          if (reg130)
            begin
              reg191 = (((-{wire121}) ~^ $unsigned({forvar177[(3'h6):(2'h2)],
                      (reg153 >>> reg179)})) ?
                  ($signed(reg154[(5'h11):(4'h8)]) - (-reg159)) : (~&reg128));
              reg192 = (~&(^reg176));
              reg193 = (~|(!(~^(reg131[(1'h0):(1'h0)] ?
                  $signed(reg170) : ((8'hbb) > reg138)))));
            end
          else
            begin
              reg191 = reg170;
              reg192 = $signed((~^(8'ha5)));
              reg193 = $unsigned(forvar143[(4'h9):(3'h7)]);
              reg194 = $unsigned(reg135);
              reg195 <= $unsigned(($signed($unsigned({(8'hb8),
                  wire121})) + $unsigned(($signed((8'h9f)) ^~ reg180[(3'h7):(2'h3)]))));
            end
          for (forvar196 = (1'h0); (forvar196 < (2'h3)); forvar196 = (forvar196 + (1'h1)))
            begin
              reg197 <= $signed({$signed($signed($signed(reg164))),
                  (+(((8'ha4) ? reg133 : wire125) ~^ (reg128 < reg132)))});
            end
          if ((({({(8'ha8), reg131} ? {reg161, reg132} : {reg144}),
                      {reg136[(1'h1):(1'h0)], ((8'hac) >>> wire121)}} ?
                  (reg158[(5'h11):(4'hf)] >> (!(&forvar184))) : reg181) ?
              (+(+forvar185)) : $unsigned(((~|forvar190) ^ $signed($unsigned(reg168))))))
            begin
              reg198 <= (reg159[(2'h3):(1'h0)] ?
                  (reg146 != (+$signed(reg142[(4'hb):(2'h2)]))) : $unsigned(reg169[(2'h2):(1'h0)]));
            end
          else
            begin
              reg198 <= (~reg188[(1'h1):(1'h0)]);
            end
          if ((8'hab))
            begin
              reg199 <= $signed($unsigned($unsigned((|(forvar143 ~^ reg146)))));
            end
          else
            begin
              reg200 = reg199[(3'h4):(1'h0)];
              reg201 <= reg161[(4'ha):(4'ha)];
              reg202 <= (!($unsigned({{(8'ha4), reg167},
                  (forvar196 && (8'hb3))}) < reg188[(4'hb):(3'h7)]));
              reg203 = reg132;
            end
        end
    end
  assign wire204 = reg136[(2'h3):(1'h0)];
  assign wire205 = (|$unsigned(((reg134 ^~ $signed(wire120)) || $signed($unsigned(reg160)))));
  assign wire206 = ($signed((reg136[(1'h0):(1'h0)] << {$signed(wire123)})) ?
                       $signed($signed(wire123)) : (($unsigned((^~reg138)) ?
                               (8'ha4) : ($unsigned((8'hac)) == $unsigned(wire127))) ?
                           (-(wire204 ?
                               $signed(reg198) : {reg182})) : reg168[(4'h8):(3'h5)]));
  assign wire207 = ($unsigned(wire124[(2'h3):(1'h1)]) != reg148);
  always
    @(posedge clk) begin
      for (forvar208 = (1'h0); (forvar208 < (1'h1)); forvar208 = (forvar208 + (1'h1)))
        begin
          if (reg167)
            begin
              reg209 <= (wire121 ?
                  (reg137 ?
                      (!(|forvar208)) : ($unsigned((~|forvar208)) ?
                          reg182 : {{(7'h42)}})) : $unsigned($unsigned($unsigned(wire122[(4'h9):(4'h9)]))));
              reg210 <= reg136[(3'h6):(3'h4)];
              reg211 = $signed(reg137);
            end
          else
            begin
              reg209 <= $signed(((forvar208[(1'h0):(1'h0)] ?
                  (reg137[(4'h8):(3'h5)] - $signed(reg209)) : ($signed(wire126) | reg158[(2'h2):(1'h0)])) ^~ (wire206[(3'h6):(2'h3)] ?
                  (~^$signed(reg141)) : reg197[(4'he):(3'h5)])));
              reg211 = wire206;
              reg212 <= reg197[(5'h10):(4'hd)];
            end
          reg213 <= (^~(^{(wire125[(1'h1):(1'h0)] ? reg186 : (~&reg159))}));
          for (forvar214 = (1'h0); (forvar214 < (3'h4)); forvar214 = (forvar214 + (1'h1)))
            begin
              reg215 = $signed($signed($unsigned((reg183 ?
                  $unsigned(wire124) : (reg187 ~^ reg157)))));
              reg216 = ((-{$unsigned(wire124[(2'h3):(1'h0)])}) == $unsigned((((forvar208 ^~ reg167) ?
                  reg134 : reg202[(1'h0):(1'h0)]) | reg201)));
              reg217 <= reg131;
              reg218 = (!($signed(reg195[(2'h3):(2'h2)]) ?
                  (!$unsigned($signed(forvar208))) : wire206));
            end
          reg219 = wire127;
        end
      if ({$signed(reg183[(4'h8):(1'h1)]),
          ((~^(~$signed(reg182))) != $signed($signed((~&reg215))))})
        begin
          if ((reg155[(4'h8):(4'h8)] * reg219[(1'h0):(1'h0)]))
            begin
              reg220 <= $unsigned($signed((&((wire122 ?
                  wire127 : reg218) == {(7'h43), reg131}))));
              reg221 = reg212;
            end
          else
            begin
              reg221 = ($unsigned($signed(wire125[(3'h7):(1'h1)])) ?
                  (((~|reg182[(1'h0):(1'h0)]) ?
                      (reg133 <= reg155[(3'h6):(1'h1)]) : forvar214) | (wire123 - $unsigned((forvar214 ?
                      reg168 : reg153)))) : $signed(((!wire123[(4'hf):(3'h4)]) >>> (8'hbd))));
              reg222 <= $unsigned($signed($unsigned($unsigned((-reg157)))));
              reg223 <= $signed((reg221[(2'h2):(2'h2)] ? {reg136} : reg148));
              reg224 <= (reg216 >>> (($signed(reg175) >>> (((8'ha9) * reg148) ?
                      $unsigned(reg131) : reg218)) ?
                  reg161 : $unsigned($signed(reg134[(1'h1):(1'h0)]))));
              reg225 <= {$unsigned($unsigned($signed(reg157[(1'h0):(1'h0)])))};
            end
        end
      else
        begin
          if ({(8'had)})
            begin
              reg220 <= $signed($signed((((reg129 | reg186) && (~reg134)) ?
                  $signed($unsigned((8'hb7))) : $unsigned(reg138))));
            end
          else
            begin
              reg221 = reg157[(2'h2):(1'h1)];
              reg222 <= (($signed(((~reg137) && reg175)) ^ reg199[(1'h1):(1'h1)]) ?
                  $signed($signed(reg138[(4'h9):(1'h0)])) : reg158);
              reg226 = reg209[(3'h4):(2'h2)];
              reg227 = {reg223};
              reg228 = reg149;
            end
          reg229 = reg220;
          if ((~^$signed(reg162)))
            begin
              reg230 = $signed($unsigned($unsigned($unsigned($unsigned(reg201)))));
              reg231 <= $signed({(~^(~|reg158))});
            end
          else
            begin
              reg231 <= forvar214;
              reg232 = wire206;
              reg233 = reg160[(2'h2):(1'h1)];
              reg234 = (+(|reg219));
              reg235 <= ((~|reg215[(4'hd):(3'h7)]) ?
                  (8'hb7) : reg155[(4'ha):(3'h6)]);
            end
          reg236 = reg131[(4'ha):(1'h0)];
          reg237 = (~|$unsigned((~wire124[(3'h5):(3'h4)])));
        end
      if (reg225)
        begin
          if (reg133)
            begin
              reg238 <= $unsigned((^$signed(reg224)));
              reg239 <= $unsigned(wire206[(1'h1):(1'h1)]);
              reg240 <= {wire207};
            end
          else
            begin
              reg238 <= reg212;
              reg239 <= (8'hb7);
            end
          reg241 <= (8'hb8);
          for (forvar242 = (1'h0); (forvar242 < (2'h3)); forvar242 = (forvar242 + (1'h1)))
            begin
              reg243 <= $unsigned(($signed(reg234) ?
                  $signed(({(8'ha9), (8'ha2)} ?
                      reg237[(4'h8):(1'h0)] : reg215)) : $signed(($signed((8'ha1)) || reg241[(2'h2):(1'h0)]))));
              reg244 <= ($unsigned($signed((+(reg240 ? reg223 : reg148)))) ?
                  reg237[(3'h7):(3'h4)] : $unsigned((&$signed($signed(reg226)))));
            end
        end
      else
        begin
          reg238 <= reg133;
          for (forvar239 = (1'h0); (forvar239 < (3'h4)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg242 = $signed(reg158);
            end
        end
    end
  assign wire245 = (8'hab);
  assign wire246 = reg238;
  assign wire247 = (reg198[(4'h8):(4'h8)] ? reg171 : wire123[(5'h12):(2'h2)]);
  assign wire248 = {reg155,
                       ({reg224} ?
                           {wire245[(1'h1):(1'h0)]} : $unsigned(({wire205} ~^ $signed(reg136))))};
  always
    @(posedge clk) begin
      for (forvar249 = (1'h0); (forvar249 < (2'h2)); forvar249 = (forvar249 + (1'h1)))
        begin
          reg250 <= (~&$signed((reg138[(3'h7):(1'h0)] ^ $unsigned(((8'hbe) ?
              reg133 : (8'ha6))))));
          for (forvar251 = (1'h0); (forvar251 < (1'h0)); forvar251 = (forvar251 + (1'h1)))
            begin
              reg252 = ((~|(^($signed(forvar251) < (~|reg138)))) ?
                  $signed(((~&$signed(reg210)) ?
                      reg186[(1'h0):(1'h0)] : reg224[(3'h6):(3'h5)])) : ($unsigned((((8'ha1) ?
                              reg235 : (8'hb8)) ?
                          ((8'ha7) - reg158) : (+reg199))) ?
                      (((^~reg129) >>> (8'hb4)) ?
                          ((reg183 ?
                              reg157 : reg168) ^ reg158) : {(reg129 & forvar249),
                              reg186[(2'h3):(1'h0)]}) : reg159));
            end
        end
      for (forvar253 = (1'h0); (forvar253 < (1'h1)); forvar253 = (forvar253 + (1'h1)))
        begin
          if ($signed($signed($signed($unsigned((^reg141))))))
            begin
              reg254 <= ($signed($signed({$signed((8'ha2))})) == (wire122 ?
                  reg171[(2'h2):(1'h0)] : reg161[(3'h4):(2'h2)]));
              reg255 <= $signed(((reg137[(1'h0):(1'h0)] ? (8'hae) : wire248) ?
                  wire205[(5'h14):(4'hf)] : reg195));
              reg256 <= reg157;
            end
          else
            begin
              reg257 = $signed($unsigned(($unsigned(reg176) ?
                  reg141[(4'hc):(4'hc)] : (reg197[(3'h6):(2'h3)] - ((8'h9f) & wire122)))));
            end
          for (forvar258 = (1'h0); (forvar258 < (2'h3)); forvar258 = (forvar258 + (1'h1)))
            begin
              reg259 <= $unsigned(wire204[(2'h2):(1'h0)]);
              reg260 <= reg160;
              reg261 <= $unsigned({$unsigned(reg240)});
              reg262 <= reg197;
              reg263 = ((~(((reg140 ? reg231 : reg168) ?
                  (wire121 && forvar251) : reg201[(1'h0):(1'h0)]) ~^ $signed($signed(reg213)))) >>> ({$signed({reg157,
                          (8'haa)})} ?
                  wire247[(3'h4):(1'h1)] : reg202[(4'ha):(1'h0)]));
            end
          if ((~|$signed(reg217)))
            begin
              reg264 <= wire207;
              reg265 = reg131[(5'h13):(4'hf)];
              reg266 <= (~&($unsigned($unsigned(reg159[(3'h5):(3'h5)])) ?
                  ((~|(wire123 - reg186)) ?
                      {$unsigned((8'ha3)),
                          (~|reg213)} : ($unsigned((8'ha2)) ~^ (reg212 ~^ reg209))) : (~reg160[(2'h3):(1'h1)])));
              reg267 = reg161[(3'h7):(3'h4)];
            end
          else
            begin
              reg264 <= $signed(((forvar251 ^ ($signed(reg149) ?
                      (reg197 ~^ (8'hae)) : (^reg217))) ?
                  reg198 : reg250[(4'h9):(3'h6)]));
              reg266 <= {$unsigned($signed(($signed(reg133) ?
                      (~&reg266) : reg240))),
                  $signed(((reg179 ?
                      $unsigned(reg157) : forvar258) || $signed(((8'hb6) >= (8'hb1)))))};
            end
          if ((|$signed($signed((reg167 <= reg212)))))
            begin
              reg268 <= $signed($signed(reg263));
              reg269 <= (~($signed($signed({reg153})) ?
                  reg186[(1'h0):(1'h0)] : {($unsigned((8'hab)) && (reg235 ?
                          (7'h42) : reg223)),
                      forvar249}));
              reg270 = ({(8'hb9)} ? wire124 : $signed(reg265[(4'h9):(4'h9)]));
              reg271 = $signed($unsigned($signed($signed((reg195 < reg212)))));
            end
          else
            begin
              reg270 = $unsigned((~&(((reg175 ^ reg171) ?
                  (7'h40) : reg176) >= $unsigned(reg195[(1'h1):(1'h1)]))));
              reg272 <= wire247[(3'h7):(3'h7)];
            end
          if ($signed(reg257))
            begin
              reg273 <= $unsigned($signed($unsigned(reg195[(2'h2):(1'h0)])));
              reg274 <= reg182;
              reg275 <= reg149[(4'h8):(3'h6)];
              reg276 = (reg254[(4'hf):(2'h3)] & wire247);
              reg277 = forvar249;
            end
          else
            begin
              reg273 <= (8'hae);
            end
        end
      for (forvar278 = (1'h0); (forvar278 < (1'h0)); forvar278 = (forvar278 + (1'h1)))
        begin
          if (forvar258[(1'h0):(1'h0)])
            begin
              reg279 = ((~(reg159[(3'h4):(3'h4)] ?
                      ((~&reg202) ?
                          (&wire207) : (reg267 > reg256)) : wire246)) ?
                  $signed((((reg235 <= (8'hb5)) - wire207) >>> ((reg162 && forvar258) ?
                      $signed(reg136) : $signed((8'ha1))))) : reg136[(3'h6):(3'h4)]);
            end
          else
            begin
              reg279 = reg141[(2'h3):(2'h3)];
              reg280 = $signed($unsigned(wire245[(1'h0):(1'h0)]));
              reg281 = $signed((+(reg243 ?
                  $signed((+reg269)) : {reg231[(1'h0):(1'h0)],
                      reg235[(4'hc):(4'hc)]})));
            end
          reg282 <= (|reg140);
          reg283 <= {$unsigned({reg239[(3'h4):(3'h4)],
                  ((wire245 != wire248) ?
                      reg141 : (reg279 ? reg187 : (8'hbf)))})};
        end
      if ($signed((reg129[(5'h10):(1'h1)] <<< $unsigned({{(8'h9e), (8'ha5)}}))))
        begin
          if ($signed(reg141[(1'h0):(1'h0)]))
            begin
              reg284 = ($unsigned((!{(reg283 == wire127)})) <= forvar278[(5'h14):(4'hc)]);
              reg285 <= (&reg198);
              reg286 <= {(~^$signed(reg183[(3'h6):(3'h4)])),
                  $unsigned($signed(reg231))};
              reg287 <= $signed((~&reg133));
            end
          else
            begin
              reg284 = {$unsigned($unsigned(reg235)),
                  $unsigned((|{((8'ha7) != (8'hb8)), $signed(reg264)}))};
              reg288 = $signed(reg131);
              reg289 <= $signed(((wire120 ^ reg217[(4'ha):(1'h0)]) ?
                  reg168 : reg239));
              reg290 <= (~|(reg255[(4'he):(2'h2)] ?
                  (!((wire123 ?
                      (8'h9e) : wire247) | $unsigned(reg238))) : reg153[(4'ha):(1'h0)]));
              reg291 <= wire246[(4'ha):(4'h8)];
            end
          if ($signed($unsigned((~$unsigned((reg271 ? reg133 : reg254))))))
            begin
              reg292 <= $signed((reg134[(2'h3):(2'h2)] && (((reg239 != reg262) ?
                  reg264 : reg260) << $unsigned($signed(reg269)))));
            end
          else
            begin
              reg292 <= ($unsigned($signed(wire122)) || ($unsigned(reg158) ?
                  reg289 : (&$signed(reg176[(4'hc):(3'h5)]))));
              reg293 = {(((!reg240[(2'h3):(1'h1)]) - ($unsigned(reg239) != reg255[(1'h0):(1'h0)])) ?
                      {$signed((reg262 ? reg284 : reg157)),
                          reg244[(4'ha):(1'h1)]} : ((reg282[(2'h3):(2'h2)] <= {reg260}) ?
                          reg260 : $signed((~|forvar258)))),
                  (-$signed((forvar258[(3'h7):(3'h4)] ?
                      {reg148, reg284} : (reg155 + reg255))))};
              reg294 = $signed(reg129);
              reg295 <= reg231;
            end
          reg296 = {reg235[(4'hf):(3'h6)]};
          reg297 = wire123;
        end
      else
        begin
          reg284 = $unsigned(reg197[(4'hc):(4'hc)]);
          if ($signed($signed(((-(~&reg266)) ?
              reg271[(1'h0):(1'h0)] : $signed((+wire248))))))
            begin
              reg285 <= {$unsigned($unsigned((~^$unsigned(reg259))))};
              reg286 <= reg149;
              reg287 <= (8'hb2);
              reg288 = (((~&($unsigned(reg274) & $signed(wire121))) * $signed(wire126)) ?
                  $signed(((((8'ha1) ? wire124 : reg276) ?
                      (reg260 | reg255) : reg199) <<< $unsigned($signed(reg271)))) : ($signed((|(wire246 + forvar251))) ?
                      {$unsigned($unsigned(reg136)),
                          $unsigned($signed(reg136))} : reg250[(4'hc):(3'h4)]));
            end
          else
            begin
              reg288 = reg255[(1'h0):(1'h0)];
            end
          if ((!{({{wire205, reg252}} ?
                  reg275[(4'h8):(2'h3)] : $unsigned(reg176[(1'h1):(1'h1)]))}))
            begin
              reg289 <= reg131;
              reg293 = {reg264};
              reg294 = reg131[(5'h13):(3'h5)];
              reg295 <= reg268;
            end
          else
            begin
              reg289 <= reg250;
              reg290 <= (^(~$unsigned($signed({(7'h43)}))));
            end
          if ({(reg197 ?
                  (reg291 * ($unsigned(forvar251) - reg168)) : {$unsigned((~|reg285))}),
              $signed((($unsigned((8'hbc)) ? reg285 : reg256) ?
                  reg289 : (reg153[(5'h11):(4'h9)] ^~ wire124)))})
            begin
              reg298 <= (~^(wire120[(5'h12):(4'he)] - $signed($unsigned(reg209[(1'h0):(1'h0)]))));
              reg299 = ((((+{wire127, (8'ha3)}) ?
                  $signed($unsigned(reg239)) : ({reg231, reg133} ?
                      reg149 : (~reg198))) ~^ reg270) >>> reg201[(1'h1):(1'h0)]);
              reg300 = $signed($unsigned(wire120[(1'h1):(1'h0)]));
              reg301 = {$unsigned((!$signed(wire125[(4'hf):(4'ha)]))),
                  {{(reg269 | (reg140 << reg267))}}};
              reg302 = {$signed({({(8'hbb), reg300} < $unsigned(reg288))}),
                  reg284[(4'hf):(4'ha)]};
            end
          else
            begin
              reg296 = $signed((-reg235));
              reg297 = (8'ha8);
              reg298 <= $signed(forvar258[(3'h7):(3'h6)]);
            end
        end
      if ($unsigned($unsigned({$unsigned($signed(reg171))})))
        begin
          reg303 <= {{($unsigned((reg276 ? reg182 : reg186)) > $signed({reg140,
                      (8'hb0)}))}};
          if (($signed(reg217) >>> reg294))
            begin
              reg304 = $unsigned($unsigned(reg279[(2'h2):(1'h1)]));
            end
          else
            begin
              reg305 <= (reg158 ? $unsigned(reg137) : reg267);
              reg306 <= ((~(~(reg276[(3'h4):(1'h1)] ?
                  (wire247 ~^ wire120) : $unsigned(reg182)))) & reg271[(2'h2):(2'h2)]);
              reg307 <= {reg276[(3'h4):(1'h0)], reg292[(3'h7):(2'h3)]};
            end
          reg308 <= $unsigned(((((&reg307) & $unsigned(reg275)) < $unsigned(reg210)) ?
              (~|(~|(reg136 ? (7'h40) : wire122))) : reg160));
        end
      else
        begin
          reg303 <= ($unsigned(($signed((wire120 != reg159)) ?
              (8'hb1) : reg291)) != (wire124 ?
              (((wire122 ? reg220 : wire204) ?
                      $signed((8'hbe)) : $signed(reg259)) ?
                  reg305[(2'h3):(2'h2)] : reg238[(4'he):(4'he)]) : $signed(reg268)));
          if ({$unsigned((~|(!{reg240, reg256})))})
            begin
              reg305 <= reg263[(3'h7):(1'h1)];
              reg309 = (8'hb7);
              reg310 <= ((+$signed(($unsigned(reg303) < $signed(reg157)))) ?
                  $signed(reg265) : ($unsigned(reg259[(3'h7):(3'h5)]) ?
                      wire205 : (($signed(reg307) ?
                              $unsigned(reg282) : $unsigned((8'ha9))) ?
                          reg255 : ((~&reg153) ?
                              reg306[(2'h3):(1'h0)] : (reg137 << reg136)))));
              reg311 = forvar278;
              reg312 <= wire120[(1'h1):(1'h0)];
            end
          else
            begin
              reg305 <= (^~$signed($signed(({reg285} > (wire121 ?
                  reg301 : reg161)))));
              reg306 <= $signed($signed($signed($unsigned(reg310[(4'hc):(2'h2)]))));
            end
        end
    end
endmodule