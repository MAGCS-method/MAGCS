(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param1094 = (&((((7'h4c) ? (!(8'hb7)) : (^~(8'hbb))) ? ({(8'ha8), (7'h51), (8'hbb)} ? ((8'ha6) | (8'hb2)) : {(7'h45)}) : (&{(8'hba), (7'h47)})) << (^{(-(8'hb8)), {(8'hb7), (8'ha2)}, (+(8'hb1))}))), 
parameter param1095 = (({((param1094 ? param1094 : (8'ha3)) || (param1094 >> param1094))} ? (|param1094) : param1094) == {{{{param1094}}, {(+param1094), (|param1094), param1094}, (^~((8'ha6) ^~ param1094))}, (param1094 ^ (+(param1094 || param1094))), param1094}))
(y, clk, wire5, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h24b8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire5;
  input wire [(5'h17):(1'h0)] wire4;
  input wire signed [(5'h12):(1'h0)] wire3;
  input wire signed [(3'h5):(1'h0)] wire2;
  input wire [(5'h1c):(1'h0)] wire1;
  input wire signed [(2'h2):(1'h0)] wire0;
  wire signed [(5'h17):(1'h0)] wire1093;
  wire signed [(4'hd):(1'h0)] wire1092;
  wire [(2'h3):(1'h0)] wire1091;
  wire [(4'hf):(1'h0)] wire1090;
  wire signed [(5'h1a):(1'h0)] wire1089;
  wire [(4'h9):(1'h0)] wire1085;
  wire signed [(5'h1e):(1'h0)] wire881;
  wire signed [(5'h1e):(1'h0)] wire880;
  wire [(5'h18):(1'h0)] wire879;
  wire [(5'h1a):(1'h0)] wire855;
  wire signed [(4'h9):(1'h0)] wire854;
  wire [(3'h5):(1'h0)] wire853;
  wire [(5'h1e):(1'h0)] wire852;
  wire signed [(4'hb):(1'h0)] wire835;
  wire signed [(5'h13):(1'h0)] wire663;
  wire [(5'h1d):(1'h0)] wire620;
  wire [(4'h9):(1'h0)] wire76;
  wire [(5'h1b):(1'h0)] wire7;
  wire [(3'h6):(1'h0)] wire6;
  reg signed [(4'h8):(1'h0)] reg1088 = (1'h0);
  reg [(3'h7):(1'h0)] reg1087 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1086 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1082 = (1'h0);
  reg [(5'h18):(1'h0)] reg1081 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1080 = (1'h0);
  reg [(4'hf):(1'h0)] reg1078 = (1'h0);
  reg [(3'h7):(1'h0)] reg1076 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1075 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1074 = (1'h0);
  reg [(5'h11):(1'h0)] reg1072 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1061 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1068 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1067 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1057 = (1'h0);
  reg [(5'h11):(1'h0)] reg1054 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1053 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1051 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1049 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1045 = (1'h0);
  reg [(5'h19):(1'h0)] reg1041 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1039 = (1'h0);
  reg [(4'he):(1'h0)] reg1038 = (1'h0);
  reg [(4'ha):(1'h0)] reg1037 = (1'h0);
  reg [(4'hc):(1'h0)] reg1036 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1035 = (1'h0);
  reg [(2'h3):(1'h0)] reg1033 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1032 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1031 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1030 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1028 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1020 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1013 = (1'h0);
  reg [(3'h6):(1'h0)] reg1009 = (1'h0);
  reg [(5'h14):(1'h0)] reg1008 = (1'h0);
  reg [(2'h2):(1'h0)] reg1007 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg987 = (1'h0);
  reg [(4'hf):(1'h0)] reg1004 = (1'h0);
  reg [(2'h3):(1'h0)] reg1003 = (1'h0);
  reg [(4'hd):(1'h0)] reg1001 = (1'h0);
  reg [(5'h12):(1'h0)] reg1000 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg999 = (1'h0);
  reg [(4'hb):(1'h0)] reg998 = (1'h0);
  reg [(4'ha):(1'h0)] reg994 = (1'h0);
  reg [(5'h19):(1'h0)] reg993 = (1'h0);
  reg [(5'h1a):(1'h0)] reg992 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg989 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg988 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg986 = (1'h0);
  reg [(5'h1b):(1'h0)] reg982 = (1'h0);
  reg [(4'h9):(1'h0)] reg979 = (1'h0);
  reg [(5'h14):(1'h0)] reg978 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg977 = (1'h0);
  reg [(5'h13):(1'h0)] reg975 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg974 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg970 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg968 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg967 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg966 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg965 = (1'h0);
  reg [(5'h12):(1'h0)] reg964 = (1'h0);
  reg [(5'h18):(1'h0)] reg962 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg961 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg959 = (1'h0);
  reg [(5'h18):(1'h0)] reg956 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg955 = (1'h0);
  reg [(5'h11):(1'h0)] reg954 = (1'h0);
  reg [(5'h1a):(1'h0)] reg947 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg944 = (1'h0);
  reg [(5'h1a):(1'h0)] reg942 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg940 = (1'h0);
  reg [(5'h12):(1'h0)] reg939 = (1'h0);
  reg [(3'h7):(1'h0)] reg938 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg934 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg933 = (1'h0);
  reg [(5'h1d):(1'h0)] reg930 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg929 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg928 = (1'h0);
  reg [(2'h2):(1'h0)] reg926 = (1'h0);
  reg [(4'hc):(1'h0)] reg925 = (1'h0);
  reg [(5'h18):(1'h0)] reg922 = (1'h0);
  reg [(5'h10):(1'h0)] reg920 = (1'h0);
  reg [(5'h17):(1'h0)] reg917 = (1'h0);
  reg [(5'h16):(1'h0)] reg916 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg912 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg910 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg909 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg908 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg901 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg895 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg894 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg891 = (1'h0);
  reg [(4'hc):(1'h0)] reg888 = (1'h0);
  reg [(5'h15):(1'h0)] reg887 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg885 = (1'h0);
  reg [(3'h6):(1'h0)] reg883 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg872 = (1'h0);
  reg [(5'h19):(1'h0)] reg871 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg870 = (1'h0);
  reg [(5'h1c):(1'h0)] reg869 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg859 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg850 = (1'h0);
  reg [(4'hf):(1'h0)] reg848 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg847 = (1'h0);
  reg [(3'h6):(1'h0)] reg846 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg845 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg844 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg843 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg842 = (1'h0);
  reg [(4'he):(1'h0)] reg838 = (1'h0);
  reg [(4'hc):(1'h0)] reg833 = (1'h0);
  reg [(5'h13):(1'h0)] reg832 = (1'h0);
  reg [(5'h1d):(1'h0)] reg831 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg830 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg819 = (1'h0);
  reg [(4'h8):(1'h0)] reg817 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg816 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg815 = (1'h0);
  reg [(3'h5):(1'h0)] reg814 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg811 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg808 = (1'h0);
  reg [(5'h1b):(1'h0)] reg807 = (1'h0);
  reg [(5'h14):(1'h0)] reg804 = (1'h0);
  reg [(3'h7):(1'h0)] reg803 = (1'h0);
  reg signed [(4'he):(1'h0)] reg801 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg795 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg794 = (1'h0);
  reg [(5'h16):(1'h0)] reg793 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg786 = (1'h0);
  reg [(5'h11):(1'h0)] reg771 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg792 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg788 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg784 = (1'h0);
  reg [(4'h8):(1'h0)] reg783 = (1'h0);
  reg [(3'h5):(1'h0)] reg782 = (1'h0);
  reg [(5'h14):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg778 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg777 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg774 = (1'h0);
  reg [(5'h12):(1'h0)] reg766 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg764 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg763 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg762 = (1'h0);
  reg [(5'h15):(1'h0)] reg761 = (1'h0);
  reg [(4'ha):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg758 = (1'h0);
  reg [(5'h18):(1'h0)] reg756 = (1'h0);
  reg [(4'he):(1'h0)] reg754 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg753 = (1'h0);
  reg [(3'h6):(1'h0)] reg751 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg750 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg745 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg743 = (1'h0);
  reg [(5'h1a):(1'h0)] reg742 = (1'h0);
  reg [(4'hf):(1'h0)] reg738 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg737 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg736 = (1'h0);
  reg [(5'h12):(1'h0)] reg734 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg733 = (1'h0);
  reg [(4'ha):(1'h0)] reg728 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg727 = (1'h0);
  reg [(5'h1c):(1'h0)] reg726 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg719 = (1'h0);
  reg [(5'h1f):(1'h0)] reg717 = (1'h0);
  reg [(4'h9):(1'h0)] reg715 = (1'h0);
  reg [(5'h12):(1'h0)] reg714 = (1'h0);
  reg [(5'h11):(1'h0)] reg712 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg708 = (1'h0);
  reg [(3'h6):(1'h0)] reg704 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg701 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg700 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg697 = (1'h0);
  reg [(5'h19):(1'h0)] reg694 = (1'h0);
  reg [(4'ha):(1'h0)] reg691 = (1'h0);
  reg [(4'h8):(1'h0)] reg686 = (1'h0);
  reg [(4'h8):(1'h0)] reg685 = (1'h0);
  reg [(5'h11):(1'h0)] reg684 = (1'h0);
  reg [(5'h1d):(1'h0)] reg683 = (1'h0);
  reg [(4'hf):(1'h0)] reg682 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg681 = (1'h0);
  reg [(4'h9):(1'h0)] reg679 = (1'h0);
  reg [(5'h17):(1'h0)] reg678 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg677 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg675 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg674 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg672 = (1'h0);
  reg [(5'h11):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg668 = (1'h0);
  reg [(5'h17):(1'h0)] reg667 = (1'h0);
  reg [(5'h1a):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg664 = (1'h0);
  reg [(5'h1e):(1'h0)] reg662 = (1'h0);
  reg [(4'hf):(1'h0)] reg660 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg657 = (1'h0);
  reg [(5'h12):(1'h0)] reg655 = (1'h0);
  reg [(5'h13):(1'h0)] reg654 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg653 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg651 = (1'h0);
  reg [(5'h13):(1'h0)] reg648 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg647 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg642 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg640 = (1'h0);
  reg [(4'he):(1'h0)] reg639 = (1'h0);
  reg [(5'h10):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg637 = (1'h0);
  reg [(2'h3):(1'h0)] reg634 = (1'h0);
  reg [(5'h1b):(1'h0)] reg631 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg629 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg626 = (1'h0);
  reg [(4'h8):(1'h0)] reg625 = (1'h0);
  reg [(4'hc):(1'h0)] reg622 = (1'h0);
  reg [(3'h4):(1'h0)] reg11 = (1'h0);
  reg [(2'h3):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg14 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg16 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg10 = (1'h0);
  reg [(5'h18):(1'h0)] reg19 = (1'h0);
  reg [(5'h16):(1'h0)] reg21 = (1'h0);
  reg [(5'h19):(1'h0)] reg25 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg27 = (1'h0);
  reg [(4'hd):(1'h0)] reg32 = (1'h0);
  reg [(4'h8):(1'h0)] reg34 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg35 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg36 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg39 = (1'h0);
  reg [(5'h1a):(1'h0)] reg41 = (1'h0);
  reg [(5'h19):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg43 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg46 = (1'h0);
  reg [(4'hd):(1'h0)] reg47 = (1'h0);
  reg [(3'h7):(1'h0)] reg49 = (1'h0);
  reg [(5'h1e):(1'h0)] reg52 = (1'h0);
  reg [(2'h2):(1'h0)] reg58 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg63 = (1'h0);
  reg [(5'h1a):(1'h0)] reg64 = (1'h0);
  reg [(5'h19):(1'h0)] reg61 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg66 = (1'h0);
  reg [(5'h14):(1'h0)] reg68 = (1'h0);
  reg [(4'hd):(1'h0)] reg71 = (1'h0);
  reg [(5'h1c):(1'h0)] reg74 = (1'h0);
  reg [(5'h10):(1'h0)] reg75 = (1'h0);
  reg [(5'h13):(1'h0)] reg1083 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1079 = (1'h0);
  reg [(4'hc):(1'h0)] reg1077 = (1'h0);
  reg [(4'hf):(1'h0)] reg1073 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1071 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1070 = (1'h0);
  reg [(4'hf):(1'h0)] reg1069 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1056 = (1'h0);
  reg [(5'h14):(1'h0)] reg1055 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1066 = (1'h0);
  reg [(4'ha):(1'h0)] reg1065 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1064 = (1'h0);
  reg [(4'h8):(1'h0)] reg1063 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1062 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1061 = (1'h0);
  reg [(2'h2):(1'h0)] reg1060 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1059 = (1'h0);
  reg [(3'h4):(1'h0)] reg1058 = (1'h0);
  reg [(4'hb):(1'h0)] reg1056 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1055 = (1'h0);
  reg [(4'ha):(1'h0)] reg1052 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1048 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1047 = (1'h0);
  reg [(4'ha):(1'h0)] reg1046 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1044 = (1'h0);
  reg [(5'h17):(1'h0)] reg1043 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1042 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1040 = (1'h0);
  reg [(4'hd):(1'h0)] reg1034 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1029 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1027 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1026 = (1'h0);
  reg [(5'h16):(1'h0)] reg1025 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1024 = (1'h0);
  reg [(3'h5):(1'h0)] reg1023 = (1'h0);
  reg [(5'h13):(1'h0)] reg1022 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1021 = (1'h0);
  reg [(4'he):(1'h0)] reg1019 = (1'h0);
  reg [(4'ha):(1'h0)] reg1018 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1017 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1016 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1015 = (1'h0);
  reg [(5'h12):(1'h0)] reg1014 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1010 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1006 = (1'h0);
  reg [(5'h17):(1'h0)] forvar993 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg990 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar979 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1005 = (1'h0);
  reg [(3'h6):(1'h0)] reg1002 = (1'h0);
  reg [(5'h14):(1'h0)] reg997 = (1'h0);
  reg [(3'h5):(1'h0)] reg996 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg995 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg991 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar990 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar987 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg985 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg984 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg983 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg981 = (1'h0);
  reg [(5'h10):(1'h0)] reg980 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg976 = (1'h0);
  reg [(4'he):(1'h0)] reg973 = (1'h0);
  reg [(5'h19):(1'h0)] reg972 = (1'h0);
  reg [(4'he):(1'h0)] reg971 = (1'h0);
  reg [(5'h16):(1'h0)] reg969 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg963 = (1'h0);
  reg [(3'h6):(1'h0)] reg960 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg958 = (1'h0);
  reg [(5'h12):(1'h0)] reg957 = (1'h0);
  reg [(3'h6):(1'h0)] forvar953 = (1'h0);
  reg [(5'h19):(1'h0)] reg952 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg951 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg950 = (1'h0);
  reg [(5'h19):(1'h0)] reg949 = (1'h0);
  reg [(5'h17):(1'h0)] reg948 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg946 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg945 = (1'h0);
  reg [(4'ha):(1'h0)] reg943 = (1'h0);
  reg [(3'h7):(1'h0)] reg941 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg931 = (1'h0);
  reg [(5'h1d):(1'h0)] reg937 = (1'h0);
  reg [(3'h7):(1'h0)] reg936 = (1'h0);
  reg [(5'h14):(1'h0)] reg935 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg932 = (1'h0);
  reg [(4'h9):(1'h0)] forvar931 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg927 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg924 = (1'h0);
  reg [(4'ha):(1'h0)] reg923 = (1'h0);
  reg [(5'h19):(1'h0)] reg921 = (1'h0);
  reg [(5'h17):(1'h0)] reg919 = (1'h0);
  reg [(5'h19):(1'h0)] reg918 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg915 = (1'h0);
  reg [(3'h7):(1'h0)] reg914 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg913 = (1'h0);
  reg [(5'h1f):(1'h0)] reg911 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg907 = (1'h0);
  reg [(5'h19):(1'h0)] reg906 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar905 = (1'h0);
  reg [(3'h4):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg896 = (1'h0);
  reg [(5'h16):(1'h0)] reg902 = (1'h0);
  reg [(5'h16):(1'h0)] reg899 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg898 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg897 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar896 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg893 = (1'h0);
  reg [(4'hb):(1'h0)] reg892 = (1'h0);
  reg [(3'h5):(1'h0)] reg890 = (1'h0);
  reg [(5'h17):(1'h0)] reg889 = (1'h0);
  reg [(5'h1e):(1'h0)] reg886 = (1'h0);
  reg [(4'h9):(1'h0)] reg884 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg882 = (1'h0);
  reg [(5'h11):(1'h0)] reg878 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg877 = (1'h0);
  reg [(4'hf):(1'h0)] reg876 = (1'h0);
  reg [(4'hd):(1'h0)] forvar875 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg874 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar873 = (1'h0);
  reg [(3'h6):(1'h0)] reg867 = (1'h0);
  reg [(5'h13):(1'h0)] forvar866 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg865 = (1'h0);
  reg [(5'h18):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg863 = (1'h0);
  reg [(5'h11):(1'h0)] forvar862 = (1'h0);
  reg [(2'h2):(1'h0)] reg861 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg860 = (1'h0);
  reg [(5'h19):(1'h0)] reg858 = (1'h0);
  reg [(5'h16):(1'h0)] forvar857 = (1'h0);
  reg [(4'hf):(1'h0)] reg856 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg851 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg849 = (1'h0);
  reg [(5'h14):(1'h0)] forvar837 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg841 = (1'h0);
  reg [(5'h1d):(1'h0)] reg840 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg839 = (1'h0);
  reg [(3'h7):(1'h0)] reg837 = (1'h0);
  reg [(5'h1e):(1'h0)] reg836 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg834 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg829 = (1'h0);
  reg [(4'h9):(1'h0)] reg828 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg827 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar826 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg825 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg824 = (1'h0);
  reg [(5'h12):(1'h0)] reg823 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg822 = (1'h0);
  reg [(2'h2):(1'h0)] forvar821 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar820 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg818 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar813 = (1'h0);
  reg [(5'h15):(1'h0)] reg812 = (1'h0);
  reg [(3'h4):(1'h0)] reg810 = (1'h0);
  reg [(4'he):(1'h0)] reg809 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg806 = (1'h0);
  reg [(5'h1c):(1'h0)] reg805 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg802 = (1'h0);
  reg [(5'h15):(1'h0)] reg800 = (1'h0);
  reg [(3'h4):(1'h0)] reg799 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar798 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg797 = (1'h0);
  reg [(5'h1d):(1'h0)] reg796 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg791 = (1'h0);
  reg [(5'h1c):(1'h0)] reg790 = (1'h0);
  reg [(5'h19):(1'h0)] reg789 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg787 = (1'h0);
  reg [(4'hc):(1'h0)] forvar786 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg785 = (1'h0);
  reg [(5'h18):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg779 = (1'h0);
  reg [(4'ha):(1'h0)] reg776 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg775 = (1'h0);
  reg [(2'h2):(1'h0)] reg773 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg772 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar771 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg770 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg769 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg768 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg767 = (1'h0);
  reg signed [(4'he):(1'h0)] reg765 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar762 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg760 = (1'h0);
  reg [(5'h19):(1'h0)] reg757 = (1'h0);
  reg signed [(4'he):(1'h0)] reg755 = (1'h0);
  reg [(5'h1a):(1'h0)] reg752 = (1'h0);
  reg [(5'h1e):(1'h0)] reg749 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar748 = (1'h0);
  reg [(4'hc):(1'h0)] reg747 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg746 = (1'h0);
  reg [(4'hc):(1'h0)] reg744 = (1'h0);
  reg [(5'h19):(1'h0)] reg741 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar740 = (1'h0);
  reg [(4'hb):(1'h0)] reg739 = (1'h0);
  reg [(5'h1f):(1'h0)] reg735 = (1'h0);
  reg [(3'h6):(1'h0)] reg732 = (1'h0);
  reg [(5'h1e):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg730 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg729 = (1'h0);
  reg [(3'h5):(1'h0)] reg725 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg724 = (1'h0);
  reg [(4'hd):(1'h0)] reg723 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg722 = (1'h0);
  reg [(4'hd):(1'h0)] reg721 = (1'h0);
  reg [(3'h5):(1'h0)] forvar720 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg718 = (1'h0);
  reg [(5'h1f):(1'h0)] reg716 = (1'h0);
  reg [(5'h13):(1'h0)] forvar713 = (1'h0);
  reg [(5'h13):(1'h0)] reg711 = (1'h0);
  reg [(5'h1d):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar709 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg707 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg706 = (1'h0);
  reg [(5'h10):(1'h0)] reg705 = (1'h0);
  reg [(4'hb):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg702 = (1'h0);
  reg [(5'h15):(1'h0)] reg699 = (1'h0);
  reg [(5'h17):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg696 = (1'h0);
  reg [(3'h7):(1'h0)] reg695 = (1'h0);
  reg [(2'h3):(1'h0)] reg693 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar692 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg690 = (1'h0);
  reg [(4'h8):(1'h0)] reg689 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg688 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg687 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg680 = (1'h0);
  reg [(4'hd):(1'h0)] forvar676 = (1'h0);
  reg [(4'h9):(1'h0)] reg673 = (1'h0);
  reg [(5'h1b):(1'h0)] reg671 = (1'h0);
  reg [(4'h9):(1'h0)] reg669 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg666 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg661 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg658 = (1'h0);
  reg [(3'h6):(1'h0)] reg656 = (1'h0);
  reg [(4'ha):(1'h0)] forvar652 = (1'h0);
  reg signed [(4'he):(1'h0)] reg650 = (1'h0);
  reg [(5'h18):(1'h0)] forvar649 = (1'h0);
  reg [(5'h1a):(1'h0)] reg627 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg646 = (1'h0);
  reg [(2'h2):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg644 = (1'h0);
  reg [(5'h17):(1'h0)] reg643 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar642 = (1'h0);
  reg [(4'hc):(1'h0)] reg641 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg636 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg635 = (1'h0);
  reg [(5'h13):(1'h0)] reg633 = (1'h0);
  reg [(5'h12):(1'h0)] reg632 = (1'h0);
  reg [(5'h10):(1'h0)] reg630 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg628 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar627 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg73 = (1'h0);
  reg [(5'h19):(1'h0)] reg72 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar67 = (1'h0);
  reg [(5'h13):(1'h0)] reg65 = (1'h0);
  reg signed [(4'he):(1'h0)] reg62 = (1'h0);
  reg [(5'h12):(1'h0)] forvar61 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg60 = (1'h0);
  reg [(4'h9):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg57 = (1'h0);
  reg [(5'h18):(1'h0)] forvar56 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg55 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg54 = (1'h0);
  reg [(4'ha):(1'h0)] forvar53 = (1'h0);
  reg [(5'h1b):(1'h0)] reg51 = (1'h0);
  reg [(4'he):(1'h0)] reg50 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg48 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg45 = (1'h0);
  reg [(2'h2):(1'h0)] reg44 = (1'h0);
  reg [(5'h16):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar38 = (1'h0);
  reg [(5'h16):(1'h0)] reg37 = (1'h0);
  reg [(5'h1b):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg31 = (1'h0);
  reg [(5'h1e):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg29 = (1'h0);
  reg [(5'h13):(1'h0)] reg28 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg23 = (1'h0);
  reg [(5'h1f):(1'h0)] reg22 = (1'h0);
  reg [(5'h1c):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar19 = (1'h0);
  reg [(4'he):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg17 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg15 = (1'h0);
  reg [(4'he):(1'h0)] reg12 = (1'h0);
  reg [(5'h11):(1'h0)] forvar10 = (1'h0);
  reg [(2'h2):(1'h0)] reg9 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg8 = (1'h0);
  assign y = {wire1093,
                 wire1092,
                 wire1091,
                 wire1090,
                 wire1089,
                 wire1085,
                 wire881,
                 wire880,
                 wire879,
                 wire855,
                 wire854,
                 wire853,
                 wire852,
                 wire835,
                 wire663,
                 wire620,
                 wire76,
                 wire7,
                 wire6,
                 reg1088,
                 reg1087,
                 reg1086,
                 reg1084,
                 reg1082,
                 reg1081,
                 reg1080,
                 reg1078,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1072,
                 reg1061,
                 reg1068,
                 reg1067,
                 reg1057,
                 reg1054,
                 reg1053,
                 reg1051,
                 reg1050,
                 reg1049,
                 reg1045,
                 reg1041,
                 reg1039,
                 reg1038,
                 reg1037,
                 reg1036,
                 reg1035,
                 reg1033,
                 reg1032,
                 reg1031,
                 reg1030,
                 reg1028,
                 reg1020,
                 reg1013,
                 reg1009,
                 reg1008,
                 reg1007,
                 reg987,
                 reg1004,
                 reg1003,
                 reg1001,
                 reg1000,
                 reg999,
                 reg998,
                 reg994,
                 reg993,
                 reg992,
                 reg989,
                 reg988,
                 reg986,
                 reg982,
                 reg979,
                 reg978,
                 reg977,
                 reg975,
                 reg974,
                 reg970,
                 reg968,
                 reg967,
                 reg966,
                 reg965,
                 reg964,
                 reg962,
                 reg961,
                 reg959,
                 reg956,
                 reg955,
                 reg954,
                 reg947,
                 reg944,
                 reg942,
                 reg940,
                 reg939,
                 reg938,
                 reg934,
                 reg933,
                 reg930,
                 reg929,
                 reg928,
                 reg926,
                 reg925,
                 reg922,
                 reg920,
                 reg917,
                 reg916,
                 reg912,
                 reg910,
                 reg909,
                 reg908,
                 reg901,
                 reg900,
                 reg895,
                 reg894,
                 reg891,
                 reg888,
                 reg887,
                 reg885,
                 reg883,
                 reg872,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 reg859,
                 reg850,
                 reg848,
                 reg847,
                 reg846,
                 reg845,
                 reg844,
                 reg843,
                 reg842,
                 reg838,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 reg819,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg811,
                 reg808,
                 reg807,
                 reg804,
                 reg803,
                 reg801,
                 reg795,
                 reg794,
                 reg793,
                 reg786,
                 reg771,
                 reg792,
                 reg788,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 reg778,
                 reg777,
                 reg774,
                 reg766,
                 reg764,
                 reg763,
                 reg762,
                 reg761,
                 reg759,
                 reg758,
                 reg756,
                 reg754,
                 reg753,
                 reg751,
                 reg750,
                 reg745,
                 reg743,
                 reg742,
                 reg738,
                 reg737,
                 reg736,
                 reg734,
                 reg733,
                 reg728,
                 reg727,
                 reg726,
                 reg719,
                 reg717,
                 reg715,
                 reg714,
                 reg712,
                 reg708,
                 reg704,
                 reg701,
                 reg700,
                 reg697,
                 reg694,
                 reg691,
                 reg686,
                 reg685,
                 reg684,
                 reg683,
                 reg682,
                 reg681,
                 reg679,
                 reg678,
                 reg677,
                 reg675,
                 reg674,
                 reg672,
                 reg670,
                 reg668,
                 reg667,
                 reg665,
                 reg664,
                 reg662,
                 reg660,
                 reg659,
                 reg657,
                 reg655,
                 reg654,
                 reg653,
                 reg651,
                 reg648,
                 reg647,
                 reg642,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg634,
                 reg631,
                 reg629,
                 reg626,
                 reg625,
                 reg622,
                 reg11,
                 reg13,
                 reg14,
                 reg16,
                 reg10,
                 reg19,
                 reg21,
                 reg25,
                 reg27,
                 reg32,
                 reg34,
                 reg35,
                 reg36,
                 reg39,
                 reg41,
                 reg42,
                 reg43,
                 reg46,
                 reg47,
                 reg49,
                 reg52,
                 reg58,
                 reg63,
                 reg64,
                 reg61,
                 reg66,
                 reg68,
                 reg71,
                 reg74,
                 reg75,
                 reg1083,
                 reg1079,
                 reg1077,
                 reg1073,
                 forvar1071,
                 forvar1070,
                 reg1069,
                 forvar1056,
                 reg1055,
                 reg1066,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 forvar1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 reg1056,
                 forvar1055,
                 reg1052,
                 reg1048,
                 reg1047,
                 reg1046,
                 reg1044,
                 reg1043,
                 reg1042,
                 reg1040,
                 reg1034,
                 reg1029,
                 reg1027,
                 reg1026,
                 reg1025,
                 reg1024,
                 reg1023,
                 reg1022,
                 reg1021,
                 reg1019,
                 reg1018,
                 forvar1017,
                 reg1016,
                 reg1015,
                 reg1014,
                 reg1012,
                 reg1011,
                 reg1010,
                 forvar1006,
                 forvar993,
                 reg990,
                 forvar979,
                 reg1005,
                 reg1002,
                 reg997,
                 reg996,
                 reg995,
                 reg991,
                 forvar990,
                 forvar987,
                 reg985,
                 reg984,
                 reg983,
                 reg981,
                 reg980,
                 reg976,
                 reg973,
                 reg972,
                 reg971,
                 reg969,
                 reg963,
                 reg960,
                 reg958,
                 reg957,
                 forvar953,
                 reg952,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 reg946,
                 reg945,
                 reg943,
                 reg941,
                 reg931,
                 reg937,
                 reg936,
                 reg935,
                 reg932,
                 forvar931,
                 reg927,
                 reg924,
                 reg923,
                 reg921,
                 reg919,
                 reg918,
                 reg915,
                 reg914,
                 reg913,
                 reg911,
                 reg907,
                 reg906,
                 forvar905,
                 reg904,
                 reg903,
                 reg896,
                 reg902,
                 reg899,
                 reg898,
                 reg897,
                 forvar896,
                 reg893,
                 reg892,
                 reg890,
                 reg889,
                 reg886,
                 reg884,
                 reg882,
                 reg878,
                 reg877,
                 reg876,
                 forvar875,
                 reg874,
                 forvar873,
                 reg867,
                 forvar866,
                 reg865,
                 reg864,
                 reg863,
                 forvar862,
                 reg861,
                 reg860,
                 reg858,
                 forvar857,
                 reg856,
                 reg851,
                 reg849,
                 forvar837,
                 reg841,
                 reg840,
                 reg839,
                 reg837,
                 reg836,
                 reg834,
                 reg829,
                 reg828,
                 reg827,
                 forvar826,
                 reg825,
                 reg824,
                 reg823,
                 reg822,
                 forvar821,
                 forvar820,
                 reg818,
                 forvar813,
                 reg812,
                 reg810,
                 reg809,
                 reg806,
                 reg805,
                 reg802,
                 reg800,
                 reg799,
                 forvar798,
                 reg797,
                 reg796,
                 reg791,
                 reg790,
                 reg789,
                 reg787,
                 forvar786,
                 reg785,
                 reg780,
                 reg779,
                 reg776,
                 reg775,
                 reg773,
                 reg772,
                 forvar771,
                 reg770,
                 reg769,
                 reg768,
                 reg767,
                 reg765,
                 forvar762,
                 reg760,
                 reg757,
                 reg755,
                 reg752,
                 reg749,
                 forvar748,
                 reg747,
                 reg746,
                 reg744,
                 reg741,
                 forvar740,
                 reg739,
                 reg735,
                 reg732,
                 reg731,
                 reg730,
                 reg729,
                 reg725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 forvar720,
                 reg718,
                 reg716,
                 forvar713,
                 reg711,
                 reg710,
                 forvar709,
                 reg707,
                 reg706,
                 reg705,
                 reg703,
                 reg702,
                 reg699,
                 reg698,
                 reg696,
                 reg695,
                 reg693,
                 forvar692,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 reg680,
                 forvar676,
                 reg673,
                 reg671,
                 reg669,
                 reg666,
                 reg661,
                 reg658,
                 reg656,
                 forvar652,
                 reg650,
                 forvar649,
                 reg627,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 forvar642,
                 reg641,
                 reg636,
                 reg635,
                 reg633,
                 reg632,
                 reg630,
                 reg628,
                 forvar627,
                 reg624,
                 reg623,
                 reg73,
                 reg72,
                 reg70,
                 reg69,
                 forvar67,
                 reg65,
                 reg62,
                 forvar61,
                 reg60,
                 reg59,
                 reg57,
                 forvar56,
                 reg55,
                 reg54,
                 forvar53,
                 reg51,
                 reg50,
                 reg48,
                 reg45,
                 reg44,
                 reg40,
                 forvar38,
                 reg37,
                 reg33,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg26,
                 reg24,
                 reg23,
                 reg22,
                 reg20,
                 forvar19,
                 reg18,
                 reg17,
                 reg15,
                 reg12,
                 forvar10,
                 reg9,
                 reg8,
                 (1'h0)};
  assign wire6 = wire3[(5'h11):(2'h3)];
  assign wire7 = $unsigned({$unsigned($unsigned((&wire1)))});
  always
    @(posedge clk) begin
      if ($signed((wire4[(3'h5):(3'h5)] >> {wire1})))
        begin
          reg8 = $unsigned($unsigned(wire0[(1'h1):(1'h0)]));
          reg9 = $signed((wire0[(1'h1):(1'h0)] + ((&{(8'hbc),
              wire4,
              (8'haa)}) >> $signed($signed(wire5)))));
          for (forvar10 = (1'h0); (forvar10 < (1'h0)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg11 <= $signed((~wire4[(4'hb):(3'h7)]));
              reg12 = wire2;
            end
          if (wire7[(3'h6):(3'h4)])
            begin
              reg13 <= ($unsigned({wire0[(1'h0):(1'h0)]}) ?
                  (((~(wire3 >>> wire7)) ~^ (wire0 << (7'h51))) ?
                      (+($signed(reg11) ?
                          {wire0} : (~^(8'hb8)))) : ($signed({wire1,
                              wire4,
                              wire1}) ?
                          ((|wire3) == $unsigned(wire6)) : ((wire5 - reg9) ?
                              (wire4 ? wire1 : wire4) : (wire5 ?
                                  wire0 : (8'had))))) : (~&($signed((~|reg9)) - wire0[(1'h1):(1'h0)])));
              reg14 <= ($signed(((~&reg9) ^ $signed((^~wire7)))) ?
                  ((~wire5) ?
                      $unsigned(forvar10[(1'h1):(1'h1)]) : $signed($unsigned((&wire3)))) : $signed(($unsigned(reg12[(3'h7):(3'h5)]) == ($signed(reg11) ?
                      (reg13 && wire2) : wire4))));
              reg15 = reg9[(2'h2):(2'h2)];
              reg16 <= (wire1[(4'ha):(1'h1)] ?
                  $signed((8'ha2)) : $signed(({{wire0, (7'h43), reg9}, reg13} ?
                      {reg8[(2'h3):(2'h3)]} : (7'h45))));
              reg17 = ((~^forvar10) ?
                  $unsigned((wire3[(2'h3):(2'h2)] ?
                      $unsigned((reg12 ?
                          (8'h9c) : forvar10)) : reg15[(4'ha):(4'h9)])) : $signed((($signed(wire1) >> ((7'h57) ?
                          wire6 : reg14)) ?
                      (~^reg11[(3'h4):(1'h1)]) : wire7)));
            end
          else
            begin
              reg15 = reg14[(4'hb):(3'h7)];
              reg17 = reg8;
              reg18 = $signed((~^$signed((8'hac))));
            end
          for (forvar19 = (1'h0); (forvar19 < (2'h2)); forvar19 = (forvar19 + (1'h1)))
            begin
              reg20 = forvar10;
            end
        end
      else
        begin
          if ((wire0[(2'h2):(2'h2)] ?
              wire1 : ($signed($signed(reg20)) ?
                  $unsigned(((7'h50) > wire5[(1'h0):(1'h0)])) : $unsigned(wire7[(4'h9):(4'h8)]))))
            begin
              reg8 = wire3;
            end
          else
            begin
              reg10 <= reg18[(3'h4):(2'h2)];
              reg12 = forvar10[(4'hc):(4'ha)];
              reg13 <= wire0;
              reg15 = ((~$unsigned(reg9)) ?
                  ((reg14 > wire4) != (($signed(reg15) ?
                          (forvar10 ~^ wire4) : reg20[(5'h19):(2'h3)]) ?
                      $unsigned({wire0,
                          reg10,
                          wire5}) : reg16[(1'h1):(1'h0)])) : wire1[(5'h1c):(4'hb)]);
              reg17 = reg17;
            end
          if (wire7)
            begin
              reg19 <= $unsigned((wire0 && $unsigned(($signed(reg15) ?
                  $unsigned(wire7) : (reg10 ? forvar19 : (8'ha9))))));
              reg21 <= reg12;
              reg22 = $signed(reg12[(4'hb):(4'hb)]);
              reg23 = ((~($unsigned(forvar10[(4'hd):(1'h0)]) ?
                      (^~(reg19 ?
                          reg15 : (8'hb5))) : $unsigned((reg14 > wire7)))) ?
                  wire2[(3'h4):(2'h2)] : wire2);
              reg24 = {{{$signed(reg11[(1'h0):(1'h0)])},
                      (reg23 ? reg19 : $unsigned((^reg10))),
                      reg11},
                  $unsigned((reg14[(4'hb):(3'h4)] ^~ ($signed(reg10) ?
                      $signed(reg13) : $unsigned(wire2)))),
                  {(reg8 ?
                          $unsigned(wire1) : ((forvar19 >= wire0) ?
                              reg8[(1'h1):(1'h1)] : (reg16 >= wire0)))}};
              reg25 <= reg9[(1'h0):(1'h0)];
              reg26 = reg24;
            end
          else
            begin
              reg18 = (reg9 ?
                  $signed({((reg8 == reg9) < (reg19 >= reg8)),
                      (|wire4[(3'h5):(3'h4)]),
                      ((reg13 <= reg14) ?
                          (wire1 ?
                              wire2 : reg15) : forvar19)}) : $unsigned(reg20[(3'h6):(3'h6)]));
              reg20 = reg11[(1'h0):(1'h0)];
            end
          reg27 <= (!$unsigned(reg10[(1'h1):(1'h1)]));
          reg28 = wire1[(2'h3):(1'h0)];
          reg29 = $signed($unsigned((7'h50)));
          reg30 = (($unsigned(((reg15 ?
                  reg13 : forvar10) - reg10[(1'h1):(1'h1)])) >> ((~&$signed(reg19)) < ($unsigned(reg29) == {wire3,
                  reg19}))) ?
              {forvar10, $signed({reg28[(1'h1):(1'h1)]})} : ((~^((reg17 ?
                      reg14 : reg26) ?
                  {reg16,
                      (8'hb5),
                      reg15} : (reg25 <<< (8'ha6)))) && $unsigned((-reg9))));
          if (($unsigned((~^$signed((|reg23)))) ?
              (((&$unsigned(wire0)) + $signed(reg12)) >> (~&$signed((8'ha3)))) : wire3[(4'hd):(3'h6)]))
            begin
              reg31 = reg24[(2'h2):(1'h1)];
              reg32 <= (&{($signed((reg30 ? reg15 : (8'hba))) ?
                      ({wire0, (7'h54)} ? (reg19 | reg28) : reg30) : wire1)});
              reg33 = ($unsigned((~&reg30)) * wire0[(1'h0):(1'h0)]);
              reg34 <= $unsigned((reg24 < ($unsigned(reg25[(3'h6):(3'h4)]) ^ wire4)));
              reg35 <= $unsigned(reg33[(4'ha):(1'h0)]);
            end
          else
            begin
              reg32 <= ($signed(($unsigned(reg26[(2'h3):(1'h1)]) ?
                  (7'h55) : $signed((reg25 || reg15)))) >> $signed($unsigned($signed(wire4))));
              reg34 <= (~^$unsigned(((reg27[(3'h7):(3'h7)] ?
                      forvar10 : reg33[(5'h15):(4'hd)]) ?
                  ($unsigned(reg15) ?
                      (-reg15) : $unsigned(reg11)) : {(-forvar10),
                      wire2[(1'h0):(1'h0)]})));
              reg35 <= wire1[(2'h3):(2'h3)];
              reg36 <= (8'h9e);
              reg37 = (~wire4[(4'hd):(4'h8)]);
            end
        end
      for (forvar38 = (1'h0); (forvar38 < (2'h3)); forvar38 = (forvar38 + (1'h1)))
        begin
          if (wire3)
            begin
              reg39 <= reg34;
              reg40 = ($signed((((reg39 ^~ forvar10) | (reg8 ?
                      wire0 : wire4)) ~^ ($unsigned((8'ha3)) ?
                      $unsigned(reg39) : (^~reg28)))) ?
                  $unsigned(reg28) : (($unsigned(reg32[(4'h9):(2'h2)]) ?
                          ((7'h4a) ?
                              $unsigned(reg35) : reg39[(4'h9):(4'h8)]) : (8'hbc)) ?
                      reg30[(4'hb):(3'h4)] : (8'hac)));
              reg41 <= $unsigned(($unsigned((^~(reg25 - (7'h54)))) ?
                  wire6 : (~wire1[(5'h10):(3'h5)])));
            end
          else
            begin
              reg40 = ((((-$unsigned(reg31)) ?
                      $unsigned($signed(reg15)) : ((reg17 ?
                          reg26 : reg19) <<< (reg34 < (7'h4d)))) ?
                  (~|reg35[(5'h11):(1'h0)]) : (~&reg24)) < (($signed(reg37) + ((~|(8'ha3)) ~^ $signed(reg14))) || {(reg40 & wire1[(4'h8):(3'h7)]),
                  (&(!reg35))}));
            end
          reg42 <= reg9[(1'h1):(1'h1)];
          if (wire3[(4'h8):(2'h3)])
            begin
              reg43 <= (7'h4e);
              reg44 = (!((|(8'h9e)) ?
                  forvar38 : ($signed(reg40[(4'hb):(3'h6)]) ~^ {(reg36 ^~ reg30)})));
            end
          else
            begin
              reg44 = {$signed(reg18[(4'hd):(4'hb)]),
                  $signed(($unsigned((!forvar19)) ?
                      $unsigned($unsigned(forvar38)) : ((8'haa) ?
                          {reg34, (8'hb0), reg44} : (reg15 >> reg11)))),
                  reg37[(4'he):(4'hd)]};
              reg45 = $unsigned(((~|$unsigned((-wire3))) ?
                  $signed(reg24[(4'he):(4'hb)]) : $signed(($unsigned(reg36) <= (reg19 ?
                      (8'hbc) : reg42)))));
              reg46 <= (reg45 * (-$unsigned(($unsigned(reg11) ~^ reg39[(4'ha):(2'h3)]))));
              reg47 <= (|($unsigned(forvar10[(4'he):(3'h5)]) ?
                  reg29[(4'hd):(4'ha)] : (&($unsigned(forvar10) < (+reg21)))));
              reg48 = $signed((reg22 > reg36));
              reg49 <= (~&($unsigned(forvar38) & $signed({(reg39 && reg11)})));
              reg50 = reg34;
            end
          reg51 = (!(reg49 >= reg27[(4'h8):(1'h1)]));
          reg52 <= {(8'hab),
              (7'h4c),
              {$signed(reg51[(4'ha):(2'h2)]), reg8[(2'h2):(2'h2)]}};
          for (forvar53 = (1'h0); (forvar53 < (1'h1)); forvar53 = (forvar53 + (1'h1)))
            begin
              reg54 = (((!(reg50 ? reg28 : $signed(reg33))) << (~|reg9)) ?
                  reg23 : reg29);
            end
        end
      reg55 = reg11[(2'h2):(2'h2)];
      for (forvar56 = (1'h0); (forvar56 < (2'h3)); forvar56 = (forvar56 + (1'h1)))
        begin
          reg57 = reg15;
          reg58 <= wire1;
        end
      if (reg10[(1'h0):(1'h0)])
        begin
          reg59 = (|wire5);
          reg60 = ({(|$unsigned($signed(reg45))),
                  $signed((reg28 * $signed(reg39)))} ?
              ($unsigned($signed((reg51 >= reg55))) ?
                  reg41 : reg30[(4'hf):(4'ha)]) : wire7[(5'h16):(4'h8)]);
          for (forvar61 = (1'h0); (forvar61 < (3'h6)); forvar61 = (forvar61 + (1'h1)))
            begin
              reg62 = reg40;
              reg63 <= $unsigned((reg42 ?
                  $unsigned({(~&(8'ha8))}) : (reg9 != ((8'h9f) - (-reg33)))));
              reg64 <= reg35;
            end
          reg65 = ((($signed({reg19}) ?
              (reg14 * $unsigned(reg54)) : ((reg25 ?
                  reg15 : (7'h57)) ~^ reg24)) || (reg63 << (reg51[(1'h1):(1'h0)] ?
              (reg25 ?
                  (7'h44) : reg31) : (~|reg62)))) ~^ ((reg13[(1'h1):(1'h0)] ?
                  ({reg58, (7'h52), reg51} == $signed(reg51)) : {(&wire4),
                      $unsigned(reg41),
                      (reg43 ? (8'hac) : (7'h42))}) ?
              ((reg28 > reg27) != ($unsigned(reg40) ^ reg32)) : (reg57[(1'h1):(1'h0)] >= (reg31 ?
                  reg26 : $unsigned(reg33)))));
        end
      else
        begin
          if (wire1)
            begin
              reg59 = $unsigned(reg32);
              reg61 <= ($signed((((reg46 >>> reg26) ?
                      reg16[(1'h1):(1'h1)] : reg63) == (forvar38[(5'h12):(5'h10)] ?
                      ((8'ha2) >> (8'ha2)) : (reg13 ? reg59 : reg46)))) ?
                  {(^~$unsigned($signed(reg20)))} : reg26);
              reg62 = {$signed(forvar61[(5'h10):(3'h5)]),
                  ((((reg46 & wire2) * (reg8 || reg21)) ?
                      wire2 : ($signed(reg29) > reg65)) - $unsigned(reg43))};
              reg63 <= {$unsigned(reg61[(4'ha):(4'h8)])};
            end
          else
            begin
              reg59 = $unsigned(((+(&(reg26 ^~ forvar61))) & (!((reg52 | reg40) ?
                  $unsigned(reg45) : $unsigned(reg49)))));
              reg60 = reg52;
            end
          reg65 = $signed(((wire1[(5'h16):(5'h13)] ?
                  {$signed(reg37), $unsigned((7'h57))} : ((forvar53 ?
                      reg44 : reg20) <= reg39)) ?
              reg58[(1'h0):(1'h0)] : {(+$unsigned(forvar56)),
                  reg33,
                  {reg21[(4'he):(2'h2)],
                      ((8'hb6) ? reg26 : (8'ha0)),
                      $unsigned(forvar19)}}));
          reg66 <= $unsigned((^reg23[(4'he):(2'h3)]));
          for (forvar67 = (1'h0); (forvar67 < (2'h3)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 <= reg43;
              reg69 = wire3;
              reg70 = reg34[(2'h2):(1'h1)];
              reg71 <= $unsigned($signed((&$signed((wire4 >= forvar67)))));
              reg72 = {$unsigned(reg71[(4'hb):(3'h6)]),
                  {forvar61, $signed(reg62)},
                  $unsigned($unsigned(((forvar61 ^ reg20) ?
                      {reg51, reg54} : wire3)))};
              reg73 = ($unsigned($unsigned(({reg31} ?
                      (8'ha1) : {reg62, reg72}))) ?
                  $unsigned((&(^~$signed(reg28)))) : (|(((reg43 > (8'hb3)) || (~reg15)) > {(^reg52)})));
              reg74 <= {(-(-(^~(7'h55))))};
            end
        end
      reg75 <= $signed(reg61[(5'h15):(4'hd)]);
    end
  assign wire76 = reg32;
  module77 #() modinst621 (.wire80(reg74), .clk(clk), .y(wire620), .wire81(reg68), .wire79(reg32), .wire78(reg61), .wire82(reg25));
  always
    @(posedge clk) begin
      if (reg32)
        begin
          if ((($signed($signed((wire76 ?
              reg32 : wire6))) >= reg64) + {(wire4 >>> ((reg13 ?
                      reg13 : reg52) ?
                  (^reg49) : (7'h53))),
              {(reg64 * (reg47 ~^ wire0))},
              (wire5[(3'h4):(3'h4)] || (~&(reg74 & (7'h4d))))}))
            begin
              reg622 <= $unsigned((({(reg34 ? wire76 : reg71), $signed(reg13)} ?
                      (|(~&(8'ha6))) : (~|(~&reg10))) ?
                  {$unsigned((reg32 ? (7'h49) : wire0)),
                      reg42[(4'ha):(4'h9)],
                      reg10[(1'h1):(1'h0)]} : {reg42,
                      $unsigned(wire3),
                      reg11}));
              reg623 = {$signed($unsigned(wire3[(5'h10):(2'h3)])),
                  reg43[(4'hb):(4'h8)],
                  {(~&reg64),
                      (((7'h52) != (reg13 << reg49)) ?
                          (((7'h51) ?
                              wire0 : (8'hbe)) != $signed(reg39)) : (8'h9e)),
                      (wire0[(1'h0):(1'h0)] & (+((8'hb7) ? reg10 : reg75)))}};
              reg624 = $unsigned($unsigned($signed((reg66 << wire2[(2'h3):(2'h3)]))));
              reg625 <= $signed($unsigned($unsigned(wire5[(2'h3):(2'h3)])));
            end
          else
            begin
              reg622 <= ({{($unsigned(wire0) || (reg11 > (8'ha0))),
                      ($signed(reg39) ? $unsigned(wire620) : (reg46 | reg14)),
                      ((reg47 ? reg52 : reg623) ?
                          (~^(8'ha4)) : reg68[(1'h0):(1'h0)])},
                  ({$signed(reg19), (reg58 >>> reg39)} ?
                      $unsigned($signed(reg47)) : {(reg68 ?
                              (8'hbf) : reg43)})} || wire1[(5'h17):(5'h13)]);
              reg623 = (((7'h4d) ?
                  $signed(reg622) : {$unsigned(reg36[(1'h1):(1'h0)]),
                      ((^reg624) ?
                          $signed(reg47) : reg61)}) <= $signed($unsigned({$signed(reg64),
                  reg21[(5'h14):(5'h10)]})));
              reg625 <= reg623[(5'h11):(4'hd)];
            end
          reg626 <= $unsigned(reg11[(2'h2):(1'h1)]);
          for (forvar627 = (1'h0); (forvar627 < (3'h5)); forvar627 = (forvar627 + (1'h1)))
            begin
              reg628 = reg66;
              reg629 <= (|$unsigned(((|$signed((8'hb9))) + reg19)));
              reg630 = $unsigned(({reg58,
                  ($unsigned(wire7) - (^~(8'hbd))),
                  (&(reg625 - reg16))} <<< reg36[(1'h0):(1'h0)]));
              reg631 <= $signed((|reg624));
            end
          if (($signed({(reg46[(2'h2):(2'h2)] == (reg622 ? wire3 : reg32)),
              $unsigned(((7'h52) ?
                  wire2 : reg35))}) <= $signed($unsigned(($unsigned(reg66) && $unsigned((8'hb2)))))))
            begin
              reg632 = $signed($signed(((|reg622[(3'h6):(3'h4)]) ?
                  ((8'hba) ?
                      (~&reg49) : (~&forvar627)) : (|wire4[(1'h0):(1'h0)]))));
              reg633 = $signed(((($signed(reg14) >>> {reg58,
                      reg61}) ~^ (~&(reg74 <= wire620))) ?
                  reg628 : (($unsigned(reg629) == $unsigned(reg27)) <<< reg11[(1'h0):(1'h0)])));
              reg634 <= (7'h43);
              reg635 = $unsigned(reg622[(3'h5):(1'h1)]);
              reg636 = $signed($unsigned($signed($unsigned({reg27, reg13}))));
              reg637 <= ($unsigned((reg631[(5'h15):(3'h4)] ?
                      (^~(&reg71)) : ({wire7, (7'h45), reg41} <= wire1))) ?
                  $signed((&$signed((reg39 ^~ wire76)))) : {$unsigned($unsigned($signed(wire0)))});
              reg638 <= (+$unsigned((|$signed((reg634 ? reg43 : reg632)))));
            end
          else
            begin
              reg632 = reg66[(2'h3):(1'h0)];
              reg634 <= reg630;
              reg637 <= wire3;
              reg638 <= wire620[(3'h4):(1'h1)];
              reg639 <= ({$unsigned(reg630[(3'h4):(2'h3)]),
                      ($unsigned(reg61) ?
                          $signed((~^wire1)) : (reg638[(4'hb):(4'h9)] | (7'h50))),
                      ((~(~^(8'ha2))) && $unsigned($signed((8'hb0))))} ?
                  ((^(&(~&reg71))) >>> $unsigned((-reg11[(1'h1):(1'h1)]))) : reg66);
              reg640 <= reg35[(4'h8):(2'h2)];
              reg641 = $unsigned((reg52 ?
                  {(wire620 ?
                          (reg64 <<< reg47) : (~^reg35))} : (($unsigned(wire3) ?
                      ((8'ha3) ?
                          reg637 : reg625) : $signed(wire2)) ^~ ($signed(reg622) ^~ (reg639 ^ reg624)))));
            end
          for (forvar642 = (1'h0); (forvar642 < (1'h1)); forvar642 = (forvar642 + (1'h1)))
            begin
              reg643 = (-wire0);
              reg644 = (($unsigned((^(reg47 ? reg11 : wire620))) ?
                  $unsigned((~&(wire620 ?
                      (8'hba) : reg27))) : $signed($unsigned($signed(reg71)))) * ((~|reg39) ^~ (8'h9d)));
              reg645 = (((~$unsigned((forvar642 < reg637))) ?
                  $signed(((reg47 << reg27) <<< reg634)) : reg625[(2'h3):(1'h0)]) == (|(reg635 ?
                  reg61[(2'h2):(1'h0)] : $unsigned({reg13}))));
              reg646 = (reg16[(1'h1):(1'h1)] ^ ({(^(reg32 ? reg32 : reg42))} ?
                  ((~&{reg631,
                      reg41}) >= (^$signed(forvar642))) : $unsigned((&{reg635,
                      reg629,
                      reg14}))));
            end
        end
      else
        begin
          if ((-$unsigned({(^~$signed(reg34))})))
            begin
              reg622 <= $signed({reg630[(2'h3):(2'h3)],
                  {$unsigned(reg64[(5'h1a):(5'h13)]),
                      {(7'h4b), $signed(reg13), (reg631 ? forvar642 : reg16)}},
                  wire3});
              reg625 <= ({$unsigned((7'h52))} ?
                  {$unsigned($unsigned((|wire2)))} : ((&$unsigned(reg634[(1'h1):(1'h1)])) << (~^$unsigned(reg640[(2'h3):(2'h3)]))));
              reg626 <= (reg646[(5'h14):(4'hc)] ?
                  $signed(($signed(((8'h9d) << reg10)) & ((reg638 != reg49) ?
                      reg633 : $signed(wire7)))) : wire3[(5'h10):(2'h2)]);
              reg627 = ((reg634[(1'h1):(1'h0)] >> $unsigned($unsigned({reg43}))) ?
                  reg16[(2'h2):(1'h0)] : ($unsigned(({reg13,
                          (8'hb3),
                          reg633} != {reg632, (8'hb7), reg42})) ?
                      (wire4 ?
                          $signed((reg634 ? reg625 : wire3)) : (&(reg636 ?
                              reg68 : (7'h4a)))) : {$unsigned({reg46, wire1}),
                          reg623}));
              reg628 = (|($signed((8'had)) * reg637[(5'h10):(4'h9)]));
              reg629 <= reg644[(4'he):(2'h2)];
            end
          else
            begin
              reg623 = (^~(({$signed(reg36),
                      $signed(reg63),
                      (7'h44)} >= reg628) ?
                  $unsigned({$unsigned(reg624),
                      $unsigned(reg646),
                      $signed((7'h54))}) : $signed(reg637[(4'hb):(1'h0)])));
              reg624 = ((&{(wire3[(1'h0):(1'h0)] && reg629[(3'h7):(3'h5)])}) + (($unsigned((~&reg63)) != $unsigned(((8'hb1) ?
                      reg622 : reg35))) ?
                  (reg71 >= reg47) : ((8'haa) > (~reg74[(3'h5):(3'h5)]))));
              reg627 = {({({forvar627, reg16} ?
                              $unsigned(reg11) : $signed(reg638)),
                          (wire620 < {reg629})} ?
                      wire4 : ($unsigned($unsigned(reg640)) >= $unsigned((reg644 ?
                          (8'hb9) : reg35))))};
              reg628 = wire2[(1'h0):(1'h0)];
              reg630 = (~|((wire2[(3'h5):(3'h4)] ?
                      ((reg35 > reg639) != reg49[(2'h3):(1'h0)]) : reg21) ?
                  reg637 : reg635));
              reg631 <= (reg32 ? wire1 : $signed($signed({$signed((7'h44))})));
              reg632 = wire620[(5'h1a):(5'h13)];
            end
          reg633 = ($unsigned($signed($unsigned(reg623))) - $signed((8'hbb)));
          if ($signed(reg639[(1'h0):(1'h0)]))
            begin
              reg634 <= {reg630[(3'h7):(2'h3)],
                  {$signed(reg625[(1'h0):(1'h0)]), (~|(8'h9c)), $signed(reg10)},
                  wire1};
              reg637 <= reg75;
              reg638 <= ($signed(reg634[(2'h2):(2'h2)]) ?
                  reg627[(4'hf):(4'ha)] : $signed(reg16));
            end
          else
            begin
              reg635 = $unsigned((~$signed(reg75[(1'h1):(1'h0)])));
              reg636 = ($signed($unsigned(($unsigned(reg36) ~^ (&(7'h58))))) ?
                  {(~reg39), reg641[(4'hc):(3'h7)]} : (!($signed(reg638) ?
                      ({(8'hb2)} ? $signed(reg19) : reg64) : ((~|reg46) ?
                          (reg624 ^~ reg636) : (!reg644)))));
              reg637 <= {reg645[(2'h2):(1'h1)]};
              reg641 = reg633;
              reg642 <= wire76[(2'h2):(2'h2)];
              reg647 <= reg19;
              reg648 <= reg74;
            end
          for (forvar649 = (1'h0); (forvar649 < (3'h4)); forvar649 = (forvar649 + (1'h1)))
            begin
              reg650 = reg633;
              reg651 <= {((($signed(reg75) ?
                          ((8'had) >>> reg644) : reg625[(1'h0):(1'h0)]) ?
                      forvar627[(1'h0):(1'h0)] : reg637) == $signed(wire5))};
            end
          for (forvar652 = (1'h0); (forvar652 < (2'h3)); forvar652 = (forvar652 + (1'h1)))
            begin
              reg653 <= reg35[(3'h7):(1'h0)];
              reg654 <= ($signed(reg14[(4'hc):(3'h5)]) * (((reg10 ?
                  (reg58 ?
                      wire2 : reg637) : reg42[(4'hb):(2'h3)]) ^~ reg19[(5'h18):(5'h11)]) && ({reg632[(3'h6):(2'h2)],
                  (reg645 ? reg13 : reg639)} > reg647[(1'h1):(1'h1)])));
              reg655 <= reg632;
              reg656 = (&((~$signed((reg624 + reg74))) || $signed(reg46[(1'h0):(1'h0)])));
              reg657 <= $signed($signed(($unsigned($signed(reg75)) ?
                  $signed(reg647[(1'h1):(1'h0)]) : (wire0 ?
                      ((8'hbe) > reg19) : reg16[(1'h1):(1'h0)]))));
              reg658 = reg32;
              reg659 <= ($unsigned($signed((~|(reg46 + reg66)))) == ({($unsigned(reg656) ?
                          reg639[(3'h4):(2'h3)] : wire1[(2'h2):(2'h2)]),
                      reg636[(2'h2):(1'h0)]} ?
                  (~^(7'h58)) : {$signed(reg656[(1'h0):(1'h0)])}));
            end
        end
    end
  always
    @(posedge clk) begin
      reg660 <= (((((~&reg13) ?
                  wire76 : $unsigned(reg637)) >= $unsigned({reg13})) ?
              $unsigned(($signed(wire620) >> reg75)) : reg13[(1'h0):(1'h0)]) ?
          $signed({({reg622, reg642} >= (^~reg47)),
              (reg16 ?
                  reg36[(1'h1):(1'h0)] : reg71[(2'h3):(1'h1)])}) : reg46[(3'h5):(2'h3)]);
      reg661 = (^(~reg58));
      reg662 <= (|reg659);
    end
  assign wire663 = (~|(reg14 & reg11));
  always
    @(posedge clk) begin
      reg664 <= $signed(reg43[(4'h8):(3'h6)]);
      reg665 <= wire620;
    end
  always
    @(posedge clk) begin
      if ($unsigned((~|($signed({reg648}) | (~|(reg19 ? reg42 : reg625))))))
        begin
          if (($signed($unsigned((reg74[(2'h3):(2'h3)] ?
              reg11[(1'h1):(1'h0)] : $signed(reg662)))) & (&{reg42,
              ((reg662 ? reg47 : reg625) | (reg36 == reg19))})))
            begin
              reg666 = ((^((~^reg655) >= wire663[(4'ha):(3'h6)])) >= $signed((~^reg634[(2'h2):(1'h1)])));
              reg667 <= reg21;
              reg668 <= reg14;
              reg669 = ($unsigned(wire2) - $unsigned((($signed(reg49) * ((7'h4e) ?
                      (7'h41) : (8'ha7))) ?
                  (~&$signed(reg66)) : $signed((reg651 ? reg42 : reg10)))));
              reg670 <= wire7;
              reg671 = $signed($signed({(7'h42), reg642}));
            end
          else
            begin
              reg666 = ({(reg671 ?
                          {(|(8'hb2)),
                              reg11[(1'h1):(1'h0)]} : $unsigned((^~reg655)))} ?
                  $signed((7'h56)) : {{(8'ha3)}});
              reg669 = (~&wire76);
              reg670 <= $signed((&($unsigned($signed(reg16)) + reg631)));
            end
          if (reg42[(3'h6):(2'h3)])
            begin
              reg672 <= reg68[(4'hc):(1'h0)];
              reg673 = (-$signed(reg19[(3'h7):(1'h1)]));
              reg674 <= reg659[(1'h0):(1'h0)];
              reg675 <= $unsigned((~|{$signed($unsigned(reg622)),
                  ($unsigned((8'hb4)) ?
                      (^reg639) : (reg66 ? reg655 : (7'h46)))}));
            end
          else
            begin
              reg673 = reg654[(4'hb):(1'h1)];
            end
          for (forvar676 = (1'h0); (forvar676 < (2'h2)); forvar676 = (forvar676 + (1'h1)))
            begin
              reg677 <= {((~((8'hb5) ?
                          (reg640 || wire663) : (reg42 >> reg16))) ?
                      reg47 : reg64),
                  $unsigned(reg634[(1'h0):(1'h0)]),
                  $signed($signed(((reg25 == reg626) >> {wire3})))};
              reg678 <= ((^~$unsigned(((reg670 * reg11) ?
                  reg668 : (reg673 ? reg648 : (8'hb5))))) + reg651);
              reg679 <= (reg21[(4'he):(2'h2)] ?
                  ({((wire5 ? wire6 : reg654) ?
                              (^reg25) : reg25[(5'h17):(4'h8)]),
                          ((+(7'h48)) | (reg625 ? wire620 : reg648)),
                          (&reg675[(4'hf):(2'h2)])} ?
                      (^~$unsigned((wire2 + reg672))) : reg651[(1'h1):(1'h0)]) : reg43);
              reg680 = ($unsigned(wire6[(1'h0):(1'h0)]) + {$signed(reg10)});
              reg681 <= (~$unsigned(reg680));
              reg682 <= (forvar676 ?
                  (~|$unsigned((-wire620))) : (+$unsigned($unsigned((reg47 ?
                      wire0 : wire663)))));
              reg683 <= $signed(reg671[(3'h4):(2'h2)]);
            end
          if ($unsigned({(^~(8'hb9)),
              reg625[(1'h1):(1'h1)],
              (reg625 != reg11[(2'h3):(2'h3)])}))
            begin
              reg684 <= ((reg43[(1'h1):(1'h1)] ?
                      (((reg19 ^~ reg75) | $unsigned((8'hb1))) >>> $signed((reg25 ?
                          reg664 : (8'hbe)))) : (~^reg52)) ?
                  reg74[(5'h15):(4'hb)] : (~&$unsigned({$signed(reg46)})));
              reg685 <= $signed((~|((~^reg75[(2'h2):(2'h2)]) ?
                  ((&reg46) > $signed(reg68)) : ((reg41 ?
                      (7'h54) : wire0) && (wire3 << reg58)))));
              reg686 <= reg659[(2'h2):(2'h2)];
              reg687 = (^((reg657[(1'h1):(1'h0)] ?
                  (~|(~|reg52)) : ((reg686 ? reg662 : reg631) ?
                      reg25 : (reg684 << reg648))) && (((~reg74) ^ $unsigned(reg683)) == (~|(wire620 && wire5)))));
              reg688 = (((((reg52 ? reg637 : reg679) ?
                      $signed(reg66) : $signed(reg680)) || ({reg34,
                      reg678} >> $unsigned((8'haa)))) ^ $unsigned((reg35[(3'h6):(3'h4)] ^ $signed((7'h50))))) ?
                  $unsigned(wire3) : $unsigned(reg648));
              reg689 = reg13[(1'h1):(1'h0)];
              reg690 = (~reg19);
            end
          else
            begin
              reg684 <= (((reg668[(4'h8):(3'h4)] >= ($unsigned(reg678) ?
                      reg673 : reg651[(1'h0):(1'h0)])) ?
                  (((reg664 ? reg74 : wire620) & (+reg689)) ?
                      $unsigned(((8'ha1) ?
                          (8'hb5) : reg622)) : reg690) : reg75[(4'hd):(4'hd)]) ^ reg690[(1'h0):(1'h0)]);
            end
        end
      else
        begin
          reg667 <= (!$unsigned($unsigned($unsigned($unsigned((8'h9f))))));
          reg668 <= reg684[(3'h5):(1'h1)];
        end
      reg691 <= (reg41[(5'h11):(4'he)] || {$signed({$unsigned(reg671)})});
      for (forvar692 = (1'h0); (forvar692 < (3'h6)); forvar692 = (forvar692 + (1'h1)))
        begin
          if (reg664[(1'h1):(1'h1)])
            begin
              reg693 = reg25;
              reg694 <= {$signed(reg25), $signed(reg64[(5'h1a):(4'hb)])};
              reg695 = (reg43 ?
                  $signed((^~reg625[(1'h1):(1'h0)])) : ($signed(wire7[(3'h4):(2'h3)]) < (^(reg10 ?
                      $signed(wire3) : wire76))));
              reg696 = $signed($signed($signed($unsigned((^reg655)))));
            end
          else
            begin
              reg694 <= ($unsigned((reg49[(3'h5):(2'h3)] <= {$signed(reg640),
                  reg664,
                  (reg681 & wire3)})) << ({reg688[(3'h7):(2'h2)],
                      reg693[(2'h2):(1'h0)],
                      (reg696 & (reg36 ? reg637 : wire663))} ?
                  (forvar676 ?
                      (reg674 || $signed(reg61)) : $signed((reg629 ?
                          reg648 : reg648))) : (~reg42)));
              reg697 <= (+$unsigned((|$signed(reg675[(5'h18):(4'he)]))));
              reg698 = (!$signed((|(reg27 ?
                  $signed(reg691) : $signed((7'h40))))));
              reg699 = $unsigned((reg19 ?
                  ($unsigned($unsigned(reg64)) < (~^reg654)) : reg680));
              reg700 <= ((~&{reg662,
                  reg21[(5'h12):(5'h12)]}) >= (reg657 ^ ($unsigned({reg639}) ?
                  reg647 : {reg662[(4'h9):(2'h3)],
                      $signed(reg698),
                      ((7'h4e) && reg35)})));
            end
          reg701 <= $unsigned($unsigned(reg684));
          if ($signed({reg74,
              reg16[(1'h0):(1'h0)],
              ($unsigned(((8'h9d) != reg626)) ?
                  $signed((~|wire663)) : reg659[(1'h0):(1'h0)])}))
            begin
              reg702 = (~^$signed((((~&reg651) ?
                      (reg688 <= reg684) : reg52[(1'h1):(1'h0)]) ?
                  $unsigned({reg39, reg678, reg667}) : (reg660 ?
                      {reg674} : $unsigned(reg688)))));
              reg703 = $unsigned(reg700);
              reg704 <= (reg684 + $signed(reg654[(4'hd):(2'h3)]));
              reg705 = ((~|$signed((wire6 ?
                  reg75[(2'h2):(1'h1)] : {reg702,
                      reg689}))) ~^ $unsigned(({reg689, reg71} ?
                  $signed(reg10[(3'h4):(1'h0)]) : reg686)));
              reg706 = $signed((~&($unsigned($unsigned(reg629)) ?
                  $signed((reg10 ? wire1 : reg68)) : {{reg63},
                      $signed(reg622)})));
              reg707 = $unsigned($signed((reg637[(1'h0):(1'h0)] == (7'h53))));
            end
          else
            begin
              reg702 = (((7'h52) ?
                      (^~{{(8'hb6), reg678, reg679},
                          wire2}) : $unsigned((~reg684))) ?
                  $unsigned((reg651 != $signed({reg11}))) : (reg631[(2'h2):(1'h1)] ?
                      reg642[(1'h1):(1'h0)] : (!$signed(reg672[(4'h9):(2'h2)]))));
              reg704 <= (reg701 ?
                  ($signed(((~^reg625) <= (-reg74))) < reg695[(1'h1):(1'h0)]) : (reg680[(3'h7):(3'h6)] << {(+(reg685 ?
                          reg25 : reg664))}));
              reg705 = (7'h52);
              reg708 <= reg698;
            end
          for (forvar709 = (1'h0); (forvar709 < (1'h0)); forvar709 = (forvar709 + (1'h1)))
            begin
              reg710 = (reg71 ?
                  {reg638[(4'hf):(4'hc)],
                      $unsigned(wire4[(5'h15):(1'h1)]),
                      ((wire3[(1'h0):(1'h0)] ? reg629 : forvar692) ?
                          (|(~^reg697)) : $unsigned({reg46,
                              reg689}))} : ({reg668} ?
                      (8'ha5) : $signed({(&reg699), (~reg46)})));
            end
          reg711 = reg708[(5'h14):(5'h11)];
          reg712 <= reg662[(5'h10):(4'ha)];
          for (forvar713 = (1'h0); (forvar713 < (1'h1)); forvar713 = (forvar713 + (1'h1)))
            begin
              reg714 <= (^~{(~|((reg46 > reg75) & ((7'h54) <<< reg673))),
                  ((~|reg671) ?
                      (reg699[(5'h14):(2'h2)] ?
                          (reg626 <= reg14) : (reg21 * reg706)) : (~&(^reg42))),
                  $unsigned($signed(reg707[(3'h4):(2'h3)]))});
              reg715 <= $signed(reg682);
              reg716 = ($unsigned(($unsigned((wire0 ? (8'hb7) : reg36)) ?
                  $signed((reg679 ^~ reg703)) : (!reg666))) || $unsigned($unsigned((-(reg653 ?
                  reg25 : (8'hac))))));
              reg717 <= ({(-((!reg667) ?
                      reg16 : (^reg662)))} | ({reg662[(5'h18):(1'h1)],
                  ($signed(reg667) * (^~reg699)),
                  (reg66[(2'h2):(1'h1)] ?
                      $unsigned(reg694) : (+reg699))} && ($unsigned({reg675,
                      reg682}) ?
                  ({reg27} | (reg697 * reg689)) : (~^(reg16 ?
                      reg682 : reg19)))));
              reg718 = (^~reg35);
              reg719 <= (reg701[(1'h1):(1'h0)] >>> reg659[(2'h2):(1'h1)]);
            end
        end
      for (forvar720 = (1'h0); (forvar720 < (1'h0)); forvar720 = (forvar720 + (1'h1)))
        begin
          reg721 = (reg674[(1'h0):(1'h0)] ?
              reg683 : ((reg685 + reg653) ?
                  $signed($unsigned(reg21)) : wire620));
          if ({(~&{(-(reg688 ^ reg703))}),
              ({$unsigned($signed(reg52)),
                  reg679,
                  $unsigned($unsigned((7'h51)))} < (reg32 + (~^forvar720)))})
            begin
              reg722 = $signed($unsigned((-((reg11 - reg708) ?
                  reg674[(3'h7):(3'h5)] : $unsigned(wire620)))));
              reg723 = ((-$unsigned(((reg16 >= (7'h45)) ^ (^~(7'h54))))) ?
                  ({((^reg682) <<< (reg674 | (7'h4a))),
                      $unsigned((|wire5))} >= (+$unsigned(reg693[(1'h1):(1'h1)]))) : reg21[(5'h10):(4'ha)]);
              reg724 = reg631;
              reg725 = (+$unsigned(forvar713));
              reg726 <= ($unsigned(((~reg629[(3'h4):(3'h4)]) ?
                  ($unsigned(reg16) - (reg689 && wire620)) : reg651[(1'h1):(1'h1)])) ^ {(~&(~reg631)),
                  (~|reg670)});
              reg727 <= reg677[(5'h15):(4'he)];
            end
          else
            begin
              reg722 = (^$unsigned(reg693[(2'h3):(2'h3)]));
              reg726 <= reg725;
              reg727 <= $signed(((~((7'h49) << $signed(reg669))) ?
                  (~|reg654[(2'h2):(1'h1)]) : (((+reg41) ?
                          reg647 : reg36[(1'h0):(1'h0)]) ?
                      $unsigned({(7'h55)}) : (~|reg703[(2'h3):(1'h0)]))));
              reg728 <= ({$unsigned($unsigned($signed(reg694)))} <= (7'h45));
              reg729 = wire6;
              reg730 = (^~reg711[(4'he):(3'h4)]);
              reg731 = $unsigned((reg16 - (+($unsigned(reg688) ?
                  reg42[(3'h7):(3'h4)] : ((7'h4b) ? reg688 : reg680)))));
            end
          if ($unsigned(($unsigned(reg729[(5'h19):(5'h19)]) & (reg689 ?
              {(wire2 ~^ reg672)} : ($unsigned(reg711) ^ ((8'hac) - reg647))))))
            begin
              reg732 = reg672[(4'he):(2'h2)];
              reg733 <= (-reg678[(3'h6):(1'h0)]);
              reg734 <= ($signed(reg712) + ($signed(reg710[(1'h0):(1'h0)]) > reg691[(4'h8):(4'h8)]));
              reg735 = ({$unsigned(((8'h9d) ? (~&reg35) : $unsigned(reg681))),
                      $unsigned((~(reg689 ^~ forvar676)))} ?
                  ((+reg46) ?
                      (reg634[(1'h1):(1'h0)] ?
                          ($signed(reg39) ?
                              $signed(wire0) : (~^reg721)) : $signed($signed(reg669))) : (7'h54)) : (((reg35 ?
                          reg49 : reg727) ?
                      $unsigned(((8'hac) | reg691)) : ($signed(reg679) ?
                          (reg19 ?
                              reg703 : reg25) : {reg25})) <<< reg27[(3'h7):(2'h3)]));
              reg736 <= ($unsigned((8'ha1)) | {$signed((!(reg648 == reg640))),
                  ((+$unsigned(reg58)) <= $unsigned((~|reg32)))});
              reg737 <= $signed(forvar709[(1'h1):(1'h0)]);
              reg738 <= reg686;
            end
          else
            begin
              reg732 = $unsigned($signed($unsigned($signed((reg671 ^ reg694)))));
            end
          reg739 = (((reg642[(3'h6):(3'h6)] ?
                  {reg669[(4'h9):(2'h3)],
                      $unsigned(reg14),
                      $signed(reg49)} : reg699) ?
              (~^(reg712 ?
                  (~reg647) : (reg732 ?
                      (7'h50) : (7'h42)))) : wire5) <<< ((&reg41[(4'hb):(3'h7)]) ^ $unsigned(reg669)));
          for (forvar740 = (1'h0); (forvar740 < (3'h6)); forvar740 = (forvar740 + (1'h1)))
            begin
              reg741 = (reg16 ?
                  $unsigned($unsigned(reg625[(3'h5):(1'h0)])) : (({$signed(reg703),
                      $unsigned(wire4)} ^~ (reg693[(1'h0):(1'h0)] ^~ reg719[(1'h1):(1'h0)])) * $signed($signed($unsigned(reg736)))));
              reg742 <= reg678;
              reg743 <= reg36[(1'h1):(1'h0)];
              reg744 = (~|(($unsigned((reg732 >> (8'ha4))) & reg64) || $signed($unsigned((~reg698)))));
              reg745 <= reg737[(5'h19):(3'h7)];
              reg746 = $signed((^~reg10[(1'h1):(1'h0)]));
              reg747 = (!$unsigned(reg43[(3'h5):(2'h2)]));
            end
          for (forvar748 = (1'h0); (forvar748 < (3'h4)); forvar748 = (forvar748 + (1'h1)))
            begin
              reg749 = ($unsigned({(7'h4a), wire4}) ?
                  ({$unsigned((reg691 ? reg675 : reg733)),
                          {reg16[(1'h0):(1'h0)], (~|wire3)}} ?
                      (~&$signed((reg25 <= reg716))) : ({$signed(reg739),
                              $unsigned(reg729),
                              ((7'h48) * reg706)} ?
                          {(reg664 ?
                                  wire2 : (8'hbf))} : $unsigned(reg680))) : wire4);
              reg750 <= reg701[(3'h4):(1'h0)];
              reg751 <= $unsigned((^reg52[(5'h1c):(5'h17)]));
              reg752 = $signed($unsigned(reg727[(1'h0):(1'h0)]));
              reg753 <= ((|($unsigned($unsigned(reg718)) >= (7'h4c))) >= ((~^$unsigned($unsigned(reg745))) ?
                  {$signed({reg11, wire4})} : ((reg660[(4'he):(4'hb)] & {reg738,
                          (7'h4f),
                          reg27}) ?
                      reg640[(3'h4):(1'h0)] : reg672)));
            end
          if (reg668[(4'hb):(4'h8)])
            begin
              reg754 <= {reg651,
                  (reg711 ?
                      reg634[(2'h2):(2'h2)] : (($signed(reg63) ?
                              reg712[(4'hc):(3'h6)] : reg42) ?
                          ($signed(reg715) <<< $unsigned(reg13)) : $signed($unsigned(reg629)))),
                  (~&reg719[(1'h0):(1'h0)])};
              reg755 = ($unsigned(reg678[(4'he):(4'hd)]) ?
                  (reg715[(1'h1):(1'h0)] ?
                      (~|$signed((reg39 >> forvar748))) : ($signed(reg682[(3'h5):(2'h2)]) ?
                          $unsigned($unsigned(reg689)) : ($signed(forvar720) ?
                              (reg684 << reg742) : reg637))) : ($unsigned(wire2[(3'h4):(1'h1)]) ?
                      ($unsigned($unsigned(reg714)) <= $signed($signed(reg691))) : {(-reg718[(3'h4):(1'h1)]),
                          reg639[(4'he):(2'h3)],
                          (~reg75[(4'hd):(2'h2)])}));
            end
          else
            begin
              reg755 = (8'ha8);
              reg756 <= ((reg678[(3'h4):(2'h2)] ?
                  ((|reg640[(1'h0):(1'h0)]) < {$signed(reg721),
                      reg678}) : (~|reg731[(2'h2):(2'h2)])) ^~ $signed(((reg39[(2'h3):(2'h2)] ?
                  {reg68} : reg735[(5'h12):(4'hc)]) ^~ wire3[(5'h12):(4'he)])));
              reg757 = $signed(reg683[(5'h1c):(5'h1a)]);
            end
        end
      reg758 <= (({({reg739, forvar692, reg688} ? (~^(7'h4b)) : (|reg728)),
              $unsigned(reg655),
              ($unsigned(reg699) ? reg684 : $signed(reg675))} ?
          {(reg634[(2'h2):(1'h0)] < (reg16 ? forvar676 : wire2)),
              $signed(reg727[(1'h0):(1'h0)])} : $unsigned((reg684 ?
              (reg66 >> wire2) : (reg728 ~^ reg696)))) ^ ($signed(reg737[(5'h11):(3'h4)]) ?
          ((^~(reg746 ?
              (7'h49) : reg723)) <<< (reg58 <= reg671)) : reg693[(2'h3):(1'h1)]));
      reg759 <= (reg52[(1'h0):(1'h0)] ? reg712 : $unsigned($unsigned(reg743)));
    end
  always
    @(posedge clk) begin
      reg760 = (^~(7'h46));
    end
  always
    @(posedge clk) begin
      reg761 <= (8'h9f);
      if ($signed(reg750))
        begin
          reg762 <= (^~$unsigned(reg19));
        end
      else
        begin
          for (forvar762 = (1'h0); (forvar762 < (2'h2)); forvar762 = (forvar762 + (1'h1)))
            begin
              reg763 <= ((+$signed($signed(reg71[(4'ha):(3'h4)]))) ?
                  ($signed(reg728) | ($unsigned(reg655[(1'h0):(1'h0)]) ?
                      $unsigned((reg75 <= reg712)) : ((reg631 ?
                              reg701 : reg678) ?
                          $unsigned(reg662) : reg42[(4'hd):(1'h1)]))) : $unsigned({reg75[(4'hb):(4'hb)]}));
              reg764 <= $unsigned($signed((reg681 > $signed($unsigned(reg684)))));
              reg765 = reg763;
              reg766 <= ((|((+((8'ha4) || forvar762)) > ($signed(reg647) ?
                      $signed(reg651) : (-reg742)))) ?
                  $signed(((((7'h40) ? reg660 : wire3) | (reg700 ?
                          reg667 : (7'h49))) ?
                      reg68[(4'h8):(3'h4)] : (~|(wire7 && reg642)))) : (wire7[(4'hf):(4'hb)] ?
                      ($signed(reg634[(2'h3):(1'h1)]) ^~ reg10[(2'h3):(1'h0)]) : reg43));
              reg767 = $unsigned(reg765);
              reg768 = {reg16,
                  (^(reg47 ?
                      reg625[(2'h2):(1'h0)] : $unsigned((reg678 >> wire5)))),
                  (((^(reg762 ^ reg668)) <<< (+(^reg64))) ?
                      $unsigned(reg756) : $unsigned($signed((reg634 <<< reg665))))};
              reg769 = $unsigned(wire76);
            end
          reg770 = $unsigned(reg626[(4'hd):(2'h2)]);
        end
      if ({(~|$unsigned(reg717)),
          $unsigned((reg27 << ((reg736 & reg679) ?
              (wire4 ? reg737 : reg58) : $unsigned(reg762)))),
          $signed($unsigned(reg761))})
        begin
          for (forvar771 = (1'h0); (forvar771 < (3'h4)); forvar771 = (forvar771 + (1'h1)))
            begin
              reg772 = ((&$unsigned($signed({reg41, reg41}))) ?
                  (($signed((~^reg677)) ?
                          ((reg742 * reg683) ~^ reg657[(1'h0):(1'h0)]) : reg665[(4'h8):(3'h7)]) ?
                      wire76 : reg742) : (((reg631 ?
                      (reg719 - reg742) : reg631) - {(reg16 > reg25),
                      reg14[(4'hd):(3'h6)]}) == reg756[(3'h6):(3'h4)]));
              reg773 = $unsigned(reg49[(3'h5):(3'h4)]);
              reg774 <= (({$unsigned((reg41 + reg74)),
                          {((8'hb7) ? reg679 : wire1)},
                          {wire6[(1'h0):(1'h0)]}} ?
                      $unsigned((!$unsigned((7'h48)))) : $signed(($signed(reg764) ?
                          reg758[(2'h2):(1'h0)] : reg759))) ?
                  reg745 : {$unsigned(((wire76 != reg701) ?
                          (reg19 <= wire6) : reg68)),
                      (~^reg717)});
              reg775 = reg664;
              reg776 = $signed($unsigned(reg13));
              reg777 <= $signed({$signed($unsigned(((8'hb2) <<< reg704))),
                  reg34[(2'h3):(1'h1)]});
            end
          if ($signed(reg772[(2'h2):(1'h0)]))
            begin
              reg778 <= (reg657 ?
                  (-reg678[(5'h12):(4'he)]) : (&$signed(reg639)));
              reg779 = reg66;
            end
          else
            begin
              reg779 = ((~^(wire620[(3'h5):(3'h5)] ?
                  (7'h4d) : $unsigned({reg61, reg761, wire2}))) < reg774);
              reg780 = (8'hb5);
              reg781 <= $signed((reg13 ^~ (reg43 * ({reg36} >> (reg679 << wire0)))));
              reg782 <= $signed(((7'h49) & reg32[(1'h1):(1'h1)]));
              reg783 <= reg727;
            end
          reg784 <= reg768[(5'h12):(4'hd)];
          reg785 = $unsigned($unsigned($signed($signed(reg754))));
          for (forvar786 = (1'h0); (forvar786 < (3'h5)); forvar786 = (forvar786 + (1'h1)))
            begin
              reg787 = (reg631 ? {$signed(reg768)} : $signed(reg777));
              reg788 <= {(!{reg58})};
              reg789 = ((reg670 + $signed((+(reg783 ?
                  reg68 : reg694)))) >> $unsigned(reg719[(1'h1):(1'h0)]));
              reg790 = reg63;
              reg791 = (reg681 <= (((~&((7'h4f) || reg670)) * (~|(~reg719))) >>> reg647[(3'h5):(3'h5)]));
              reg792 <= (+$unsigned((^~{$unsigned(reg43)})));
            end
        end
      else
        begin
          reg771 <= reg651;
          if ((reg766[(3'h4):(2'h2)] >= ((reg639[(1'h1):(1'h1)] <<< ((reg668 ?
                  reg719 : (8'ha5)) ?
              (-reg14) : {wire663, reg761, reg39})) - reg753)))
            begin
              reg772 = ($unsigned($signed(reg697[(3'h5):(2'h2)])) <= (($unsigned($signed((8'hb0))) ?
                      (~&$signed(wire0)) : ((~reg640) ~^ (reg764 && reg717))) ?
                  (($signed(reg681) ?
                      (!reg625) : (reg679 ?
                          reg770 : reg659)) ~^ {reg785[(3'h5):(1'h1)],
                      {reg46},
                      $signed(reg790)}) : $unsigned(reg763)));
              reg773 = ($signed((~reg753[(1'h0):(1'h0)])) ^ reg784);
            end
          else
            begin
              reg772 = reg758;
              reg773 = (|($signed((|(8'h9e))) >>> $signed($signed((reg651 != reg638)))));
              reg774 <= reg622;
            end
          if (wire76)
            begin
              reg777 <= reg691[(3'h7):(3'h4)];
              reg779 = reg736[(5'h11):(5'h10)];
              reg781 <= (-reg659);
            end
          else
            begin
              reg775 = reg767;
              reg776 = $unsigned(((&($unsigned(reg765) << $signed(reg766))) != (~&((reg657 - (8'ha2)) ?
                  reg682[(4'h9):(2'h2)] : reg765))));
              reg779 = forvar771[(4'he):(3'h4)];
              reg780 = reg10[(2'h2):(1'h1)];
            end
          reg782 <= (+$signed($signed(reg681)));
          if (forvar771)
            begin
              reg785 = $unsigned(({$signed($unsigned(reg664)),
                      $signed((reg653 ? reg792 : reg672))} ?
                  ($unsigned(((8'ha4) ? wire620 : reg701)) ?
                      ((reg742 ? wire620 : reg704) << {forvar786,
                          reg667,
                          reg785}) : {reg742,
                          {reg791, reg41},
                          reg653[(2'h3):(1'h0)]}) : ($unsigned($signed(reg694)) ?
                      reg622[(4'ha):(1'h1)] : (8'h9c))));
              reg786 <= (8'hb7);
              reg787 = {{$unsigned(reg625),
                      $unsigned({$signed(reg13)}),
                      ((-$signed((7'h53))) != {$signed(reg684)})},
                  $signed(reg677[(5'h16):(4'ha)]),
                  (~&$unsigned($unsigned(reg42[(5'h14):(3'h7)])))};
              reg789 = (reg648[(4'h9):(4'h9)] && reg763);
              reg790 = $signed($unsigned((reg642[(4'h8):(3'h6)] ^~ (^~$signed(wire663)))));
              reg792 <= reg781;
              reg793 <= reg682[(4'hd):(2'h3)];
            end
          else
            begin
              reg783 <= $signed($signed(reg634[(2'h2):(2'h2)]));
              reg785 = $unsigned(reg43);
              reg786 <= ((reg14 ?
                      reg13 : ({reg773[(2'h2):(2'h2)],
                              {reg634, reg750, reg14},
                              (reg769 ? wire4 : wire620)} ?
                          ((wire5 != reg68) ?
                              $unsigned(reg63) : $unsigned(reg783)) : ((reg659 ?
                                  (7'h44) : reg779) ?
                              reg733[(3'h4):(1'h0)] : ((8'h9c) ?
                                  reg61 : reg770)))) ?
                  (^($unsigned($unsigned(reg670)) ?
                      $unsigned((+reg779)) : reg737)) : (^(&$unsigned($signed(reg785)))));
              reg788 <= (reg751[(3'h6):(3'h6)] || (reg659 ?
                  reg785[(3'h7):(3'h4)] : reg762));
              reg789 = $unsigned($unsigned(({$unsigned(reg764)} ?
                  $signed(wire7[(4'ha):(2'h3)]) : forvar786[(1'h0):(1'h0)])));
            end
          reg794 <= reg717;
        end
      reg795 <= $unsigned($signed({(^wire0),
          (~(~^reg794)),
          reg43[(2'h3):(2'h2)]}));
      reg796 = $unsigned((~((&{reg790, reg701, wire663}) ?
          (7'h57) : (!(reg679 ? wire4 : reg785)))));
      reg797 = reg679;
    end
  always
    @(posedge clk) begin
      for (forvar798 = (1'h0); (forvar798 < (2'h2)); forvar798 = (forvar798 + (1'h1)))
        begin
          if (reg651[(3'h6):(3'h5)])
            begin
              reg799 = {$unsigned((({reg648, reg657} ?
                          ((8'hb4) & reg794) : $signed(reg32)) ?
                      reg625 : reg637[(4'h9):(3'h7)]))};
              reg800 = (8'h9d);
              reg801 <= (+($unsigned($unsigned($signed(reg784))) && (reg686[(2'h2):(1'h0)] ?
                  reg675[(3'h5):(2'h3)] : ({reg734} ?
                      $signed(reg783) : $unsigned(reg737)))));
              reg802 = (|({reg733[(5'h12):(1'h0)]} ?
                  reg47[(1'h1):(1'h1)] : (|(&(reg788 >> reg758)))));
              reg803 <= {({((~|wire2) ? $signed(reg672) : $unsigned(reg783))} ?
                      reg36 : {reg717, reg664})};
              reg804 <= (!{reg686[(3'h6):(3'h4)],
                  reg751,
                  (^~(^((8'ha3) > reg670)))});
              reg805 = reg792[(3'h4):(1'h1)];
            end
          else
            begin
              reg799 = $signed({($signed((reg793 ? reg743 : reg637)) ?
                      (wire1 || (~reg675)) : (^~(8'ha8)))});
              reg800 = $unsigned((reg794 ?
                  (($unsigned(reg762) ^ (~|(7'h54))) >>> (|(reg737 ?
                      wire7 : reg782))) : ($signed((reg756 ~^ (7'h45))) ?
                      (|(reg41 + reg804)) : ((reg784 ? reg700 : wire3) ?
                          {reg804} : ((8'haf) | (7'h4c))))));
            end
          if ($unsigned(reg14[(4'hc):(4'hc)]))
            begin
              reg806 = $signed((((reg800[(5'h13):(4'hb)] ?
                          $signed((8'hb2)) : (reg766 ^~ reg677)) ?
                      reg697 : (~|(8'h9f))) ?
                  {(~&$unsigned(reg622))} : reg675[(4'hf):(1'h0)]));
              reg807 <= ({{($unsigned(reg762) & (~reg762)),
                      reg701[(2'h3):(2'h2)]}} < ($unsigned(($signed(reg715) ?
                      reg738[(3'h5):(2'h2)] : (reg49 ^ reg737))) ?
                  reg640[(3'h7):(1'h1)] : (&((~&reg753) ? reg16 : (+reg786)))));
              reg808 <= (($unsigned(reg27[(3'h7):(1'h1)]) ?
                      $unsigned((wire76[(2'h2):(2'h2)] ?
                          (reg677 ?
                              reg726 : reg660) : (~^wire5))) : $signed($signed((~|reg32)))) ?
                  reg670[(1'h1):(1'h1)] : (reg21[(4'hd):(4'hd)] ?
                      (^($signed(reg784) * $signed(reg41))) : ($unsigned(reg781[(5'h10):(3'h5)]) ?
                          $signed(reg782) : ($unsigned(reg795) <<< reg788))));
              reg809 = (~^((&reg651[(1'h1):(1'h1)]) ?
                  reg712 : $signed(((~&reg700) ? (|reg46) : (^reg719)))));
              reg810 = $signed((($signed((reg653 || reg677)) * $unsigned(((8'ha4) ?
                      reg74 : reg675))) ?
                  ($signed($unsigned(reg777)) ?
                      ($signed(reg14) > (reg16 || reg758)) : $unsigned(reg64)) : $signed($unsigned((reg66 ?
                      reg677 : (7'h4c))))));
              reg811 <= (reg16[(2'h2):(1'h0)] ^~ (!$signed({(reg788 <<< reg58)})));
              reg812 = reg659;
            end
          else
            begin
              reg806 = ((&$unsigned(((-reg812) ? (8'ha6) : (7'h49)))) ?
                  ($signed({(reg745 || reg727), reg781, reg25}) ?
                      ((&$signed((8'haa))) & ($signed(wire76) ?
                          (~reg771) : (~|reg622))) : $signed({(8'hb7),
                          $signed(reg64),
                          (reg750 <<< reg766)})) : $unsigned($signed((!reg660))));
              reg807 <= $unsigned($unsigned(reg21[(2'h3):(1'h1)]));
              reg809 = ((^~(~^$signed((reg802 ? reg734 : reg637)))) ?
                  reg46[(1'h1):(1'h0)] : $unsigned($unsigned(reg631)));
              reg810 = (^(($signed((wire2 ? reg781 : reg737)) < {(+(7'h55)),
                  (~&reg11)}) <= $signed($signed((reg806 ? reg629 : reg637)))));
            end
          for (forvar813 = (1'h0); (forvar813 < (3'h5)); forvar813 = (forvar813 + (1'h1)))
            begin
              reg814 <= $signed(($unsigned($unsigned($unsigned(reg694))) == reg13[(1'h1):(1'h1)]));
              reg815 <= {(~^reg751[(3'h6):(1'h0)]),
                  ({{$unsigned(reg766)}, wire3} + reg58[(1'h1):(1'h0)])};
              reg816 <= $unsigned((~^(~&{$unsigned(reg759),
                  (reg13 ? reg657 : reg717)})));
            end
          if ($unsigned(($unsigned($signed({reg66})) ^ reg10)))
            begin
              reg817 <= (!(($signed({(8'hbf), reg639}) ?
                  $signed(reg52) : (~&reg727)) & $unsigned(reg75[(4'hd):(3'h7)])));
            end
          else
            begin
              reg817 <= ((8'ha6) ?
                  ((~reg46[(3'h4):(3'h4)]) + (((reg685 << reg804) - reg738[(4'h8):(3'h5)]) >>> $signed((reg808 + reg753)))) : (^~$signed((~&$signed((8'hb2))))));
              reg818 = (reg681 ?
                  {reg64,
                      reg704} : ((wire0[(2'h2):(1'h1)] >>> (^$signed((7'h49)))) ~^ $unsigned(reg677)));
            end
        end
      reg819 <= (reg670[(1'h1):(1'h1)] ?
          reg750[(4'hd):(3'h5)] : (reg648 >> reg34));
      for (forvar820 = (1'h0); (forvar820 < (3'h4)); forvar820 = (forvar820 + (1'h1)))
        begin
          for (forvar821 = (1'h0); (forvar821 < (3'h4)); forvar821 = (forvar821 + (1'h1)))
            begin
              reg822 = {$unsigned((~$unsigned(reg32[(4'hc):(3'h7)]))),
                  $unsigned(($signed(reg761[(2'h2):(2'h2)]) && ($unsigned(forvar813) ?
                      reg766[(2'h2):(1'h0)] : reg27)))};
            end
          reg823 = reg784;
          reg824 = {(($unsigned((reg66 - reg812)) < reg19) ^~ $unsigned(wire0)),
              reg778[(5'h13):(4'hd)],
              {$unsigned(reg694),
                  reg818,
                  $unsigned($signed((reg704 >>> reg810)))}};
          reg825 = {$unsigned($unsigned(({wire1} ^ (reg66 >> (8'hbe))))),
              ($unsigned((reg737[(4'he):(2'h3)] && $unsigned(reg14))) | (($unsigned((7'h4c)) - (^reg809)) ?
                  reg805 : reg66))};
          for (forvar826 = (1'h0); (forvar826 < (2'h2)); forvar826 = (forvar826 + (1'h1)))
            begin
              reg827 = $signed({(^reg762[(3'h7):(3'h6)])});
              reg828 = (reg771[(5'h10):(2'h3)] ?
                  $signed((((~^reg777) == $signed((8'hb4))) >= (&(reg734 + reg701)))) : ((reg61[(4'hc):(4'h8)] ?
                          reg75[(3'h4):(3'h4)] : ({reg670,
                              reg714,
                              reg808} > (reg805 ^~ reg774))) ?
                      wire4[(5'h12):(2'h2)] : $unsigned($signed((reg733 <= reg691)))));
              reg829 = $unsigned(reg691[(4'h8):(1'h0)]);
              reg830 <= (wire4 ^~ ($signed(reg727[(2'h2):(1'h0)]) > (forvar798[(1'h0):(1'h0)] >> reg682[(3'h5):(2'h2)])));
              reg831 <= (~|$unsigned($unsigned(reg34)));
              reg832 <= reg13;
            end
          reg833 <= ((($unsigned($unsigned(reg750)) && (reg743 || reg665)) ?
                  (~&((reg659 ? forvar820 : reg761) ^~ (reg777 ?
                      wire0 : (7'h53)))) : $unsigned((7'h45))) ?
              $signed({$signed((reg816 < reg807))}) : reg63);
        end
      reg834 = (~|{reg685});
    end
  assign wire835 = ((~|reg691[(2'h2):(1'h0)]) ^ reg766[(3'h7):(3'h5)]);
  always
    @(posedge clk) begin
      reg836 = reg832;
      if ((+$signed(reg36)))
        begin
          reg837 = {$signed(reg13[(1'h0):(1'h0)]),
              ($signed($unsigned($unsigned(reg701))) > {reg36[(2'h3):(1'h1)],
                  (^~(reg622 * (7'h52))),
                  reg814[(2'h3):(2'h3)]}),
              {$unsigned(($signed(reg811) ?
                      (reg46 == reg795) : reg58[(1'h0):(1'h0)]))}};
          if ((reg793[(5'h15):(5'h11)] & reg784))
            begin
              reg838 <= $signed((-$unsigned(reg701[(1'h1):(1'h1)])));
              reg839 = $signed((reg742[(5'h18):(4'hb)] & reg764));
              reg840 = reg763;
              reg841 = reg679[(4'h8):(3'h6)];
            end
          else
            begin
              reg838 <= ({(reg19 ? reg754[(1'h0):(1'h0)] : (+wire5)),
                      $signed(reg836[(5'h18):(5'h16)]),
                      $unsigned((8'hbc))} ?
                  (^~({$signed(reg665),
                      (reg717 ?
                          reg728 : reg803)} - $signed(reg771[(4'he):(4'he)]))) : {$signed(reg840),
                      reg738[(3'h4):(2'h2)]});
              reg839 = $signed(reg781);
            end
        end
      else
        begin
          for (forvar837 = (1'h0); (forvar837 < (3'h5)); forvar837 = (forvar837 + (1'h1)))
            begin
              reg838 <= $unsigned((|$signed({{reg759}, $signed((8'h9c))})));
              reg839 = reg793[(4'h9):(3'h6)];
              reg840 = (~&{(^$unsigned(reg61[(4'ha):(2'h2)]))});
              reg841 = (($signed(reg32[(4'h8):(4'h8)]) ?
                  {reg778} : reg808) == {(reg629 | $signed($signed(reg674))),
                  ({$signed((7'h58)),
                      reg728,
                      (reg14 - reg700)} ~^ ((reg647 || reg761) - (reg819 ?
                      (8'h9c) : reg675)))});
              reg842 <= $unsigned((7'h40));
              reg843 <= (((!reg66) ^~ reg674[(3'h6):(3'h5)]) <<< reg762);
            end
          reg844 <= $signed(reg35[(4'hd):(2'h2)]);
          reg845 <= $signed(((~&({(7'h48)} ?
              $signed(reg41) : (reg667 * reg657))) == ($signed(((8'ha9) ?
              reg701 : reg701)) <= reg39[(3'h5):(3'h5)])));
          if (reg801)
            begin
              reg846 <= {$unsigned(reg764), wire1[(3'h4):(2'h2)]};
              reg847 <= (+reg846);
              reg848 <= reg839;
            end
          else
            begin
              reg846 <= {reg736};
              reg847 <= {(&reg74[(5'h1c):(5'h14)])};
              reg848 <= (((+(reg42 >= $unsigned(reg642))) ?
                  reg637 : $signed(wire5)) != (reg626 + ($unsigned((^wire7)) << $unsigned((wire835 ?
                  reg660 : reg32)))));
              reg849 = ($signed($unsigned($signed((reg657 ?
                  reg13 : reg817)))) ^~ (&$signed(reg734)));
              reg850 <= reg25[(5'h12):(2'h2)];
            end
        end
      reg851 = reg733[(5'h12):(3'h5)];
    end
  assign wire852 = wire663;
  assign wire853 = (8'ha1);
  assign wire854 = wire0[(1'h1):(1'h0)];
  assign wire855 = $signed($signed($unsigned({(+reg58),
                       reg659,
                       $signed(reg778)})));
  always
    @(posedge clk) begin
      reg856 = $unsigned(reg659);
      for (forvar857 = (1'h0); (forvar857 < (1'h0)); forvar857 = (forvar857 + (1'h1)))
        begin
          if (reg64[(4'he):(1'h1)])
            begin
              reg858 = (+$signed($signed(({reg686, reg634} ?
                  (reg792 ? reg19 : reg843) : reg75))));
              reg859 <= ((((reg647[(3'h5):(3'h4)] && reg808[(3'h5):(2'h3)]) ?
                      reg762 : $signed($unsigned(reg761))) ?
                  $unsigned({$signed(reg754),
                      $signed((8'ha9))}) : $signed(forvar857[(5'h16):(4'hf)])) & (~&(+((8'ha8) ?
                  reg736 : $signed(reg683)))));
            end
          else
            begin
              reg858 = {reg625, reg804[(1'h1):(1'h0)]};
              reg860 = reg719[(1'h1):(1'h1)];
              reg861 = reg778[(5'h11):(3'h4)];
            end
          for (forvar862 = (1'h0); (forvar862 < (1'h0)); forvar862 = (forvar862 + (1'h1)))
            begin
              reg863 = (($signed(reg19) ?
                      $signed(reg629[(5'h14):(4'hb)]) : $unsigned((wire76[(3'h7):(1'h1)] ?
                          reg10[(3'h4):(2'h2)] : (~reg766)))) ?
                  ({(&((8'ha5) ?
                          reg842 : forvar862))} && $signed($signed((+reg850)))) : {(&((-reg781) ~^ reg794[(3'h5):(1'h0)])),
                      {$signed((reg842 ? reg49 : reg808)),
                          (~^{(7'h47), reg691}),
                          reg784[(3'h6):(3'h5)]},
                      reg41});
              reg864 = ($signed(wire663) ?
                  reg750[(4'hc):(3'h7)] : reg860[(4'he):(2'h3)]);
            end
          reg865 = reg651[(3'h4):(1'h1)];
          for (forvar866 = (1'h0); (forvar866 < (3'h6)); forvar866 = (forvar866 + (1'h1)))
            begin
              reg867 = $signed($unsigned(reg847[(1'h1):(1'h0)]));
              reg868 <= $signed({$unsigned((+(reg778 | wire76))),
                  (reg867[(2'h2):(1'h1)] > ($signed(reg21) != $unsigned(reg71))),
                  $unsigned((^$signed(reg761)))});
              reg869 <= reg626;
              reg870 <= $unsigned(($unsigned(($unsigned(reg814) > (reg784 ^~ reg850))) >>> (+{(reg786 == reg844),
                  wire7[(3'h7):(1'h1)],
                  reg629})));
              reg871 <= forvar862[(4'hc):(2'h2)];
              reg872 <= (reg804[(4'hb):(3'h7)] ?
                  {($unsigned((reg701 ?
                          reg704 : reg674)) > ($unsigned(reg758) ^~ $unsigned(reg733)))} : (~^((7'h44) != $unsigned(reg662[(5'h1a):(5'h13)]))));
            end
          for (forvar873 = (1'h0); (forvar873 < (3'h4)); forvar873 = (forvar873 + (1'h1)))
            begin
              reg874 = reg25;
            end
          for (forvar875 = (1'h0); (forvar875 < (2'h2)); forvar875 = (forvar875 + (1'h1)))
            begin
              reg876 = reg782[(3'h4):(2'h3)];
              reg877 = $unsigned((((-$unsigned(reg728)) ?
                  ($unsigned(reg66) ^ (^~reg74)) : {$signed(reg683)}) == $unsigned(reg719)));
              reg878 = {$unsigned((forvar857[(5'h15):(3'h6)] ?
                      reg691[(3'h6):(1'h0)] : $signed((|reg801))))};
            end
        end
    end
  assign wire879 = $signed(reg794[(2'h3):(1'h0)]);
  assign wire880 = $unsigned((|reg719));
  assign wire881 = (^~($unsigned($signed($unsigned(reg764))) == (+(reg672 ?
                       $unsigned(wire1) : {reg845, reg64, reg657}))));
  always
    @(posedge clk) begin
      if (wire835)
        begin
          if (wire6)
            begin
              reg882 = $signed(reg848);
              reg883 <= ($signed(reg778[(2'h2):(2'h2)]) >> reg631);
              reg884 = $signed(reg63);
              reg885 <= $unsigned(wire663[(4'h9):(4'h9)]);
            end
          else
            begin
              reg882 = wire854[(1'h1):(1'h1)];
              reg884 = wire835;
              reg885 <= $signed($signed(reg816));
              reg886 = wire663;
              reg887 <= (reg712[(4'hc):(4'h9)] ?
                  reg872[(1'h1):(1'h0)] : $unsigned(($unsigned(wire663) ?
                      {reg804[(1'h0):(1'h0)],
                          $unsigned(reg831),
                          $signed(reg638)} : ((reg728 ?
                          wire853 : (7'h54)) | ((8'hbc) || reg846)))));
              reg888 <= $signed((7'h4d));
            end
          if ((&{{(reg846[(3'h5):(1'h0)] ? {reg742} : (reg793 >>> reg71)),
                  $unsigned(reg647)},
              reg885[(2'h2):(1'h1)]}))
            begin
              reg889 = $signed(($signed($unsigned(wire879)) * reg49));
              reg890 = reg759[(1'h0):(1'h0)];
              reg891 <= {(^$signed({$unsigned(reg838),
                      $unsigned(wire0),
                      $unsigned(reg831)})),
                  (^(-(reg817 > $unsigned(wire879))))};
            end
          else
            begin
              reg889 = $signed(reg678[(4'he):(3'h4)]);
              reg890 = (reg777[(5'h11):(4'hb)] ?
                  $signed(($signed((reg677 ? reg782 : reg728)) | ({reg743} ?
                      $signed(reg889) : (reg691 ?
                          reg782 : reg683)))) : ((reg685[(3'h4):(2'h2)] ?
                      $unsigned(reg816[(2'h3):(2'h3)]) : reg846) <<< reg811[(4'ha):(1'h1)]));
              reg892 = ((reg52[(3'h6):(2'h2)] ?
                      $unsigned($unsigned($signed(reg691))) : reg751[(2'h3):(2'h3)]) ?
                  {(~^((~|reg629) & reg662))} : reg61);
              reg893 = reg753;
              reg894 <= reg754;
              reg895 <= ((^~(|{(^reg655), {(8'ha6)}, reg10[(2'h2):(1'h1)]})) ?
                  {reg833[(3'h6):(1'h1)],
                      $unsigned(((reg893 ?
                          reg892 : reg738) <<< $signed((8'hab)))),
                      $unsigned($unsigned($unsigned((8'ha6))))} : (8'hb6));
            end
          for (forvar896 = (1'h0); (forvar896 < (1'h1)); forvar896 = (forvar896 + (1'h1)))
            begin
              reg897 = wire853[(2'h2):(2'h2)];
              reg898 = {reg47[(3'h4):(2'h3)],
                  {reg21,
                      (~^{$unsigned(reg19),
                          $unsigned(reg887),
                          (reg654 ? wire620 : reg626)}),
                      (~^$signed((reg884 ? reg850 : forvar896)))},
                  ((7'h4e) >>> $unsigned((&$signed((8'hac)))))};
              reg899 = $signed((~^(&reg58[(1'h0):(1'h0)])));
              reg900 <= (^(reg742[(5'h14):(5'h10)] ?
                  ($unsigned({(7'h52), reg25, wire5}) ?
                      reg887[(4'hf):(4'hd)] : {((8'haa) ?
                              reg52 : reg893)}) : $unsigned(($signed(reg781) ?
                      $unsigned(reg894) : (reg683 ? reg886 : reg845)))));
              reg901 <= reg694;
            end
          reg902 = (((~^($unsigned(reg764) >= reg726[(4'h9):(3'h6)])) ?
                  (&((reg786 ?
                      reg736 : reg844) || reg47[(2'h3):(1'h1)])) : ((^$signed((8'haa))) ?
                      reg678 : (reg894 ?
                          $unsigned(reg682) : reg678[(5'h12):(4'hb)]))) ?
              reg640 : reg659);
        end
      else
        begin
          reg882 = ({(8'hbc),
              (((~|reg887) ? {reg738, (8'hb3)} : reg625) ?
                  reg781[(5'h12):(5'h10)] : ($unsigned((8'had)) >> reg670[(1'h1):(1'h1)])),
              reg759[(1'h0):(1'h0)]} * reg742[(3'h7):(2'h3)]);
          reg883 <= (^~reg694);
          reg884 = ((~(~$unsigned((-(7'h56))))) ?
              $unsigned((reg898 << (((8'ha2) >>> reg758) <<< {reg674,
                  reg844,
                  (7'h42)}))) : {{{((8'ha4) ~^ reg786)}, $signed(reg665)},
                  {$signed($unsigned(reg634)),
                      ($signed(reg39) ?
                          ((7'h56) ?
                              reg784 : reg719) : wire76[(2'h3):(2'h3)])}});
          if ($unsigned($signed($signed({((8'hb1) > (8'hae)),
              reg66[(3'h5):(1'h0)],
              $signed(reg814)}))))
            begin
              reg886 = reg736[(2'h2):(2'h2)];
              reg889 = (^$unsigned({reg681, reg893}));
              reg891 <= reg891;
              reg894 <= $unsigned($signed(({$signed(wire852)} >>> {(reg71 + reg816),
                  {(8'hb9), reg626},
                  (~&reg743)})));
              reg895 <= reg691;
              reg896 = {reg25,
                  $signed((reg782[(1'h1):(1'h0)] == $unsigned((reg626 != wire853))))};
            end
          else
            begin
              reg886 = $unsigned((&(^(7'h44))));
              reg889 = $unsigned((~&(((reg870 ? (8'haa) : reg708) ^~ (reg761 ?
                  reg719 : reg788)) || reg674[(4'h8):(1'h1)])));
              reg890 = {(({((8'ha8) || (8'ha1)),
                      $unsigned(reg833)} <= reg631[(3'h6):(3'h6)]) - ({(reg883 ?
                          reg872 : wire76),
                      (reg651 ? (7'h46) : reg882),
                      reg887} ~^ ((reg733 ~^ reg647) ^ reg714[(3'h5):(2'h2)]))),
                  {(7'h57),
                      reg10,
                      (^~{$signed(reg753), $signed(reg681), (~reg683)})},
                  forvar896};
              reg892 = reg901[(3'h4):(1'h1)];
              reg894 <= $unsigned(reg727);
              reg895 <= (wire854 && $signed(reg35[(4'hf):(1'h0)]));
              reg896 = {reg678[(5'h16):(1'h0)]};
            end
          if ($unsigned($signed({$unsigned((~^reg13)),
              reg63[(5'h13):(5'h11)]})))
            begin
              reg897 = (7'h46);
              reg900 <= reg759;
              reg902 = $unsigned($signed((^{(~&reg708)})));
            end
          else
            begin
              reg897 = $unsigned(wire853[(1'h1):(1'h0)]);
              reg898 = {{reg774},
                  $signed({((^~reg697) <= reg814[(2'h3):(2'h2)]),
                      reg34[(3'h4):(2'h2)]})};
              reg899 = reg14;
              reg902 = reg844;
              reg903 = reg848[(4'h8):(1'h1)];
              reg904 = (reg736[(1'h0):(1'h0)] && (+($unsigned((reg708 || reg700)) == $unsigned({reg36,
                  reg714,
                  (7'h4b)}))));
            end
          for (forvar905 = (1'h0); (forvar905 < (1'h0)); forvar905 = (forvar905 + (1'h1)))
            begin
              reg906 = ((~|($signed($signed(reg903)) > (~&$unsigned(reg792)))) | $unsigned(reg727[(2'h2):(1'h0)]));
              reg907 = $signed(reg885[(2'h3):(1'h1)]);
              reg908 <= (wire881 ? $signed(reg890) : reg647[(1'h0):(1'h0)]);
              reg909 <= ((8'hb2) ?
                  (($unsigned((reg637 ?
                      wire0 : reg870)) ^~ (^~$signed(reg734))) ^~ ($unsigned($unsigned((7'h4f))) >> reg642)) : ($signed((reg742 ?
                      (reg719 ? reg882 : (7'h4e)) : (reg678 ?
                          reg694 : reg871))) <= reg651[(2'h3):(1'h1)]));
              reg910 <= {reg39[(3'h7):(3'h7)],
                  $unsigned(reg763[(3'h4):(3'h4)])};
              reg911 = reg870[(3'h6):(1'h0)];
            end
          if ($unsigned($unsigned($signed(($signed(wire5) >= $signed(reg694))))))
            begin
              reg912 <= wire852;
              reg913 = {($signed(reg762[(1'h1):(1'h1)]) <= ($unsigned(reg685) ?
                      $signed($signed(reg653)) : ((~reg662) ?
                          wire2[(1'h1):(1'h0)] : (reg778 ? reg708 : reg637)))),
                  $signed((reg788 <<< ($unsigned(reg694) ?
                      ((8'haf) + reg832) : $signed(wire663)))),
                  {(~|((reg889 & reg715) ?
                          $unsigned(reg848) : $signed(reg754))),
                      {reg651[(1'h0):(1'h0)],
                          (~|(reg766 * (8'ha0))),
                          ((&reg75) ? $signed(reg869) : $signed(reg870))},
                      ($signed(((7'h4d) & reg46)) >= ({(7'h43), reg750, wire0} ?
                          (reg833 ^~ reg788) : reg714[(4'h8):(2'h2)]))}};
              reg914 = $unsigned(reg68[(4'he):(2'h2)]);
              reg915 = (($unsigned((!reg715)) ?
                  (|{$unsigned(reg886), $signed(reg648)}) : {$unsigned(reg794),
                      reg654}) + {$unsigned((-$signed(reg814))),
                  $unsigned(reg637[(4'hc):(3'h5)])});
            end
          else
            begin
              reg912 <= (-reg36[(2'h2):(1'h0)]);
              reg916 <= (~^$unsigned((!((reg830 ?
                  reg679 : (7'h57)) ~^ reg781))));
              reg917 <= $signed(((8'ha2) ?
                  ($unsigned($signed(reg655)) ?
                      reg830[(4'hb):(3'h7)] : ((~|reg793) != (reg914 ?
                          reg884 : reg19))) : ($unsigned(((8'ha5) ?
                          reg637 : reg651)) ?
                      ((~|reg634) || $signed(reg891)) : {(8'hb3)})));
              reg918 = reg738[(4'hf):(1'h0)];
              reg919 = reg717[(4'hf):(4'hf)];
            end
        end
      reg920 <= reg904[(2'h3):(2'h2)];
      if ($signed(reg10[(3'h4):(1'h1)]))
        begin
          if ((~|{$signed((|(~reg651))), reg674[(4'h9):(3'h5)]}))
            begin
              reg921 = ((+((^$signed(reg634)) ?
                  wire852 : ((~^(7'h50)) ?
                      reg912[(4'h9):(2'h3)] : (!reg915)))) == $unsigned(reg66));
              reg922 <= (reg794[(1'h1):(1'h1)] ?
                  ((-($signed(reg909) << {reg61,
                      (7'h49),
                      reg795})) || reg758[(3'h4):(1'h0)]) : reg782[(2'h2):(1'h0)]);
              reg923 = ($signed((reg869 ?
                      (wire3[(1'h1):(1'h0)] + {reg870}) : ($signed(reg653) ?
                          $unsigned((7'h54)) : {reg833, reg897, reg793}))) ?
                  (wire620[(4'h8):(4'h8)] == $unsigned(reg704[(1'h0):(1'h0)])) : reg631[(5'h11):(2'h3)]);
              reg924 = reg734;
              reg925 <= reg814[(1'h1):(1'h1)];
              reg926 <= wire7[(4'hf):(4'hb)];
              reg927 = ((-wire5) ? reg843[(3'h7):(3'h7)] : reg819);
            end
          else
            begin
              reg921 = ($signed(reg622[(3'h5):(2'h3)]) ?
                  ($signed(reg891) < reg906) : reg651);
              reg923 = $signed(reg659);
              reg924 = (reg830 ?
                  $signed((({(8'hbe), reg681, reg675} ?
                          $signed(reg903) : {reg762}) ?
                      (reg668[(5'h10):(3'h5)] ^~ {reg919,
                          reg889,
                          reg763}) : wire663)) : reg792[(3'h7):(2'h2)]);
              reg925 <= (7'h53);
              reg926 <= $signed(reg75);
              reg928 <= ($signed(reg64) ?
                  reg726 : $signed(reg895[(5'h17):(5'h11)]));
              reg929 <= reg914;
            end
          reg930 <= (($unsigned($signed(reg631[(5'h13):(3'h5)])) ?
                  (reg892 ?
                      reg914 : ((reg848 ?
                          reg74 : reg11) >>> (reg850 < (7'h54)))) : reg919[(2'h3):(1'h1)]) ?
              reg848[(2'h3):(1'h1)] : (~|(((!reg11) & wire5[(1'h0):(1'h0)]) ?
                  $signed((-reg761)) : (~$signed(reg43)))));
          for (forvar931 = (1'h0); (forvar931 < (2'h2)); forvar931 = (forvar931 + (1'h1)))
            begin
              reg932 = reg868[(3'h4):(2'h3)];
              reg933 <= reg622;
              reg934 <= reg917[(2'h2):(2'h2)];
              reg935 = reg832[(4'hb):(2'h3)];
              reg936 = reg803[(2'h3):(2'h3)];
              reg937 = ($unsigned($unsigned(((8'hac) ?
                      (wire854 ? reg728 : reg914) : (reg909 >>> reg654)))) ?
                  reg764 : ((|{reg68, $unsigned(reg10)}) ?
                      $signed(reg845) : (((reg625 ?
                          (8'ha2) : reg927) <<< $signed(reg784)) + $signed($unsigned((7'h56))))));
            end
          reg938 <= (|{reg41[(1'h1):(1'h0)], reg935[(4'hf):(3'h4)]});
          reg939 <= (reg937[(4'hb):(4'ha)] == (~&{$unsigned((reg647 - wire1))}));
          reg940 <= reg39[(4'ha):(4'h9)];
        end
      else
        begin
          reg922 <= reg899;
          reg923 = ($unsigned($unsigned(reg774[(2'h2):(1'h0)])) ?
              ((~$unsigned((!wire1))) ?
                  ((~&(reg655 > reg889)) > reg672) : (~reg640[(4'h8):(3'h4)])) : (&$unsigned((~&(reg733 ~^ reg674)))));
          if ((^~(7'h4d)))
            begin
              reg925 <= $unsigned(reg927[(3'h7):(2'h3)]);
              reg927 = ((reg647 ?
                  reg665[(4'h8):(3'h5)] : $unsigned($signed($unsigned(reg61)))) > (($signed($signed(reg700)) < (reg816 + ((8'hb8) == reg888))) == $unsigned(((reg686 != reg745) ?
                  $signed(reg660) : $unsigned((7'h4c))))));
              reg931 = reg659[(1'h0):(1'h0)];
            end
          else
            begin
              reg925 <= $unsigned((($unsigned((-(8'hb7))) != ((7'h53) ?
                  ((8'hb5) > reg847) : reg910[(1'h0):(1'h0)])) >>> ((~|{reg42,
                  (8'hbb)}) * (^(wire835 & reg898)))));
              reg927 = {$signed($unsigned(reg803[(1'h1):(1'h0)])),
                  {reg719[(2'h2):(1'h1)], reg843[(4'h8):(3'h6)]},
                  reg850};
              reg931 = $unsigned($signed($unsigned(reg71[(1'h1):(1'h0)])));
              reg932 = reg647;
              reg933 <= reg670;
              reg934 <= reg811;
              reg938 <= reg893[(4'h8):(3'h5)];
            end
          if ((-($signed((-reg653)) >> $signed({(reg870 | reg907),
              reg902,
              (^reg847)}))))
            begin
              reg941 = reg891[(2'h2):(1'h0)];
            end
          else
            begin
              reg941 = ($unsigned($signed($signed(((8'hb4) ?
                  reg933 : reg64)))) ~^ (reg738[(4'h9):(4'h8)] <<< (((~^(8'hb4)) ?
                  (reg774 ?
                      reg937 : reg46) : (reg672 <<< reg916)) && $unsigned(reg625[(2'h3):(2'h2)]))));
              reg942 <= $signed(($unsigned($signed(reg728[(2'h2):(1'h0)])) & (^~($unsigned(reg32) ?
                  ((8'hbf) ? reg845 : wire835) : (reg909 ? reg930 : reg71)))));
            end
          reg943 = (|reg766);
          if ((reg727 ? $unsigned(reg932) : reg925))
            begin
              reg944 <= $unsigned($signed(($unsigned($unsigned((8'had))) ?
                  (~|(reg41 ? reg814 : reg64)) : reg774)));
              reg945 = ((~^forvar896[(5'h14):(1'h0)]) ?
                  reg889 : (^~(|reg943[(1'h1):(1'h1)])));
              reg946 = {reg916[(5'h12):(1'h1)]};
              reg947 <= reg634[(2'h2):(1'h0)];
              reg948 = ({(-$signed((~reg694))),
                  $unsigned(({reg907, reg672, reg625} != ((7'h4d) ?
                      (8'hab) : (7'h44)))),
                  $signed(($signed(reg888) ?
                      reg916 : $signed(reg754)))} & reg832[(5'h10):(2'h2)]);
            end
          else
            begin
              reg944 <= $signed($unsigned(reg756));
              reg947 <= {$unsigned((reg845[(2'h2):(1'h1)] ?
                      $signed({reg685, wire835}) : (~&(^~reg631))))};
              reg948 = $signed({wire6,
                  (((7'h49) ? $unsigned(reg774) : (reg817 ? reg25 : (8'hbf))) ?
                      $signed((|reg727)) : reg754[(4'hd):(4'hd)]),
                  $signed(reg807)});
              reg949 = (8'hbb);
              reg950 = (|reg694);
              reg951 = {((&$unsigned((reg870 > reg672))) == $unsigned($signed((~reg19))))};
              reg952 = reg947[(1'h1):(1'h1)];
            end
        end
      for (forvar953 = (1'h0); (forvar953 < (2'h3)); forvar953 = (forvar953 + (1'h1)))
        begin
          reg954 <= $unsigned((!(($signed((8'haa)) ?
                  $unsigned(reg714) : reg908) ?
              ((reg869 ? wire2 : reg648) >>> (|reg938)) : reg886)));
          if ({(($unsigned(reg742) - {$signed(reg884),
                      reg64[(5'h18):(5'h14)],
                      reg717[(4'h8):(3'h6)]}) ?
                  $signed(((reg738 >>> reg737) >>> (reg814 >= (8'ha8)))) : (8'hae)),
              ($signed($unsigned(reg892[(3'h4):(2'h2)])) + (-$unsigned(wire6[(3'h6):(3'h5)]))),
              $unsigned($signed($unsigned(wire6)))})
            begin
              reg955 <= {forvar905[(4'hd):(4'hd)],
                  $signed({(~^(reg715 ~^ (7'h54))), $signed(reg946)}),
                  (~^({$signed(reg937), (-(7'h41)), reg945} ?
                      $signed((!reg885)) : (7'h45)))};
              reg956 <= wire855[(5'h19):(5'h14)];
              reg957 = ($signed((((|reg654) - $unsigned(reg761)) ?
                      wire663 : (8'hab))) ?
                  reg951[(5'h18):(2'h2)] : $signed(($signed((^~reg908)) ?
                      $unsigned((reg36 < reg908)) : reg659)));
              reg958 = $signed($signed(reg786));
              reg959 <= reg844;
              reg960 = reg667[(4'hc):(1'h0)];
              reg961 <= ($signed(($unsigned((7'h4e)) && ($unsigned((8'ha2)) ?
                      (reg811 ? reg774 : reg897) : (reg887 & forvar905)))) ?
                  reg75 : $signed(reg742));
            end
          else
            begin
              reg955 <= reg890;
              reg956 <= (($signed(((reg771 ^ reg39) <<< (&reg838))) >> $signed((reg662[(4'he):(3'h6)] & (reg751 ?
                  (8'hb5) : reg801)))) ^~ (^reg959[(4'h8):(3'h7)]));
              reg957 = reg625[(3'h4):(1'h0)];
              reg959 <= $signed($signed($signed(reg957[(4'he):(4'h9)])));
              reg961 <= $unsigned({$signed($unsigned(reg784[(5'h12):(5'h12)]))});
              reg962 <= (&reg944);
            end
        end
      reg963 = (~^reg814[(2'h3):(2'h2)]);
      reg964 <= reg915;
      if ($unsigned(($signed($signed((8'hb9))) < reg782)))
        begin
          if ($signed($unsigned((~^wire881))))
            begin
              reg965 <= $signed((!({{wire6},
                  {reg52, (8'ha4)}} >= $signed($unsigned(wire5)))));
              reg966 <= ((-{(|(reg640 ? reg815 : reg842)),
                      reg908[(3'h5):(1'h0)]}) ?
                  (reg71[(4'hb):(3'h5)] ?
                      $signed(reg792[(5'h15):(5'h13)]) : $unsigned(reg640[(4'hb):(3'h6)])) : $unsigned(reg962[(5'h18):(5'h18)]));
              reg967 <= (~(7'h46));
              reg968 <= $unsigned((($unsigned($unsigned(reg738)) + {((8'haf) ?
                      (8'hbc) : reg885),
                  $unsigned(reg909)}) < reg961[(2'h3):(1'h0)]));
              reg969 = reg672;
              reg970 <= reg795;
            end
          else
            begin
              reg969 = $signed({$signed($signed(reg771[(4'hb):(3'h6)])),
                  (-reg920[(4'hc):(2'h2)]),
                  ((~|reg670[(2'h2):(1'h1)]) ?
                      {reg640[(4'ha):(4'h9)],
                          (reg899 ? reg638 : reg21),
                          (reg61 == reg664)} : (~&(reg943 & reg900)))});
              reg970 <= reg909[(4'he):(3'h6)];
              reg971 = reg750[(2'h2):(2'h2)];
              reg972 = (&({$signed($signed(reg35)),
                      (!(reg846 ? reg717 : reg704))} ?
                  ((8'hab) ^ $unsigned((+reg782))) : (~^($signed(reg61) + $unsigned(reg21)))));
            end
          reg973 = (~&reg58[(2'h2):(1'h1)]);
          reg974 <= reg714;
        end
      else
        begin
          reg965 <= reg937[(4'ha):(3'h7)];
          reg966 <= (reg25 >> ($signed(((reg804 ? reg640 : reg950) ?
              $signed(reg872) : (^~reg948))) | ((wire880[(2'h2):(2'h2)] ^~ reg964[(4'hb):(4'h9)]) ^~ {(!(7'h52)),
              (reg936 ? reg39 : reg756)})));
          if ((((7'h58) ?
                  (reg714[(4'he):(4'h9)] ?
                      (^~$signed(reg682)) : {reg13,
                          $unsigned(reg762),
                          $unsigned(reg913)}) : (~^(~|reg742))) ?
              (^~(reg969[(5'h16):(3'h6)] ?
                  ((reg631 <= reg46) ?
                      (reg949 ~^ reg750) : ((8'hbe) ^ reg945)) : $unsigned((reg727 ?
                      reg956 : wire6)))) : reg924))
            begin
              reg967 <= (wire7[(4'hf):(1'h0)] ?
                  reg925 : ((&reg14) ?
                      $signed(reg933) : (reg954 ?
                          reg638[(5'h10):(3'h6)] : {$unsigned((8'hb8)),
                              (reg920 >>> reg964)})));
              reg969 = (~^$unsigned(reg933));
            end
          else
            begin
              reg969 = reg869[(2'h2):(1'h0)];
              reg971 = (reg884[(3'h6):(3'h6)] ?
                  $signed({(reg963[(5'h13):(4'hb)] == (reg842 >> wire2)),
                      $unsigned($signed(reg942))}) : $signed((((reg801 ?
                          reg930 : reg913) ?
                      ((7'h4f) ? (7'h4b) : reg885) : {reg960,
                          wire5}) || $unsigned((reg36 ? reg665 : reg920)))));
              reg974 <= reg784[(4'hb):(3'h4)];
              reg975 <= {{$signed(forvar896[(1'h1):(1'h1)])}, reg842};
              reg976 = (~|$signed($signed({{reg19, reg898},
                  {reg13, reg42, wire6},
                  (reg19 ? reg68 : reg908)})));
              reg977 <= $unsigned(($unsigned($signed((&reg895))) * (({(8'ha5),
                      reg907} ?
                  (reg908 > reg932) : {reg951, reg960}) | ($unsigned(reg893) ?
                  (reg930 < wire663) : (reg975 ? reg901 : reg788)))));
              reg978 <= reg786[(4'hf):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      if ((reg58 <= (reg670[(5'h10):(4'hf)] ?
          $unsigned(({reg682} ?
              (8'hb7) : (reg761 >>> reg634))) : $unsigned($signed((&reg940))))))
        begin
          if ((7'h56))
            begin
              reg979 <= reg52;
            end
          else
            begin
              reg980 = $unsigned(reg870);
              reg981 = (7'h46);
              reg982 <= (7'h55);
              reg983 = ($signed((((-reg888) ^~ reg677[(5'h11):(4'hc)]) < {wire663,
                  $unsigned(reg655)})) * reg700[(4'he):(4'he)]);
              reg984 = (|(($signed($signed((7'h4f))) ^~ reg783[(1'h1):(1'h0)]) ?
                  ($signed((~|reg795)) ?
                      $signed((reg870 < reg979)) : $signed(((7'h4b) != (8'ha5)))) : wire1[(3'h6):(3'h6)]));
              reg985 = $unsigned(reg900[(1'h1):(1'h1)]);
              reg986 <= reg910;
            end
          for (forvar987 = (1'h0); (forvar987 < (3'h6)); forvar987 = (forvar987 + (1'h1)))
            begin
              reg988 <= ($signed(($signed($unsigned((8'hae))) <= reg42)) >>> (-reg968));
              reg989 <= reg759;
            end
          for (forvar990 = (1'h0); (forvar990 < (2'h3)); forvar990 = (forvar990 + (1'h1)))
            begin
              reg991 = {$signed($unsigned(reg753)), (^~$unsigned(reg920))};
              reg992 <= $unsigned($unsigned($signed(reg668)));
              reg993 <= (wire879[(2'h2):(1'h0)] ?
                  (($unsigned(reg766) ?
                      $signed({reg966,
                          reg830}) : ((reg928 * reg684) <<< (!reg848))) >>> (7'h4f)) : $signed($signed(reg61[(5'h17):(4'hc)])));
              reg994 <= (~^(~|$signed($signed((~|(7'h4d))))));
            end
          if ((reg13[(2'h3):(1'h0)] ~^ wire2))
            begin
              reg995 = reg970;
            end
          else
            begin
              reg995 = (&(&(reg783 ? reg977 : reg784)));
              reg996 = (reg974[(5'h1a):(4'hc)] ?
                  (!($unsigned($unsigned(reg979)) ?
                      (reg831[(5'h17):(3'h6)] ?
                          (~^(7'h49)) : (wire3 ?
                              reg933 : reg989)) : reg922)) : $unsigned((^$unsigned((reg11 && reg14)))));
              reg997 = {((reg683[(4'h9):(3'h7)] ?
                      $unsigned((8'hb4)) : (^(reg14 ?
                          reg970 : reg980))) == (&(~^(~&reg728)))),
                  (-reg683),
                  $unsigned((((-reg751) ?
                      (reg859 ? (7'h43) : reg685) : reg988) || reg900))};
              reg998 <= (((^~(+$unsigned(reg887))) ?
                      $unsigned(reg974[(5'h14):(4'he)]) : reg679[(2'h2):(2'h2)]) ?
                  $signed(reg908) : (&(~|(reg929 * (~&reg14)))));
            end
          reg999 <= ({reg634[(1'h0):(1'h0)],
                  $unsigned($signed($unsigned(reg653)))} ?
              forvar990[(4'h9):(3'h7)] : $unsigned(((!reg984) >> (+(reg954 > reg833)))));
          if (({reg956[(4'he):(4'hc)]} <<< (8'ha4)))
            begin
              reg1000 <= $signed(reg970);
              reg1001 <= reg737;
              reg1002 = $signed($signed(({reg32,
                  reg625[(4'h8):(3'h6)]} | $signed((reg967 ?
                  reg956 : reg653)))));
              reg1003 <= {$signed((((+reg19) ?
                          (~reg966) : (reg895 ? (8'hb6) : reg10)) ?
                      (reg681[(3'h4):(3'h4)] ?
                          {reg660} : $unsigned(reg68)) : $signed(reg908[(2'h2):(2'h2)]))),
                  (!$unsigned($signed(reg968))),
                  (reg700[(1'h1):(1'h0)] != ({{reg638, reg43},
                      $unsigned(reg888)} == $unsigned(reg625)))};
              reg1004 <= $signed($signed($unsigned($signed(reg774[(1'h0):(1'h0)]))));
              reg1005 = $unsigned(((((~^reg14) - reg1003[(2'h3):(1'h1)]) < ($unsigned(reg993) ?
                      reg68 : $signed(forvar987))) ?
                  $unsigned((^$unsigned((8'ha9)))) : (+({reg850,
                          reg845,
                          reg814} ?
                      wire854 : reg25))));
            end
          else
            begin
              reg1002 = (reg774[(2'h2):(1'h0)] ?
                  wire5 : ($signed(reg719[(2'h2):(2'h2)]) ?
                      reg34 : reg678[(4'hc):(1'h1)]));
            end
        end
      else
        begin
          for (forvar979 = (1'h0); (forvar979 < (2'h2)); forvar979 = (forvar979 + (1'h1)))
            begin
              reg982 <= reg678[(5'h11):(3'h6)];
              reg986 <= reg783;
            end
          if ({reg657[(4'ha):(3'h5)], (!reg764[(4'h8):(3'h5)]), reg778})
            begin
              reg987 <= (~&(|reg981));
              reg990 = {((($signed(reg982) <= (reg977 + wire881)) ?
                      forvar990[(4'hc):(2'h2)] : ($signed(wire7) != ((8'ha8) ?
                          reg647 : reg850))) ~^ $unsigned(reg52[(5'h14):(4'hc)])),
                  {reg43, (^$signed(reg819))},
                  reg788};
              reg991 = $unsigned({reg684,
                  (^$signed($signed(forvar987))),
                  {$signed($unsigned((7'h54))), $unsigned($unsigned(reg737))}});
              reg992 <= reg63;
            end
          else
            begin
              reg987 <= ($signed((reg759 ?
                      ($unsigned(reg681) ?
                          (7'h4b) : reg657[(5'h15):(5'h12)]) : ($signed(reg784) ?
                          {(7'h4f)} : {(7'h49)}))) ?
                  reg764 : (^$signed($signed($unsigned(reg759)))));
            end
          for (forvar993 = (1'h0); (forvar993 < (3'h6)); forvar993 = (forvar993 + (1'h1)))
            begin
              reg995 = (8'ha8);
              reg998 <= ($signed((((reg966 <<< reg870) ?
                          (8'hb4) : (reg979 ? reg68 : reg981)) ?
                      wire852[(1'h0):(1'h0)] : (!$unsigned(reg917)))) ?
                  (!(&(|reg901))) : {reg920[(4'hf):(4'he)],
                      $signed((+reg781))});
              reg1002 = reg955[(4'hd):(3'h7)];
              reg1003 <= $unsigned($unsigned($unsigned((+$unsigned(reg681)))));
            end
          reg1005 = ($unsigned(reg974[(4'hc):(4'h9)]) <= $unsigned((reg47 ?
              reg761[(2'h3):(1'h1)] : ((^~reg916) ?
                  reg714[(4'hd):(3'h5)] : $unsigned(reg985)))));
          for (forvar1006 = (1'h0); (forvar1006 < (1'h1)); forvar1006 = (forvar1006 + (1'h1)))
            begin
              reg1007 <= wire663[(4'h9):(3'h4)];
              reg1008 <= wire854;
              reg1009 <= reg700;
              reg1010 = ((8'ha7) > ($unsigned(reg1008) && reg869));
              reg1011 = {(($signed((reg980 < reg966)) && reg778) ?
                      $unsigned($unsigned($unsigned(reg43))) : (^~reg783[(1'h1):(1'h0)]))};
            end
          if (reg648)
            begin
              reg1012 = reg968[(4'hd):(4'ha)];
              reg1013 <= ($signed(reg717) << $unsigned($unsigned((^{reg942}))));
              reg1014 = ($signed(reg679) ?
                  $signed(((~$signed(reg21)) ?
                      ((wire835 ? reg758 : reg19) > {reg36}) : {{reg975,
                              reg885},
                          reg52})) : {$signed($unsigned((forvar993 ?
                          reg928 : (7'h47))))});
              reg1015 = (reg992 < $signed(reg966[(3'h6):(3'h4)]));
              reg1016 = reg816[(3'h5):(2'h3)];
            end
          else
            begin
              reg1013 <= $unsigned(reg801[(2'h2):(1'h0)]);
              reg1014 = (reg1013[(5'h10):(1'h0)] ?
                  {reg58[(2'h2):(2'h2)],
                      reg1003[(2'h3):(2'h2)]} : ($signed(reg68) | (^~reg959)));
              reg1015 = reg962;
            end
          for (forvar1017 = (1'h0); (forvar1017 < (3'h4)); forvar1017 = (forvar1017 + (1'h1)))
            begin
              reg1018 = reg11;
              reg1019 = $signed(wire879[(4'hc):(2'h2)]);
              reg1020 <= ((reg964 ?
                      reg1005[(4'h9):(2'h3)] : $signed((!{reg961,
                          reg778,
                          reg665}))) ?
                  $signed(reg998[(3'h4):(1'h0)]) : reg637[(3'h6):(2'h3)]);
              reg1021 = ((($unsigned((reg981 == (7'h49))) >= ($signed(reg925) - (reg742 << reg677))) ?
                  reg642 : $unsigned({reg622[(4'h8):(1'h0)],
                      (reg782 ? reg883 : (8'h9c))})) + {reg19});
              reg1022 = (+((reg638 ?
                      $unsigned((reg942 ? reg726 : reg19)) : ((reg49 ?
                          (7'h43) : reg814) >= $signed(reg928))) ?
                  ({$unsigned(reg764), $signed(reg777), {reg13}} >= {reg868,
                      $unsigned((8'h9e))}) : ($unsigned((reg894 + reg1016)) * reg49[(2'h3):(1'h0)])));
            end
        end
      if ((reg962 >> reg660[(4'he):(3'h5)]))
        begin
          if ((reg926 ?
              $unsigned((($unsigned(reg41) == reg678[(5'h11):(4'hb)]) ?
                  reg701 : ((reg743 < reg983) ?
                      (wire854 > reg801) : (reg940 ?
                          (8'hbe) : reg1014)))) : $unsigned((($signed(reg763) >= $signed(reg653)) | reg742))))
            begin
              reg1023 = ((-$unsigned((~(~wire2)))) ?
                  $unsigned($signed(reg970[(4'ha):(3'h5)])) : $signed((($unsigned((7'h56)) ?
                          ((8'hb4) ? (8'hae) : reg667) : $unsigned(reg1011)) ?
                      ({reg838, reg920, reg35} ?
                          reg962 : $signed(reg726)) : (&(reg975 ?
                          wire0 : reg672)))));
              reg1024 = reg629[(5'h18):(4'h9)];
              reg1025 = (|reg1007);
              reg1026 = reg783;
              reg1027 = ($unsigned($unsigned({reg727})) + $signed((|reg47[(3'h7):(2'h2)])));
              reg1028 <= reg708;
              reg1029 = reg734[(4'hb):(3'h6)];
            end
          else
            begin
              reg1023 = $unsigned($unsigned(($unsigned((reg52 == reg961)) ?
                  $signed((reg715 ? wire620 : reg1018)) : reg859)));
              reg1028 <= $unsigned(reg983[(3'h5):(1'h1)]);
              reg1030 <= $signed(reg922);
              reg1031 <= $unsigned($signed($signed(reg27)));
              reg1032 <= (reg942[(3'h4):(1'h1)] == $signed($signed(reg1018)));
            end
          reg1033 <= $unsigned((!(~&reg933[(2'h3):(1'h1)])));
          reg1034 = (reg1013[(4'ha):(2'h3)] ? reg1021 : reg678);
          reg1035 <= $unsigned(reg1018[(4'ha):(3'h5)]);
          if (((-reg939[(5'h11):(4'hc)]) ?
              $unsigned(((|(reg708 * reg938)) || (((7'h46) ?
                  reg638 : wire5) | (!reg712)))) : reg804))
            begin
              reg1036 <= ({(((reg1018 ? wire0 : forvar1006) ?
                      reg764[(3'h7):(2'h2)] : $unsigned(reg694)) ^ ($signed(wire4) || (7'h4e))),
                  $unsigned(((reg819 ? reg980 : reg733) ?
                      $signed(reg763) : (reg922 ? reg967 : reg43))),
                  (({reg1002} ?
                      (reg647 ?
                          reg888 : reg1002) : (reg916 ~^ reg52)) >>> reg885[(1'h0):(1'h0)])} ~^ (reg984[(4'h8):(3'h5)] ^~ $unsigned({reg1007})));
              reg1037 <= reg638;
              reg1038 <= reg19[(4'hc):(4'hb)];
              reg1039 <= (~^((7'h45) != $signed((+(~&reg1034)))));
              reg1040 = (~|reg679);
              reg1041 <= ((&reg777) != $signed(wire663[(2'h3):(2'h2)]));
              reg1042 = (^~(~|$signed((8'ha4))));
            end
          else
            begin
              reg1040 = (((~&($signed(reg788) ?
                      $unsigned(reg928) : $signed((8'hb7)))) - $signed((+(reg966 ?
                      (8'hb3) : (8'ha2))))) ?
                  (reg901 == $signed((reg74 ?
                      $unsigned(reg1028) : (!reg1016)))) : $unsigned((^reg74[(3'h4):(1'h1)])));
              reg1041 <= $unsigned(reg838);
              reg1042 = reg626;
              reg1043 = ((-($signed(reg992[(4'hc):(1'h0)]) ?
                  {(!reg13)} : (~|$unsigned((8'hb1))))) + ($signed(((|reg640) ^ reg1033)) & (^~reg738[(3'h7):(3'h4)])));
              reg1044 = {$unsigned(reg1023)};
              reg1045 <= ($unsigned($unsigned($signed($unsigned(reg1026)))) || (^$signed(((reg784 ~^ reg751) ?
                  ((7'h43) ? reg1001 : reg751) : (reg847 && (8'h9d))))));
              reg1046 = reg751[(1'h1):(1'h1)];
            end
          reg1047 = reg994;
          if ((^({reg847[(4'he):(3'h5)],
              reg783[(4'h8):(4'h8)]} && (!$unsigned({reg1030, (8'ha3)})))))
            begin
              reg1048 = $unsigned($signed((-reg869[(4'he):(4'h8)])));
              reg1049 <= $signed({(reg679 + $signed(reg712))});
              reg1050 <= (&(^~$unsigned($signed(reg784[(5'h15):(4'ha)]))));
              reg1051 <= $signed($unsigned(reg929[(5'h11):(5'h10)]));
              reg1052 = {$unsigned($signed(reg901[(2'h2):(2'h2)])),
                  reg996[(3'h5):(3'h5)],
                  {(~^($unsigned(reg653) ? {wire1} : reg700))}};
            end
          else
            begin
              reg1048 = reg832[(4'hb):(3'h5)];
              reg1049 <= reg900;
              reg1050 <= ($unsigned(reg1033[(1'h0):(1'h0)]) <= reg697[(2'h3):(2'h2)]);
              reg1051 <= (((7'h4d) > $signed($signed($unsigned((8'hb2))))) ?
                  ((reg966 ?
                      reg845[(1'h0):(1'h0)] : reg801[(4'ha):(4'h9)]) >>> (~|{(^(8'hbe))})) : (((wire5 ?
                          (reg781 ? reg1000 : reg793) : $signed(reg660)) ?
                      (reg1047[(2'h2):(2'h2)] ?
                          $signed(wire881) : (~reg817)) : $signed((reg979 <= reg625))) > $signed(reg1025[(4'he):(4'ha)])));
              reg1052 = {$unsigned(reg675[(4'h8):(4'h8)])};
              reg1053 <= ({$signed(((^~reg1045) ?
                      $signed(reg742) : ((7'h40) == reg979)))} >= ($signed({reg956,
                      $signed(reg925),
                      {reg978, reg955, reg1028}}) ?
                  $signed(($signed(reg727) * $signed(reg984))) : reg929[(4'h9):(2'h3)]));
              reg1054 <= $signed({((7'h4a) ~^ ((reg988 >> (8'ha5)) ?
                      reg664 : (reg653 * reg964))),
                  $unsigned(($signed(reg1044) ?
                      reg1021[(4'h9):(2'h3)] : reg682[(3'h6):(3'h5)]))});
            end
        end
      else
        begin
          reg1023 = (~&$signed(reg39[(3'h7):(3'h5)]));
        end
      if ($unsigned(((({reg901} ? $unsigned(reg843) : (reg1003 && reg634)) ?
          (~reg801[(4'hc):(3'h6)]) : {$unsigned(reg928),
              wire881}) * forvar990[(1'h1):(1'h0)])))
        begin
          for (forvar1055 = (1'h0); (forvar1055 < (2'h3)); forvar1055 = (forvar1055 + (1'h1)))
            begin
              reg1056 = {(~(wire855 ?
                      ($unsigned(forvar990) && reg25[(4'h8):(1'h0)]) : (reg917[(2'h2):(1'h1)] | reg756)))};
              reg1057 <= (~(^reg701));
              reg1058 = ($unsigned({($signed((8'hb2)) ?
                      (reg1050 ?
                          forvar987 : reg733) : $unsigned(reg738))}) <= reg640[(3'h4):(2'h2)]);
              reg1059 = (7'h47);
            end
          reg1060 = reg728;
          for (forvar1061 = (1'h0); (forvar1061 < (1'h0)); forvar1061 = (forvar1061 + (1'h1)))
            begin
              reg1062 = $signed(reg1015[(5'h10):(3'h5)]);
              reg1063 = $unsigned(($unsigned((7'h57)) < ((reg1044 ?
                  (reg847 ~^ reg788) : $unsigned(reg727)) || ($signed(reg665) ?
                  $signed((7'h58)) : {reg998, reg1048}))));
              reg1064 = (-($signed((7'h4f)) > (-($unsigned(reg965) ?
                  (|reg683) : (^~reg58)))));
              reg1065 = $signed({((^~(reg994 - reg831)) <= $unsigned(reg801[(3'h4):(3'h4)]))});
              reg1066 = $signed((&((reg843[(3'h6):(2'h2)] ?
                  {reg929} : {reg49,
                      reg940,
                      reg691}) && $signed(reg714[(3'h6):(3'h4)]))));
              reg1067 <= (^$signed(((~&(reg885 ? reg999 : forvar1061)) ?
                  reg979 : wire7)));
              reg1068 <= $unsigned((+(((reg846 >= reg640) ?
                      $unsigned((7'h42)) : reg39) ?
                  ((^forvar1061) ?
                      (reg682 ?
                          reg648 : reg795) : (reg819 ^~ wire7)) : $unsigned($signed(reg654)))));
            end
        end
      else
        begin
          reg1055 = reg19[(3'h7):(3'h5)];
          for (forvar1056 = (1'h0); (forvar1056 < (2'h2)); forvar1056 = (forvar1056 + (1'h1)))
            begin
              reg1058 = ((reg1000 ?
                      (^wire1[(3'h6):(3'h4)]) : (+reg1021[(5'h14):(4'hb)])) ?
                  (reg634[(1'h0):(1'h0)] ?
                      ($unsigned((reg764 >>> reg845)) || reg888) : reg781) : ($signed(reg667) && $signed($unsigned(wire835[(4'hb):(2'h2)]))));
              reg1059 = reg651;
            end
          if ((^(8'hbd)))
            begin
              reg1061 <= reg832;
              reg1062 = wire6[(3'h5):(1'h1)];
            end
          else
            begin
              reg1061 <= (~&(~^reg847));
              reg1062 = ($unsigned(reg930) < {$unsigned(reg956[(5'h15):(4'he)])});
              reg1063 = (-$unsigned((!$unsigned((&(7'h4c))))));
              reg1064 = $signed($signed($unsigned(((reg1036 ?
                  reg1066 : reg1022) << reg908[(3'h7):(2'h3)]))));
            end
          reg1065 = $unsigned($unsigned((reg759 ?
              (~|{reg675, reg871, reg1068}) : (reg64 ?
                  {reg794, reg942, reg686} : reg1057[(1'h0):(1'h0)]))));
          reg1066 = $unsigned(reg670);
          reg1069 = $unsigned((|(7'h4d)));
        end
      for (forvar1070 = (1'h0); (forvar1070 < (2'h2)); forvar1070 = (forvar1070 + (1'h1)))
        begin
          for (forvar1071 = (1'h0); (forvar1071 < (3'h6)); forvar1071 = (forvar1071 + (1'h1)))
            begin
              reg1072 <= ($unsigned({reg811[(5'h18):(5'h16)]}) ^ reg888[(4'h8):(2'h2)]);
            end
          if (($unsigned({(~&$unsigned((8'hbc))),
              ($signed(reg981) ? $signed(reg654) : (reg16 ? reg845 : reg908)),
              (+$unsigned(reg1050))}) <<< {{reg984[(4'ha):(3'h6)],
                  {$unsigned(reg784)},
                  $unsigned(((8'hab) ? (8'ha2) : reg883))}}))
            begin
              reg1073 = $signed(reg626[(4'h9):(2'h3)]);
            end
          else
            begin
              reg1074 <= {$signed((reg1014[(2'h3):(1'h0)] ?
                      {((8'hbe) ? reg657 : (8'ha9)),
                          $signed((8'hb5))} : $signed((reg909 >= reg831)))),
                  reg39[(4'ha):(4'h8)]};
              reg1075 <= forvar1017[(4'he):(3'h5)];
              reg1076 <= $signed(reg983);
              reg1077 = $unsigned($unsigned((7'h46)));
              reg1078 <= (($signed(reg1002) ?
                  (~^(|(^~(8'ha3)))) : {reg883,
                      (^(reg655 >> reg47))}) | reg660[(4'ha):(3'h7)]);
            end
        end
      if ($unsigned(($signed(reg771[(4'hb):(3'h4)]) | $signed($unsigned($signed(reg938))))))
        begin
          if (wire2)
            begin
              reg1079 = (reg642[(4'h9):(3'h5)] && ($unsigned((&{(8'hba),
                      reg804})) ?
                  reg42[(1'h0):(1'h0)] : $unsigned((~^reg901[(2'h3):(1'h0)]))));
              reg1080 <= reg1068[(2'h3):(1'h1)];
              reg1081 <= (&$signed({reg1008[(4'ha):(3'h5)]}));
            end
          else
            begin
              reg1080 <= (~&($signed($unsigned(reg1057[(1'h1):(1'h1)])) ?
                  (7'h44) : ((^$unsigned(reg1059)) > (~^$signed(reg648)))));
              reg1081 <= $unsigned((reg728[(1'h0):(1'h0)] <<< reg980));
              reg1082 <= $unsigned(((((^reg1074) ?
                      reg1069[(1'h1):(1'h0)] : forvar1061) ?
                  (8'hab) : (+(!reg926))) == $unsigned(($unsigned(reg63) > {reg1055,
                  (8'haf),
                  reg934}))));
            end
        end
      else
        begin
          if ((!forvar993))
            begin
              reg1079 = ($signed((($signed(reg966) ?
                      $unsigned(reg1051) : reg926) ?
                  $unsigned(((7'h49) ?
                      reg869 : reg938)) : reg954[(3'h7):(3'h4)])) - $signed((((^reg1079) & wire2[(1'h1):(1'h1)]) ?
                  $unsigned((reg1007 ?
                      reg1075 : (8'hbd))) : (^reg928[(4'h8):(3'h4)]))));
            end
          else
            begin
              reg1079 = (~&reg975[(4'h8):(3'h6)]);
              reg1080 <= $unsigned($unsigned($signed((((7'h4d) >= reg901) ?
                  reg991 : reg1062[(3'h5):(1'h1)]))));
              reg1083 = (((+reg909[(2'h3):(2'h2)]) ?
                  reg792 : forvar1017[(1'h1):(1'h0)]) ^~ $signed((reg1073 ?
                  (|reg887) : reg43)));
              reg1084 <= (((7'h46) <= (+$unsigned(reg910))) ?
                  reg1001[(1'h1):(1'h1)] : (~&reg831[(2'h2):(2'h2)]));
            end
        end
    end
  assign wire1085 = reg648[(4'he):(1'h1)];
  always
    @(posedge clk) begin
      reg1086 <= {(|{(~&(reg970 >= (8'hab)))}),
          (({(reg63 >= reg844), (-reg1001), ((8'ha7) != reg639)} ?
              reg1076[(2'h3):(1'h1)] : ((reg637 ?
                  reg734 : reg964) >> $unsigned(reg75))) < (&$unsigned(reg947)))};
      reg1087 <= $unsigned(((+$unsigned(reg1028[(1'h1):(1'h1)])) && $signed((reg1080[(4'hc):(1'h0)] ?
          {reg631, reg940} : (reg684 ? reg967 : wire855)))));
      reg1088 <= (^~(!$signed($unsigned((+reg846)))));
    end
  assign wire1089 = $unsigned({reg734[(2'h3):(2'h3)], (reg34 ~^ reg1074)});
  assign wire1090 = ($unsigned(reg761[(5'h14):(2'h3)]) < $unsigned(((reg654 == reg784) ?
                        $unsigned((reg762 ? reg811 : reg803)) : (8'hab))));
  assign wire1091 = $unsigned(reg975[(1'h1):(1'h1)]);
  assign wire1092 = ((7'h42) ?
                        $unsigned((!$unsigned({reg762,
                            reg764}))) : $signed($signed(((+reg25) + {reg887,
                            (8'haf)}))));
  assign wire1093 = $unsigned(reg734);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module77
#(parameter param618 = {{(~^(((7'h41) ? (8'hb3) : (8'hab)) * (~&(8'ha7)))), (^~((~&(8'hba)) ? ((8'h9f) ^ (8'had)) : (-(7'h52))))}}, 
parameter param619 = ((param618 ? param618 : (param618 ? (+{param618, param618}) : (param618 ? (param618 ? (8'h9f) : param618) : {param618}))) ? {{param618, (+{param618, param618, param618})}} : {{param618, (((7'h55) ? param618 : param618) - (^~param618))}, ((&(param618 == param618)) == {(param618 <= param618), param618, param618})}))
(y, clk, wire82, wire81, wire80, wire79, wire78);
  output wire [(32'h23d6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire82;
  input wire [(5'h14):(1'h0)] wire81;
  input wire signed [(5'h1c):(1'h0)] wire80;
  input wire [(4'h9):(1'h0)] wire79;
  input wire [(4'hc):(1'h0)] wire78;
  wire [(5'h12):(1'h0)] wire617;
  wire signed [(2'h2):(1'h0)] wire525;
  wire signed [(4'hc):(1'h0)] wire511;
  wire signed [(4'ha):(1'h0)] wire471;
  wire signed [(5'h1f):(1'h0)] wire470;
  wire [(4'he):(1'h0)] wire469;
  wire [(4'h8):(1'h0)] wire468;
  wire [(3'h7):(1'h0)] wire467;
  wire [(3'h7):(1'h0)] wire344;
  wire signed [(5'h12):(1'h0)] wire266;
  wire [(4'ha):(1'h0)] wire265;
  wire signed [(5'h12):(1'h0)] wire233;
  wire signed [(5'h15):(1'h0)] wire121;
  wire signed [(5'h13):(1'h0)] wire83;
  reg [(5'h17):(1'h0)] reg616 = (1'h0);
  reg [(5'h1e):(1'h0)] reg614 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg609 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg607 = (1'h0);
  reg [(2'h3):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg596 = (1'h0);
  reg [(4'he):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg594 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg590 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg588 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg585 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg583 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg581 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg580 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg577 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg567 = (1'h0);
  reg [(4'hf):(1'h0)] reg566 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg565 = (1'h0);
  reg [(5'h1c):(1'h0)] reg562 = (1'h0);
  reg [(2'h2):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg557 = (1'h0);
  reg [(4'hc):(1'h0)] reg556 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg555 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg553 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg552 = (1'h0);
  reg [(2'h2):(1'h0)] reg549 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg547 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg546 = (1'h0);
  reg [(5'h11):(1'h0)] reg545 = (1'h0);
  reg [(2'h3):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg538 = (1'h0);
  reg [(5'h18):(1'h0)] reg537 = (1'h0);
  reg signed [(4'he):(1'h0)] reg536 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg535 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg533 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg528 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg521 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg517 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg516 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg513 = (1'h0);
  reg [(5'h1d):(1'h0)] reg510 = (1'h0);
  reg [(5'h1a):(1'h0)] reg506 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg505 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg502 = (1'h0);
  reg [(4'hc):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg496 = (1'h0);
  reg [(4'ha):(1'h0)] reg494 = (1'h0);
  reg [(4'he):(1'h0)] reg493 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg486 = (1'h0);
  reg [(4'h9):(1'h0)] reg483 = (1'h0);
  reg [(5'h10):(1'h0)] reg481 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg477 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg476 = (1'h0);
  reg [(5'h12):(1'h0)] reg473 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg466 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg465 = (1'h0);
  reg [(3'h4):(1'h0)] reg464 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg463 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg462 = (1'h0);
  reg [(5'h1b):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg453 = (1'h0);
  reg [(5'h19):(1'h0)] reg451 = (1'h0);
  reg [(5'h19):(1'h0)] reg449 = (1'h0);
  reg [(5'h11):(1'h0)] reg448 = (1'h0);
  reg [(4'hd):(1'h0)] reg446 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg443 = (1'h0);
  reg [(4'hf):(1'h0)] reg441 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg440 = (1'h0);
  reg [(5'h1f):(1'h0)] reg437 = (1'h0);
  reg [(2'h2):(1'h0)] reg438 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg435 = (1'h0);
  reg [(5'h1a):(1'h0)] reg434 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg431 = (1'h0);
  reg [(4'hc):(1'h0)] reg427 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg426 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg424 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg422 = (1'h0);
  reg [(5'h1c):(1'h0)] reg421 = (1'h0);
  reg [(4'hf):(1'h0)] reg419 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg412 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg410 = (1'h0);
  reg [(5'h11):(1'h0)] reg409 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg402 = (1'h0);
  reg [(2'h3):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg398 = (1'h0);
  reg [(5'h12):(1'h0)] reg396 = (1'h0);
  reg signed [(4'he):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg394 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg393 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg392 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg387 = (1'h0);
  reg [(3'h7):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg382 = (1'h0);
  reg [(4'h8):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg380 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg376 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg371 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg369 = (1'h0);
  reg [(4'h9):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg363 = (1'h0);
  reg [(5'h14):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg361 = (1'h0);
  reg [(4'h8):(1'h0)] reg359 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg355 = (1'h0);
  reg [(4'h9):(1'h0)] reg354 = (1'h0);
  reg [(5'h1d):(1'h0)] reg353 = (1'h0);
  reg [(5'h11):(1'h0)] reg352 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg347 = (1'h0);
  reg [(5'h10):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg343 = (1'h0);
  reg [(5'h1f):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg339 = (1'h0);
  reg [(4'he):(1'h0)] reg336 = (1'h0);
  reg [(4'hc):(1'h0)] reg332 = (1'h0);
  reg signed [(4'he):(1'h0)] reg330 = (1'h0);
  reg [(5'h1e):(1'h0)] reg329 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg324 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg322 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg321 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg320 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg318 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg313 = (1'h0);
  reg [(5'h1e):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg309 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg307 = (1'h0);
  reg [(4'he):(1'h0)] reg298 = (1'h0);
  reg [(5'h12):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg293 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg289 = (1'h0);
  reg signed [(4'he):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg286 = (1'h0);
  reg [(5'h1d):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg284 = (1'h0);
  reg [(5'h17):(1'h0)] reg281 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg280 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg279 = (1'h0);
  reg [(4'h8):(1'h0)] reg277 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg274 = (1'h0);
  reg [(3'h5):(1'h0)] reg270 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg262 = (1'h0);
  reg [(4'ha):(1'h0)] reg260 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg258 = (1'h0);
  reg [(5'h17):(1'h0)] reg255 = (1'h0);
  reg [(5'h10):(1'h0)] reg254 = (1'h0);
  reg [(4'hb):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg251 = (1'h0);
  reg [(4'ha):(1'h0)] reg250 = (1'h0);
  reg [(5'h1a):(1'h0)] reg249 = (1'h0);
  reg [(4'he):(1'h0)] reg246 = (1'h0);
  reg [(5'h1d):(1'h0)] reg241 = (1'h0);
  reg [(5'h12):(1'h0)] reg239 = (1'h0);
  reg [(5'h1a):(1'h0)] reg236 = (1'h0);
  reg [(5'h11):(1'h0)] reg232 = (1'h0);
  reg [(5'h1a):(1'h0)] reg229 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg227 = (1'h0);
  reg [(5'h15):(1'h0)] reg226 = (1'h0);
  reg [(4'hf):(1'h0)] reg224 = (1'h0);
  reg [(5'h19):(1'h0)] reg219 = (1'h0);
  reg [(5'h12):(1'h0)] reg218 = (1'h0);
  reg [(2'h3):(1'h0)] reg216 = (1'h0);
  reg [(5'h14):(1'h0)] reg215 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg213 = (1'h0);
  reg [(2'h2):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg211 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg210 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg208 = (1'h0);
  reg [(5'h12):(1'h0)] reg206 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg205 = (1'h0);
  reg [(4'h9):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg202 = (1'h0);
  reg [(5'h18):(1'h0)] reg192 = (1'h0);
  reg [(5'h1f):(1'h0)] reg191 = (1'h0);
  reg [(5'h15):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg187 = (1'h0);
  reg [(5'h13):(1'h0)] reg186 = (1'h0);
  reg [(5'h11):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg178 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg175 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg174 = (1'h0);
  reg [(3'h5):(1'h0)] reg167 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg164 = (1'h0);
  reg [(5'h11):(1'h0)] reg162 = (1'h0);
  reg [(3'h4):(1'h0)] reg157 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg156 = (1'h0);
  reg [(5'h1d):(1'h0)] reg154 = (1'h0);
  reg [(5'h11):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg150 = (1'h0);
  reg [(5'h1f):(1'h0)] reg149 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg146 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg143 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg142 = (1'h0);
  reg [(5'h14):(1'h0)] reg139 = (1'h0);
  reg [(5'h10):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg125 = (1'h0);
  reg [(2'h3):(1'h0)] reg124 = (1'h0);
  reg [(5'h1c):(1'h0)] reg122 = (1'h0);
  reg [(5'h1d):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg119 = (1'h0);
  reg [(4'ha):(1'h0)] reg115 = (1'h0);
  reg [(5'h14):(1'h0)] reg114 = (1'h0);
  reg [(5'h1b):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg101 = (1'h0);
  reg [(4'he):(1'h0)] reg99 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg97 = (1'h0);
  reg [(5'h10):(1'h0)] reg96 = (1'h0);
  reg [(3'h6):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg92 = (1'h0);
  reg [(4'h8):(1'h0)] reg88 = (1'h0);
  reg [(4'hc):(1'h0)] reg87 = (1'h0);
  reg [(4'h8):(1'h0)] reg85 = (1'h0);
  reg [(5'h17):(1'h0)] reg84 = (1'h0);
  reg [(5'h1b):(1'h0)] reg615 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg613 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar612 = (1'h0);
  reg [(5'h17):(1'h0)] forvar611 = (1'h0);
  reg [(4'hc):(1'h0)] reg610 = (1'h0);
  reg [(4'hd):(1'h0)] reg606 = (1'h0);
  reg [(2'h3):(1'h0)] forvar605 = (1'h0);
  reg [(3'h5):(1'h0)] reg603 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg602 = (1'h0);
  reg [(5'h17):(1'h0)] reg601 = (1'h0);
  reg [(4'ha):(1'h0)] reg599 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg598 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar597 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg593 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg592 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar591 = (1'h0);
  reg [(5'h17):(1'h0)] reg589 = (1'h0);
  reg [(2'h3):(1'h0)] reg587 = (1'h0);
  reg [(5'h10):(1'h0)] forvar586 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar584 = (1'h0);
  reg [(2'h3):(1'h0)] reg584 = (1'h0);
  reg [(4'hf):(1'h0)] reg582 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg579 = (1'h0);
  reg [(4'h9):(1'h0)] reg578 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg576 = (1'h0);
  reg [(3'h6):(1'h0)] reg575 = (1'h0);
  reg [(5'h18):(1'h0)] reg573 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg572 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg571 = (1'h0);
  reg [(5'h16):(1'h0)] reg570 = (1'h0);
  reg [(5'h15):(1'h0)] reg569 = (1'h0);
  reg [(5'h1d):(1'h0)] reg568 = (1'h0);
  reg [(2'h2):(1'h0)] reg564 = (1'h0);
  reg [(4'hb):(1'h0)] reg563 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg561 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg560 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg554 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar551 = (1'h0);
  reg [(3'h4):(1'h0)] forvar550 = (1'h0);
  reg [(4'hb):(1'h0)] reg548 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar543 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg542 = (1'h0);
  reg [(4'hf):(1'h0)] reg541 = (1'h0);
  reg [(3'h5):(1'h0)] reg540 = (1'h0);
  reg [(5'h16):(1'h0)] reg539 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg534 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar531 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg530 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg529 = (1'h0);
  reg [(2'h3):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar526 = (1'h0);
  reg [(5'h19):(1'h0)] reg524 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg523 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar522 = (1'h0);
  reg [(4'ha):(1'h0)] reg520 = (1'h0);
  reg [(3'h7):(1'h0)] reg519 = (1'h0);
  reg [(2'h2):(1'h0)] reg518 = (1'h0);
  reg [(5'h1a):(1'h0)] reg515 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar514 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg512 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg508 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar507 = (1'h0);
  reg [(5'h13):(1'h0)] reg503 = (1'h0);
  reg [(5'h14):(1'h0)] reg501 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg500 = (1'h0);
  reg [(4'hd):(1'h0)] reg498 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar497 = (1'h0);
  reg [(4'h9):(1'h0)] reg495 = (1'h0);
  reg [(5'h14):(1'h0)] forvar491 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg490 = (1'h0);
  reg [(4'h9):(1'h0)] reg489 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg488 = (1'h0);
  reg [(5'h10):(1'h0)] forvar487 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg485 = (1'h0);
  reg [(4'hc):(1'h0)] forvar484 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg482 = (1'h0);
  reg [(3'h5):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg479 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg478 = (1'h0);
  reg [(5'h19):(1'h0)] reg475 = (1'h0);
  reg [(5'h17):(1'h0)] reg474 = (1'h0);
  reg [(5'h17):(1'h0)] forvar472 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar455 = (1'h0);
  reg [(3'h4):(1'h0)] forvar448 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar441 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar460 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg459 = (1'h0);
  reg [(5'h1b):(1'h0)] reg457 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg455 = (1'h0);
  reg [(3'h5):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg452 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg450 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg447 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg445 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg444 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg442 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg439 = (1'h0);
  reg [(5'h17):(1'h0)] forvar437 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg436 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar433 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg432 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg430 = (1'h0);
  reg [(5'h1b):(1'h0)] reg429 = (1'h0);
  reg [(3'h6):(1'h0)] forvar428 = (1'h0);
  reg [(5'h1d):(1'h0)] reg425 = (1'h0);
  reg [(5'h1b):(1'h0)] reg423 = (1'h0);
  reg [(5'h12):(1'h0)] forvar421 = (1'h0);
  reg [(3'h6):(1'h0)] forvar407 = (1'h0);
  reg [(5'h1b):(1'h0)] reg420 = (1'h0);
  reg [(4'hd):(1'h0)] reg417 = (1'h0);
  reg [(4'h8):(1'h0)] reg416 = (1'h0);
  reg [(3'h6):(1'h0)] reg415 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg413 = (1'h0);
  reg [(5'h12):(1'h0)] reg411 = (1'h0);
  reg [(5'h19):(1'h0)] reg407 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg399 = (1'h0);
  reg [(3'h5):(1'h0)] reg405 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg403 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar399 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg397 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg391 = (1'h0);
  reg [(3'h6):(1'h0)] reg390 = (1'h0);
  reg [(5'h1e):(1'h0)] reg389 = (1'h0);
  reg [(5'h1f):(1'h0)] reg388 = (1'h0);
  reg [(4'hd):(1'h0)] reg386 = (1'h0);
  reg [(5'h12):(1'h0)] reg385 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg384 = (1'h0);
  reg [(4'hc):(1'h0)] forvar374 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg379 = (1'h0);
  reg [(5'h1b):(1'h0)] reg378 = (1'h0);
  reg [(5'h17):(1'h0)] reg377 = (1'h0);
  reg [(4'hf):(1'h0)] forvar376 = (1'h0);
  reg [(3'h4):(1'h0)] reg375 = (1'h0);
  reg [(5'h15):(1'h0)] reg374 = (1'h0);
  reg [(5'h17):(1'h0)] reg373 = (1'h0);
  reg [(4'ha):(1'h0)] reg372 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg368 = (1'h0);
  reg [(4'hd):(1'h0)] reg366 = (1'h0);
  reg [(5'h17):(1'h0)] reg365 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar364 = (1'h0);
  reg [(5'h16):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg358 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg357 = (1'h0);
  reg [(4'hd):(1'h0)] reg356 = (1'h0);
  reg [(5'h13):(1'h0)] reg351 = (1'h0);
  reg [(4'hd):(1'h0)] reg350 = (1'h0);
  reg [(4'ha):(1'h0)] reg349 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg348 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar345 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar318 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg341 = (1'h0);
  reg [(5'h11):(1'h0)] forvar340 = (1'h0);
  reg [(5'h11):(1'h0)] forvar338 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg337 = (1'h0);
  reg [(4'hc):(1'h0)] reg335 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar334 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg333 = (1'h0);
  reg [(5'h19):(1'h0)] reg331 = (1'h0);
  reg [(5'h18):(1'h0)] forvar327 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg326 = (1'h0);
  reg [(5'h18):(1'h0)] reg325 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg323 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg319 = (1'h0);
  reg [(5'h16):(1'h0)] reg316 = (1'h0);
  reg [(5'h1e):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg312 = (1'h0);
  reg [(5'h1f):(1'h0)] reg310 = (1'h0);
  reg [(5'h1a):(1'h0)] reg308 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg306 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar305 = (1'h0);
  reg [(5'h1f):(1'h0)] reg304 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg303 = (1'h0);
  reg [(5'h14):(1'h0)] reg302 = (1'h0);
  reg [(4'ha):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar300 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg299 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg297 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar295 = (1'h0);
  reg [(3'h7):(1'h0)] reg292 = (1'h0);
  reg [(3'h6):(1'h0)] reg290 = (1'h0);
  reg [(5'h1c):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar285 = (1'h0);
  reg [(5'h19):(1'h0)] reg283 = (1'h0);
  reg [(3'h4):(1'h0)] reg282 = (1'h0);
  reg [(5'h12):(1'h0)] reg278 = (1'h0);
  reg [(4'hf):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg272 = (1'h0);
  reg [(4'h9):(1'h0)] reg271 = (1'h0);
  reg signed [(4'he):(1'h0)] reg269 = (1'h0);
  reg [(3'h6):(1'h0)] forvar267 = (1'h0);
  reg [(4'hc):(1'h0)] reg261 = (1'h0);
  reg [(4'hb):(1'h0)] forvar259 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar248 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg247 = (1'h0);
  reg [(5'h1b):(1'h0)] reg245 = (1'h0);
  reg [(5'h18):(1'h0)] reg244 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar243 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg242 = (1'h0);
  reg [(4'hf):(1'h0)] reg240 = (1'h0);
  reg [(5'h1a):(1'h0)] reg238 = (1'h0);
  reg [(4'he):(1'h0)] forvar237 = (1'h0);
  reg [(4'hb):(1'h0)] reg235 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar234 = (1'h0);
  reg [(5'h18):(1'h0)] reg231 = (1'h0);
  reg [(5'h1b):(1'h0)] reg230 = (1'h0);
  reg [(3'h5):(1'h0)] reg228 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar225 = (1'h0);
  reg [(5'h16):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg222 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar221 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar220 = (1'h0);
  reg [(3'h7):(1'h0)] reg217 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg214 = (1'h0);
  reg [(5'h12):(1'h0)] reg209 = (1'h0);
  reg [(5'h1a):(1'h0)] reg207 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg199 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar198 = (1'h0);
  reg [(5'h12):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg201 = (1'h0);
  reg [(4'ha):(1'h0)] reg200 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar199 = (1'h0);
  reg [(5'h17):(1'h0)] reg198 = (1'h0);
  reg [(3'h5):(1'h0)] reg197 = (1'h0);
  reg [(5'h1d):(1'h0)] reg196 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar195 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg194 = (1'h0);
  reg [(4'hb):(1'h0)] reg193 = (1'h0);
  reg [(5'h1c):(1'h0)] reg190 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg188 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar185 = (1'h0);
  reg [(2'h3):(1'h0)] reg184 = (1'h0);
  reg [(2'h3):(1'h0)] reg183 = (1'h0);
  reg signed [(4'he):(1'h0)] reg181 = (1'h0);
  reg [(4'hd):(1'h0)] reg180 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg177 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg172 = (1'h0);
  reg [(5'h11):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar170 = (1'h0);
  reg [(5'h1e):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg168 = (1'h0);
  reg [(5'h10):(1'h0)] forvar165 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg163 = (1'h0);
  reg [(5'h14):(1'h0)] forvar161 = (1'h0);
  reg [(4'h9):(1'h0)] reg160 = (1'h0);
  reg [(3'h6):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar152 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg151 = (1'h0);
  reg [(4'ha):(1'h0)] reg147 = (1'h0);
  reg [(2'h2):(1'h0)] reg145 = (1'h0);
  reg [(4'hc):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg140 = (1'h0);
  reg [(3'h5):(1'h0)] reg138 = (1'h0);
  reg [(4'hb):(1'h0)] reg137 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg135 = (1'h0);
  reg [(5'h1d):(1'h0)] reg133 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar132 = (1'h0);
  reg [(5'h11):(1'h0)] reg131 = (1'h0);
  reg [(3'h6):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg129 = (1'h0);
  reg [(3'h6):(1'h0)] reg126 = (1'h0);
  reg [(3'h5):(1'h0)] forvar123 = (1'h0);
  reg [(3'h6):(1'h0)] reg118 = (1'h0);
  reg [(4'he):(1'h0)] reg117 = (1'h0);
  reg [(5'h1b):(1'h0)] reg116 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg113 = (1'h0);
  reg [(4'hf):(1'h0)] reg112 = (1'h0);
  reg [(5'h17):(1'h0)] reg111 = (1'h0);
  reg [(5'h15):(1'h0)] reg110 = (1'h0);
  reg [(5'h1e):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg108 = (1'h0);
  reg [(5'h11):(1'h0)] reg106 = (1'h0);
  reg [(4'h9):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar103 = (1'h0);
  reg [(5'h17):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg100 = (1'h0);
  reg [(5'h13):(1'h0)] reg98 = (1'h0);
  reg [(5'h14):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg93 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg91 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg90 = (1'h0);
  reg [(4'he):(1'h0)] forvar89 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar86 = (1'h0);
  assign y = {wire617,
                 wire525,
                 wire511,
                 wire471,
                 wire470,
                 wire469,
                 wire468,
                 wire467,
                 wire344,
                 wire266,
                 wire265,
                 wire233,
                 wire121,
                 wire83,
                 reg616,
                 reg614,
                 reg609,
                 reg608,
                 reg607,
                 reg604,
                 reg600,
                 reg596,
                 reg595,
                 reg594,
                 reg590,
                 reg588,
                 reg585,
                 reg583,
                 reg581,
                 reg580,
                 reg577,
                 reg574,
                 reg567,
                 reg566,
                 reg565,
                 reg562,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg553,
                 reg552,
                 reg549,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 reg533,
                 reg532,
                 reg528,
                 reg521,
                 reg517,
                 reg516,
                 reg513,
                 reg510,
                 reg506,
                 reg505,
                 reg504,
                 reg502,
                 reg499,
                 reg496,
                 reg494,
                 reg493,
                 reg492,
                 reg486,
                 reg483,
                 reg481,
                 reg477,
                 reg476,
                 reg473,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg458,
                 reg456,
                 reg453,
                 reg451,
                 reg449,
                 reg448,
                 reg446,
                 reg443,
                 reg441,
                 reg440,
                 reg437,
                 reg438,
                 reg435,
                 reg434,
                 reg431,
                 reg427,
                 reg426,
                 reg424,
                 reg422,
                 reg421,
                 reg419,
                 reg418,
                 reg412,
                 reg410,
                 reg409,
                 reg408,
                 reg406,
                 reg404,
                 reg402,
                 reg400,
                 reg398,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg387,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg376,
                 reg371,
                 reg370,
                 reg369,
                 reg367,
                 reg363,
                 reg362,
                 reg361,
                 reg359,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg347,
                 reg346,
                 reg343,
                 reg342,
                 reg339,
                 reg336,
                 reg332,
                 reg330,
                 reg329,
                 reg328,
                 reg324,
                 reg322,
                 reg321,
                 reg320,
                 reg318,
                 reg317,
                 reg313,
                 reg311,
                 reg309,
                 reg307,
                 reg298,
                 reg294,
                 reg293,
                 reg291,
                 reg289,
                 reg288,
                 reg286,
                 reg285,
                 reg284,
                 reg281,
                 reg280,
                 reg279,
                 reg277,
                 reg275,
                 reg274,
                 reg270,
                 reg268,
                 reg264,
                 reg263,
                 reg262,
                 reg260,
                 reg258,
                 reg255,
                 reg254,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg246,
                 reg241,
                 reg239,
                 reg236,
                 reg232,
                 reg229,
                 reg227,
                 reg226,
                 reg224,
                 reg219,
                 reg218,
                 reg216,
                 reg215,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg208,
                 reg206,
                 reg205,
                 reg203,
                 reg202,
                 reg192,
                 reg191,
                 reg189,
                 reg187,
                 reg186,
                 reg182,
                 reg178,
                 reg175,
                 reg174,
                 reg167,
                 reg166,
                 reg164,
                 reg162,
                 reg157,
                 reg156,
                 reg154,
                 reg153,
                 reg150,
                 reg149,
                 reg148,
                 reg146,
                 reg143,
                 reg142,
                 reg139,
                 reg136,
                 reg134,
                 reg128,
                 reg127,
                 reg125,
                 reg124,
                 reg122,
                 reg120,
                 reg119,
                 reg115,
                 reg114,
                 reg107,
                 reg105,
                 reg101,
                 reg99,
                 reg97,
                 reg96,
                 reg95,
                 reg92,
                 reg88,
                 reg87,
                 reg85,
                 reg84,
                 reg615,
                 reg613,
                 forvar612,
                 forvar611,
                 reg610,
                 reg606,
                 forvar605,
                 reg603,
                 reg602,
                 reg601,
                 reg599,
                 reg598,
                 forvar597,
                 reg593,
                 reg592,
                 forvar591,
                 reg589,
                 reg587,
                 forvar586,
                 forvar584,
                 reg584,
                 reg582,
                 reg579,
                 reg578,
                 reg576,
                 reg575,
                 reg573,
                 reg572,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 reg564,
                 reg563,
                 reg561,
                 reg560,
                 reg559,
                 reg554,
                 forvar551,
                 forvar550,
                 reg548,
                 forvar543,
                 reg542,
                 reg541,
                 reg540,
                 reg539,
                 reg534,
                 forvar531,
                 reg530,
                 reg529,
                 reg527,
                 forvar526,
                 reg524,
                 reg523,
                 forvar522,
                 reg520,
                 reg519,
                 reg518,
                 reg515,
                 forvar514,
                 reg512,
                 reg509,
                 reg508,
                 forvar507,
                 reg503,
                 reg501,
                 reg500,
                 reg498,
                 forvar497,
                 reg495,
                 forvar491,
                 reg490,
                 reg489,
                 reg488,
                 forvar487,
                 reg485,
                 forvar484,
                 reg482,
                 reg480,
                 reg479,
                 reg478,
                 reg475,
                 reg474,
                 forvar472,
                 forvar455,
                 forvar448,
                 forvar441,
                 forvar460,
                 reg459,
                 reg457,
                 reg455,
                 reg454,
                 reg452,
                 reg450,
                 reg447,
                 reg445,
                 reg444,
                 reg442,
                 reg433,
                 reg439,
                 forvar437,
                 reg436,
                 forvar433,
                 reg432,
                 reg430,
                 reg429,
                 forvar428,
                 reg425,
                 reg423,
                 forvar421,
                 forvar407,
                 reg420,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg411,
                 reg407,
                 reg399,
                 reg405,
                 reg403,
                 reg401,
                 forvar399,
                 reg397,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg386,
                 reg385,
                 reg384,
                 forvar374,
                 reg379,
                 reg378,
                 reg377,
                 forvar376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg368,
                 reg366,
                 reg365,
                 forvar364,
                 reg360,
                 reg358,
                 reg357,
                 reg356,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 forvar345,
                 forvar318,
                 reg341,
                 forvar340,
                 forvar338,
                 reg337,
                 reg335,
                 forvar334,
                 reg333,
                 reg331,
                 forvar327,
                 reg326,
                 reg325,
                 reg323,
                 reg319,
                 reg316,
                 reg315,
                 reg314,
                 reg312,
                 reg310,
                 reg308,
                 reg306,
                 forvar305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 forvar300,
                 reg299,
                 reg297,
                 reg296,
                 forvar295,
                 reg292,
                 reg290,
                 reg287,
                 forvar285,
                 reg283,
                 reg282,
                 reg278,
                 reg276,
                 reg273,
                 reg272,
                 reg271,
                 reg269,
                 forvar267,
                 reg261,
                 forvar259,
                 reg257,
                 reg256,
                 reg253,
                 forvar248,
                 reg247,
                 reg245,
                 reg244,
                 forvar243,
                 reg242,
                 reg240,
                 reg238,
                 forvar237,
                 reg235,
                 forvar234,
                 reg231,
                 reg230,
                 reg228,
                 forvar225,
                 reg223,
                 reg222,
                 forvar221,
                 forvar220,
                 reg217,
                 reg214,
                 reg209,
                 reg207,
                 reg199,
                 forvar198,
                 reg204,
                 reg201,
                 reg200,
                 forvar199,
                 reg198,
                 reg197,
                 reg196,
                 forvar195,
                 reg194,
                 reg193,
                 reg190,
                 reg188,
                 forvar185,
                 reg184,
                 reg183,
                 reg181,
                 reg180,
                 reg179,
                 reg177,
                 reg176,
                 reg173,
                 reg172,
                 reg171,
                 forvar170,
                 reg169,
                 reg168,
                 forvar165,
                 reg163,
                 forvar161,
                 reg160,
                 reg159,
                 reg158,
                 reg155,
                 forvar152,
                 reg151,
                 reg147,
                 reg145,
                 reg144,
                 reg141,
                 reg140,
                 reg138,
                 reg137,
                 reg135,
                 reg133,
                 forvar132,
                 reg131,
                 reg130,
                 reg129,
                 reg126,
                 forvar123,
                 reg118,
                 reg117,
                 reg116,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg106,
                 reg104,
                 forvar103,
                 reg102,
                 reg100,
                 reg98,
                 reg94,
                 reg93,
                 reg91,
                 reg90,
                 forvar89,
                 forvar86,
                 (1'h0)};
  assign wire83 = wire79[(3'h5):(3'h4)];
  always
    @(posedge clk) begin
      reg84 <= wire83[(5'h11):(4'hc)];
      reg85 <= $signed({$signed({$signed(reg84)}),
          (|(wire79 >> $signed(wire79)))});
      for (forvar86 = (1'h0); (forvar86 < (3'h4)); forvar86 = (forvar86 + (1'h1)))
        begin
          reg87 <= {wire82,
              $signed(($unsigned($unsigned(wire79)) >= $signed($signed(reg85))))};
          reg88 <= reg84;
          for (forvar89 = (1'h0); (forvar89 < (3'h6)); forvar89 = (forvar89 + (1'h1)))
            begin
              reg90 = wire79;
              reg91 = reg85[(3'h5):(2'h3)];
              reg92 <= (~((wire79 ?
                  {wire83,
                      (+reg84)} : ($unsigned(wire83) - $signed(wire82))) ^~ (~^wire83)));
              reg93 = wire79;
              reg94 = (|(reg90 ?
                  reg84[(5'h16):(4'ha)] : (wire81 ?
                      (((8'h9c) ? wire81 : reg90) ?
                          (wire78 ?
                              reg93 : reg91) : $signed(forvar89)) : $signed((|reg93)))));
              reg95 <= (+reg88);
              reg96 <= (!((|((~forvar89) * reg88[(3'h7):(3'h6)])) ?
                  (wire80[(5'h12):(3'h6)] + {reg90,
                      (|reg87),
                      forvar86[(2'h3):(1'h0)]}) : wire78));
            end
          if (((|(reg85 || $signed((reg92 ? wire83 : wire79)))) + reg92))
            begin
              reg97 <= (7'h58);
              reg98 = $signed($signed((((reg95 ?
                  wire82 : wire80) - (~&wire80)) << $signed((wire82 ?
                  forvar86 : reg84)))));
            end
          else
            begin
              reg97 <= reg91[(3'h5):(2'h3)];
              reg99 <= $unsigned(forvar86[(3'h4):(3'h4)]);
              reg100 = reg84;
              reg101 <= (~(^~$unsigned($unsigned((&wire83)))));
              reg102 = {(^$unsigned(reg85[(2'h3):(1'h0)])),
                  $signed((($signed((8'ha3)) == $unsigned(forvar86)) ?
                      $unsigned((!reg100)) : wire83))};
            end
          for (forvar103 = (1'h0); (forvar103 < (3'h4)); forvar103 = (forvar103 + (1'h1)))
            begin
              reg104 = ((reg102 ?
                      $signed(($signed((8'had)) ~^ reg87[(4'hc):(4'h8)])) : (reg102[(5'h16):(4'hc)] ?
                          {$signed(reg95)} : $signed((wire81 ?
                              wire81 : wire83)))) ?
                  $unsigned(((((8'hb5) ~^ reg84) && {reg88,
                      forvar86}) != {$signed(wire81)})) : (reg96[(4'h8):(3'h6)] <<< reg92));
              reg105 <= (reg100 >= $signed($signed((reg85[(3'h7):(3'h5)] <<< (reg104 || reg85)))));
              reg106 = (~|{{$signed((~&wire82)),
                      reg105[(3'h6):(2'h3)],
                      $signed(reg96[(4'hf):(4'h8)])},
                  ($signed($unsigned((8'ha7))) || wire80)});
              reg107 <= ($unsigned($unsigned(reg93)) ^~ {(^~(reg93[(4'h8):(2'h3)] ?
                      (wire81 >= wire82) : $unsigned(forvar89))),
                  $signed($unsigned(wire83)),
                  $signed(reg94)});
              reg108 = (!(~&$unsigned(reg104[(4'h9):(3'h6)])));
            end
          if ($unsigned((wire79[(4'h9):(2'h2)] <= reg93)))
            begin
              reg109 = {$signed($signed((~^{wire82, (8'hac), reg107})))};
              reg110 = $unsigned(({wire80[(4'h9):(3'h4)]} | reg99));
              reg111 = wire79;
              reg112 = $unsigned(wire79[(3'h6):(3'h6)]);
              reg113 = (((8'hb7) <= $signed($signed({reg108}))) + wire82[(1'h1):(1'h0)]);
              reg114 <= reg93[(3'h7):(2'h3)];
            end
          else
            begin
              reg114 <= $unsigned($signed({$signed($unsigned(reg107))}));
              reg115 <= $signed($signed({reg110[(2'h3):(2'h2)]}));
              reg116 = $unsigned(wire78);
              reg117 = ((wire81[(3'h5):(3'h4)] ?
                  reg97 : $unsigned(reg101[(3'h6):(2'h2)])) - $signed((($signed(reg100) * reg100[(3'h5):(3'h4)]) ?
                  reg115 : $signed(reg111))));
              reg118 = (^reg114);
              reg119 <= ((~|({$unsigned((8'had)),
                      $unsigned(reg118),
                      (wire81 || (7'h51))} ?
                  ((~|(8'hbd)) ?
                      (-(8'hab)) : $signed(reg104)) : {(8'hbc)})) - reg97[(2'h2):(2'h2)]);
              reg120 <= $unsigned($unsigned($unsigned(reg109[(4'hf):(1'h1)])));
            end
        end
    end
  assign wire121 = (reg97 >> $signed((wire78 ?
                       (|$signed(reg96)) : $unsigned(reg87[(4'h9):(3'h7)]))));
  always
    @(posedge clk) begin
      reg122 <= reg84[(1'h1):(1'h0)];
      for (forvar123 = (1'h0); (forvar123 < (1'h0)); forvar123 = (forvar123 + (1'h1)))
        begin
          reg124 <= $signed(((((wire81 ?
              wire81 : reg84) ^ {reg119}) < $unsigned(wire121)) * wire82[(4'hb):(3'h4)]));
          reg125 <= ($signed((({reg95,
              (8'h9d)} - reg97) * $signed($unsigned(wire83)))) >>> (reg107[(3'h5):(2'h2)] || wire78));
        end
      if ({reg96[(4'hc):(3'h5)]})
        begin
          if ($signed(reg124[(1'h0):(1'h0)]))
            begin
              reg126 = $signed((((reg95 ? {wire81} : (reg120 ^ reg84)) ?
                  reg87[(3'h5):(1'h0)] : (reg96 ?
                      {reg96,
                          (7'h4e),
                          reg105} : $unsigned(reg114))) == (&(reg124 >> wire121[(4'hb):(4'ha)]))));
            end
          else
            begin
              reg127 <= (7'h4c);
              reg128 <= wire81[(5'h13):(5'h11)];
              reg129 = (wire83 - (^~($signed(reg122[(5'h19):(5'h17)]) ?
                  ($signed(reg105) ?
                      (reg119 ?
                          reg124 : reg107) : $signed((7'h53))) : reg125)));
              reg130 = reg119[(1'h1):(1'h0)];
              reg131 = (&{$unsigned($signed((^reg88))),
                  $signed({(reg96 * reg101)}),
                  (&reg84)});
            end
          for (forvar132 = (1'h0); (forvar132 < (1'h0)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 = $signed(reg129);
              reg134 <= ((($unsigned((!reg105)) + $signed({(7'h52)})) && wire81[(5'h11):(3'h6)]) ?
                  forvar132 : ($signed($signed($signed((7'h51)))) ?
                      wire83 : {$unsigned((~^reg115)),
                          {(forvar123 ? (8'ha1) : (8'ha9))}}));
              reg135 = reg124[(1'h0):(1'h0)];
              reg136 <= reg87[(4'hc):(4'h9)];
              reg137 = $unsigned($unsigned(((~reg124) != wire121)));
              reg138 = (!($unsigned({reg130}) & (+(!(~^reg96)))));
              reg139 <= reg135;
            end
          reg140 = (($signed($signed($signed((7'h4a)))) ?
              (reg122[(5'h1c):(4'h9)] <<< reg114) : $signed(wire78[(2'h3):(1'h1)])) && reg92);
          if ($unsigned((^(((|reg133) ? $unsigned(reg134) : wire82) - reg128))))
            begin
              reg141 = reg92;
              reg142 <= $signed((!(~&wire78)));
              reg143 <= $unsigned((~|$signed(((wire81 < wire82) ~^ (~reg115)))));
              reg144 = reg137;
            end
          else
            begin
              reg141 = (7'h4a);
              reg144 = reg131[(4'hb):(2'h3)];
              reg145 = (reg140 ^ {(wire78[(4'hb):(2'h2)] ?
                      (+(^~wire82)) : $signed(reg138[(2'h3):(2'h3)])),
                  $signed($unsigned(((8'hbb) == reg107))),
                  (|$unsigned(reg101))});
            end
          reg146 <= $signed(reg144);
          if (((wire83[(3'h4):(3'h4)] << (&reg84[(4'h8):(3'h7)])) <<< $signed((forvar132[(4'ha):(3'h4)] ?
              $unsigned($unsigned((8'ha8))) : $signed((~^reg135))))))
            begin
              reg147 = forvar132[(5'h19):(5'h16)];
              reg148 <= $signed(reg134[(4'hd):(4'hb)]);
              reg149 <= $unsigned(((!$signed($signed(forvar123))) ?
                  (|reg142[(1'h1):(1'h0)]) : (!$unsigned(reg144))));
              reg150 <= $unsigned($signed(($unsigned({reg136, forvar123}) ?
                  (7'h4b) : reg146)));
              reg151 = $unsigned((reg139[(4'he):(4'h8)] & ((^~$signed(reg134)) ?
                  $unsigned(reg122) : ((reg143 ? reg97 : reg125) == (8'hb4)))));
            end
          else
            begin
              reg147 = ((~^$signed({$unsigned(reg148),
                  (reg130 ^~ reg125)})) ^ wire78[(2'h2):(1'h1)]);
              reg148 <= $signed((-(^reg143)));
              reg151 = $unsigned(($unsigned($unsigned($signed((7'h43)))) ?
                  (reg87[(4'h9):(3'h5)] + reg137[(3'h4):(2'h3)]) : (7'h49)));
            end
        end
      else
        begin
          reg126 = reg126;
          reg127 <= {{$unsigned($signed($unsigned(reg107))),
                  (~^{(reg101 >> reg96), reg148})},
              (((reg101 ?
                      reg126[(2'h2):(1'h0)] : (~^reg126)) == $signed($signed((8'ha5)))) ?
                  {((reg88 > reg140) && {reg140}),
                      ($signed(forvar123) <<< $unsigned((7'h53)))} : (((forvar132 ?
                          reg142 : reg139) ?
                      reg115[(3'h6):(3'h6)] : (+reg122)) & (~|$signed(reg85)))),
              (+(((reg105 << reg88) | (7'h42)) ~^ reg88[(3'h5):(2'h3)]))};
        end
    end
  always
    @(posedge clk) begin
      for (forvar152 = (1'h0); (forvar152 < (2'h2)); forvar152 = (forvar152 + (1'h1)))
        begin
          if ((!$signed($signed($signed(reg127[(3'h7):(3'h4)])))))
            begin
              reg153 <= ((wire79[(4'h8):(3'h6)] & (reg127 >= ({(8'ha4),
                          reg146} ?
                      (reg99 ? (8'haa) : (8'h9f)) : $signed(reg124)))) ?
                  reg124[(1'h0):(1'h0)] : (({(!(7'h40))} ?
                          (7'h40) : reg143[(1'h0):(1'h0)]) ?
                      reg127 : (-({reg119, wire82} ^ (reg119 ?
                          reg99 : reg96)))));
              reg154 <= ((($signed(wire79[(1'h0):(1'h0)]) ?
                          $unsigned($signed(reg124)) : reg136[(4'hb):(4'hb)]) ?
                      reg96[(5'h10):(1'h0)] : $signed(($signed(reg95) ?
                          {(7'h4a), (8'hbc)} : (reg85 < reg85)))) ?
                  wire82[(4'hb):(2'h3)] : $unsigned({reg146[(4'hb):(3'h5)],
                      reg136}));
              reg155 = (reg114 && (|$unsigned($unsigned((!(8'h9f))))));
              reg156 <= ($signed({({wire80, reg128} ?
                          $signed((7'h52)) : (reg97 - wire83)),
                      $signed((^reg114))}) ?
                  (reg143 <<< reg146) : (reg139 >= $signed((reg155[(3'h6):(1'h0)] + (~&reg127)))));
              reg157 <= $signed((($unsigned((~^reg128)) ?
                  ((-(8'hb0)) < {reg155,
                      reg148,
                      reg119}) : reg107) < ({$unsigned(reg114),
                  {reg156, reg124}} < $signed($unsigned(reg136)))));
              reg158 = ($signed(reg150[(2'h3):(2'h3)]) ? reg105 : reg96);
              reg159 = reg85[(3'h6):(3'h6)];
            end
          else
            begin
              reg153 <= (^~(8'hbc));
              reg155 = wire79;
              reg158 = reg107[(5'h10):(1'h0)];
              reg159 = $unsigned(({{{(8'ha6)},
                      reg150[(1'h1):(1'h1)]}} & reg128[(5'h10):(4'h8)]));
            end
          reg160 = $signed(reg142);
          for (forvar161 = (1'h0); (forvar161 < (3'h5)); forvar161 = (forvar161 + (1'h1)))
            begin
              reg162 <= ((+((reg128[(5'h12):(2'h2)] ?
                      reg146[(3'h4):(2'h3)] : $unsigned(wire82)) ?
                  $unsigned((^reg119)) : reg156)) != reg95);
              reg163 = (8'ha5);
              reg164 <= reg96[(4'he):(1'h1)];
            end
        end
      for (forvar165 = (1'h0); (forvar165 < (3'h5)); forvar165 = (forvar165 + (1'h1)))
        begin
          reg166 <= $unsigned(($signed(wire81) ?
              (8'ha4) : {($unsigned((7'h55)) ?
                      ((7'h42) ? forvar161 : forvar165) : (reg125 ?
                          reg95 : (8'hb0)))}));
          if ($unsigned(reg150[(2'h3):(1'h0)]))
            begin
              reg167 <= (|((reg97 ?
                      ((~^reg146) ?
                          {reg154} : reg96[(4'he):(4'h8)]) : (-(wire121 ?
                          (7'h52) : reg101))) ?
                  $unsigned($unsigned((|reg87))) : ($signed($signed(reg124)) ^ ($unsigned((8'hb2)) < reg114[(5'h12):(4'hf)]))));
              reg168 = (&reg160);
              reg169 = ((+((reg128[(2'h3):(2'h3)] - (reg134 ?
                      wire80 : wire82)) ?
                  ((~&reg107) * (|reg148)) : $signed(reg160[(4'h9):(2'h2)]))) && ($unsigned($unsigned(reg154[(1'h1):(1'h1)])) + ((7'h40) ^~ $unsigned((wire81 ?
                  (8'hb1) : wire78)))));
            end
          else
            begin
              reg167 <= (~|$unsigned(reg92[(5'h1b):(4'hc)]));
            end
          for (forvar170 = (1'h0); (forvar170 < (3'h4)); forvar170 = (forvar170 + (1'h1)))
            begin
              reg171 = reg153;
              reg172 = $signed((reg96 ?
                  (reg92 ?
                      reg164 : wire79[(2'h2):(1'h1)]) : $unsigned(wire81)));
              reg173 = ($signed(reg99) ?
                  (((+reg157[(3'h4):(2'h3)]) ?
                      ((|reg146) ?
                          $signed((8'h9d)) : (reg172 << reg134)) : {forvar165,
                          $signed(reg166)}) <<< $unsigned(reg159)) : (!$unsigned(reg107[(4'he):(1'h0)])));
              reg174 <= $unsigned((reg164 ?
                  ($signed((reg119 && forvar152)) ^ reg168[(4'hb):(1'h1)]) : forvar165[(4'ha):(1'h1)]));
              reg175 <= (^~(($signed((wire121 ^~ reg143)) ?
                      ((reg166 ?
                          wire121 : reg156) || wire80) : $unsigned({reg99,
                          reg136,
                          reg125})) ?
                  $unsigned(($signed(reg167) ?
                      (&forvar161) : (reg97 >= reg169))) : $signed(reg107)));
              reg176 = $unsigned((($signed(reg156[(4'he):(1'h0)]) ?
                  (reg159[(1'h0):(1'h0)] ?
                      reg163[(1'h1):(1'h1)] : $unsigned(reg167)) : reg169[(5'h1a):(5'h11)]) >>> reg156[(4'hf):(4'h8)]));
              reg177 = (($unsigned((~&(7'h54))) ?
                  ((+(8'h9c)) - {reg134,
                      reg163,
                      (^~reg125)}) : (((!(8'had)) == forvar170) ?
                      $unsigned({wire82,
                          reg146,
                          reg155}) : ($signed(forvar170) ?
                          ((8'ha4) ?
                              reg166 : (7'h52)) : $unsigned(reg142)))) > $signed($unsigned((((7'h45) & reg159) ?
                  reg85 : {wire80}))));
            end
          if ($unsigned((~&{reg119[(3'h7):(3'h4)]})))
            begin
              reg178 <= reg163[(1'h0):(1'h0)];
              reg179 = $signed(reg150);
              reg180 = reg169[(2'h2):(2'h2)];
              reg181 = reg163;
              reg182 <= ({wire121[(3'h4):(1'h1)]} ?
                  $signed((^$unsigned((reg92 + reg177)))) : $signed(reg153[(4'hf):(2'h2)]));
            end
          else
            begin
              reg179 = ((-(&($signed(reg167) < (~(7'h51))))) ?
                  reg128[(4'ha):(3'h5)] : reg119[(5'h19):(5'h16)]);
              reg180 = ($unsigned(($signed({reg150}) > (reg159 ?
                  (reg181 ?
                      (8'hba) : (8'ha5)) : reg119[(2'h2):(1'h1)]))) + reg149[(5'h13):(5'h13)]);
              reg182 <= {reg173};
            end
          reg183 = {reg169, $unsigned(reg99[(4'hc):(4'hb)]), reg119};
          reg184 = {(+$unsigned($signed($unsigned(reg128))))};
        end
      for (forvar185 = (1'h0); (forvar185 < (2'h2)); forvar185 = (forvar185 + (1'h1)))
        begin
          if ($unsigned($unsigned(reg178)))
            begin
              reg186 <= reg122[(5'h18):(5'h11)];
              reg187 <= reg107;
            end
          else
            begin
              reg188 = (($signed((forvar170[(1'h0):(1'h0)] && reg175)) == {({reg154} - reg174),
                      reg92[(4'ha):(3'h7)]}) ?
                  $signed($signed((^~{(7'h4d)}))) : $unsigned(wire79[(1'h1):(1'h1)]));
              reg189 <= reg188;
              reg190 = reg156;
              reg191 <= reg164[(5'h1b):(4'hf)];
              reg192 <= $unsigned(reg166);
              reg193 = (-$signed({reg184,
                  {reg182[(4'h9):(2'h3)], (reg157 ^ reg143)}}));
              reg194 = $signed(((reg175[(1'h1):(1'h1)] ?
                  (reg84[(5'h17):(5'h10)] ?
                      {reg163} : $unsigned(reg150)) : reg192[(5'h16):(3'h5)]) && ((^$unsigned(reg146)) ?
                  ((^~reg168) ?
                      $signed(reg171) : (reg146 ?
                          reg142 : reg155)) : ($signed(reg178) && {reg120,
                      reg163}))));
            end
          for (forvar195 = (1'h0); (forvar195 < (2'h2)); forvar195 = (forvar195 + (1'h1)))
            begin
              reg196 = reg187;
              reg197 = $unsigned(reg146[(4'hb):(2'h2)]);
            end
        end
      if ($signed($signed($unsigned(wire82))))
        begin
          reg198 = (~^$signed($signed(((!reg150) ? (8'hb7) : (8'had)))));
          for (forvar199 = (1'h0); (forvar199 < (2'h2)); forvar199 = (forvar199 + (1'h1)))
            begin
              reg200 = reg155;
              reg201 = reg114;
              reg202 <= (-wire83);
              reg203 <= (($unsigned(((~(8'hb0)) ?
                      (reg150 <<< reg196) : (~reg146))) || ((+((8'hb7) ?
                      reg87 : reg156)) == {(reg172 ? (7'h40) : (8'h9d))})) ?
                  (~&({{reg166,
                          forvar170,
                          reg200}} == reg169)) : ($signed(reg157) >> ((~((8'h9d) - reg175)) ?
                      forvar185[(1'h0):(1'h0)] : (~|$unsigned(reg191)))));
              reg204 = (~$signed(((wire81[(3'h4):(1'h1)] ?
                      (forvar185 ? reg166 : reg180) : (~^reg190)) ?
                  $unsigned((reg160 + (8'ha6))) : reg92[(2'h2):(1'h0)])));
              reg205 <= reg178[(4'hf):(3'h7)];
            end
          reg206 <= $unsigned((-{(!reg193[(3'h7):(1'h1)]),
              (-$unsigned((7'h48))),
              {((8'ha6) ? reg115 : (7'h42)),
                  forvar170,
                  reg164[(4'ha):(4'h9)]}}));
        end
      else
        begin
          for (forvar198 = (1'h0); (forvar198 < (2'h2)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 = (7'h53);
              reg200 = reg177;
            end
          if ({(7'h4d),
              (+$unsigned($signed({(8'hb3), (8'hb0), reg107}))),
              reg180[(4'hb):(1'h1)]})
            begin
              reg201 = reg197[(1'h0):(1'h0)];
              reg204 = (reg156 ?
                  $signed(reg95) : ({reg160[(4'h9):(2'h3)],
                      ((-reg92) || $signed(reg177))} ^ reg156));
              reg205 <= $unsigned((($unsigned($unsigned(reg162)) & reg198) ?
                  reg176 : $signed(wire78)));
            end
          else
            begin
              reg202 <= reg134[(2'h2):(1'h0)];
              reg204 = (+(^(((^~reg128) | $signed(wire82)) <<< $unsigned((8'ha9)))));
              reg207 = $unsigned(reg122[(2'h3):(2'h2)]);
              reg208 <= {($unsigned(((~^reg172) ?
                      (reg120 ?
                          reg200 : (7'h41)) : (reg95 >= (7'h50)))) ^~ reg169)};
              reg209 = {reg134,
                  ({$unsigned($unsigned(reg181))} ? reg88 : reg105),
                  $unsigned((~&reg169[(4'hf):(4'h9)]))};
              reg210 <= ($signed(forvar161[(3'h4):(2'h2)]) ?
                  $unsigned({reg197,
                      (reg188 ?
                          ((8'hb2) || reg153) : $unsigned(forvar152))}) : {reg96});
              reg211 <= (&(~|(8'hbf)));
            end
          if ((^~reg199))
            begin
              reg212 <= (^~$unsigned($signed((-$signed(reg204)))));
              reg213 <= {((&reg207[(4'hc):(4'hc)]) ?
                      reg180[(4'h9):(3'h7)] : (^~(&$unsigned(reg92)))),
                  (|($unsigned($signed(reg87)) ?
                      $unsigned((reg85 ^ reg119)) : {$signed(reg197)})),
                  {$signed(reg208),
                      (((8'had) ?
                          $signed((8'hae)) : (reg163 ?
                              (8'hae) : (7'h4a))) > $unsigned($signed(reg212))),
                      $signed({(~reg196),
                          $unsigned((7'h46)),
                          $unsigned((7'h43))})}};
              reg214 = reg194[(4'h8):(1'h1)];
              reg215 <= $signed((&(reg210 ? reg209[(4'hc):(4'hb)] : reg84)));
              reg216 <= $unsigned(reg183[(2'h2):(1'h1)]);
              reg217 = (reg186 ?
                  ((8'hb1) ?
                      $signed((~^(8'ha4))) : (~^$unsigned($unsigned((7'h49))))) : reg194[(3'h5):(1'h1)]);
              reg218 <= (wire83[(4'he):(4'h8)] ?
                  reg115[(2'h2):(1'h1)] : {(^(forvar152[(5'h15):(3'h7)] - $signed(reg160)))});
            end
          else
            begin
              reg214 = {{(^~($unsigned((7'h4d)) * $unsigned(reg143))),
                      $signed($unsigned({reg189, (7'h4c)}))}};
              reg215 <= $unsigned((^~(^$unsigned((8'hb6)))));
              reg217 = (~^reg202[(4'h8):(3'h7)]);
              reg218 <= ($signed(reg105) != $signed(reg99[(3'h4):(2'h3)]));
            end
        end
      reg219 <= reg154;
      for (forvar220 = (1'h0); (forvar220 < (2'h3)); forvar220 = (forvar220 + (1'h1)))
        begin
          for (forvar221 = (1'h0); (forvar221 < (3'h6)); forvar221 = (forvar221 + (1'h1)))
            begin
              reg222 = reg175[(3'h4):(1'h1)];
            end
          reg223 = reg218;
          reg224 <= {(8'hb0)};
          for (forvar225 = (1'h0); (forvar225 < (2'h2)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 <= (8'ha1);
              reg227 <= (8'hac);
              reg228 = reg196[(5'h18):(4'hc)];
              reg229 <= $unsigned(reg227);
            end
          reg230 = ({reg177} ?
              $unsigned($signed(reg157[(1'h0):(1'h0)])) : ($unsigned(($signed(reg219) & reg172)) ?
                  (((reg166 <= reg124) ?
                      {reg134} : reg172[(4'h9):(2'h2)]) || ((reg208 | (8'hbb)) <<< $signed(reg205))) : reg188));
        end
      reg231 = ($unsigned(reg85[(1'h0):(1'h0)]) != $signed({(!{reg213,
              reg199})}));
    end
  always
    @(posedge clk) begin
      reg232 <= $unsigned(reg157);
    end
  assign wire233 = $unsigned($unsigned($signed(reg150)));
  always
    @(posedge clk) begin
      for (forvar234 = (1'h0); (forvar234 < (3'h5)); forvar234 = (forvar234 + (1'h1)))
        begin
          reg235 = $unsigned($unsigned($signed({wire80[(4'ha):(4'h9)],
              reg136[(4'ha):(4'h8)],
              reg85})));
          reg236 <= (-reg175);
          for (forvar237 = (1'h0); (forvar237 < (1'h0)); forvar237 = (forvar237 + (1'h1)))
            begin
              reg238 = $unsigned((~(($signed(reg175) & $unsigned(wire78)) ?
                  wire83 : ($unsigned(reg122) || {reg101}))));
              reg239 <= reg127[(3'h6):(1'h0)];
              reg240 = $signed(reg97);
              reg241 <= (^~{(^~reg205)});
              reg242 = $unsigned(((($unsigned(wire233) ?
                          (wire121 ? (8'h9c) : wire78) : {wire121,
                              reg136,
                              (7'h40)}) ?
                      (8'hb6) : (|$signed(reg125))) ?
                  (reg205 ?
                      reg154 : ((reg143 ? reg125 : reg227) ?
                          (~^reg212) : reg240[(4'hc):(3'h5)])) : $signed(reg240[(4'h9):(1'h0)])));
            end
          for (forvar243 = (1'h0); (forvar243 < (1'h1)); forvar243 = (forvar243 + (1'h1)))
            begin
              reg244 = ((~reg115) ?
                  (~&{((~reg218) ? {wire80, reg239} : (reg226 - reg213)),
                      ((8'ha7) ?
                          $signed(reg206) : (reg162 ?
                              (8'ha2) : reg174))}) : {$signed($unsigned({reg186,
                          reg153})),
                      {$signed(((8'hb3) ~^ wire81)), (~|$unsigned(reg95))}});
              reg245 = reg95;
              reg246 <= $unsigned($unsigned($signed({$signed(reg227),
                  ((7'h56) * reg154),
                  reg146[(4'hd):(4'ha)]})));
              reg247 = reg240;
            end
        end
      for (forvar248 = (1'h0); (forvar248 < (3'h6)); forvar248 = (forvar248 + (1'h1)))
        begin
          reg249 <= $unsigned(forvar248);
          reg250 <= $signed((|reg229[(5'h12):(4'hb)]));
          reg251 <= reg107[(5'h19):(2'h3)];
          if (reg114[(4'he):(4'hb)])
            begin
              reg252 <= (-{($signed(reg87) ?
                      (reg251 ?
                          {(8'ha2),
                              (8'ha6),
                              (8'ha5)} : reg186[(3'h7):(3'h6)]) : {(reg241 - reg119),
                          reg215,
                          $unsigned(reg84)}),
                  reg84});
              reg253 = ($unsigned(reg95) * reg134);
              reg254 <= $signed(wire80[(5'h10):(2'h3)]);
              reg255 <= $unsigned((~&$signed((!$unsigned(reg240)))));
              reg256 = $unsigned((|($unsigned((^reg174)) ?
                  ($unsigned((8'hb3)) ^~ (7'h4f)) : $unsigned((reg119 ?
                      (8'ha2) : (8'hbc))))));
              reg257 = (reg97[(1'h1):(1'h0)] ?
                  ((wire121 ? (reg210 ? (8'ha2) : $signed(reg124)) : reg242) ?
                      $signed($signed($signed(reg240))) : reg235) : reg122);
            end
          else
            begin
              reg252 <= ($unsigned(reg154) ?
                  (+({reg101[(3'h7):(3'h6)],
                      (reg125 << (7'h4a))} < wire79[(2'h2):(2'h2)])) : $signed(((|((8'ha9) * reg211)) != $signed($signed(reg238)))));
            end
          reg258 <= reg92[(1'h0):(1'h0)];
          for (forvar259 = (1'h0); (forvar259 < (3'h6)); forvar259 = (forvar259 + (1'h1)))
            begin
              reg260 <= (reg136[(4'ha):(2'h2)] >= wire121);
              reg261 = ($unsigned({wire233,
                  ($signed(reg124) * (reg208 >>> reg191))}) & reg87);
            end
        end
      reg262 <= (reg157[(1'h1):(1'h0)] && {(~|$signed(reg261)),
          $signed((8'hbb)),
          (reg97 ~^ ((reg244 ? reg143 : reg260) <<< $unsigned(reg154)))});
      reg263 <= (((((reg246 << reg142) ? $signed(reg249) : {reg241, reg124}) ?
          reg236[(5'h15):(5'h12)] : (~{reg87,
              (8'ha2)})) >>> $unsigned((~|(reg120 ?
          reg99 : reg224)))) - reg251[(5'h10):(4'he)]);
      reg264 <= reg87;
    end
  assign wire265 = reg246;
  assign wire266 = wire233[(5'h11):(3'h4)];
  always
    @(posedge clk) begin
      for (forvar267 = (1'h0); (forvar267 < (3'h5)); forvar267 = (forvar267 + (1'h1)))
        begin
          if ($unsigned($signed(reg95)))
            begin
              reg268 <= ((($unsigned({(8'ha7), reg125}) << (~&{(8'hbd),
                      reg157})) ?
                  $unsigned({(reg224 ? reg213 : wire81),
                      $signed((8'had))}) : $unsigned($unsigned(reg162[(2'h2):(2'h2)]))) - (^(&(-((8'hab) ?
                  reg187 : reg239)))));
              reg269 = $signed($unsigned($signed($signed($signed((7'h46))))));
              reg270 <= $unsigned($signed($unsigned($unsigned($unsigned((8'hbf))))));
              reg271 = (7'h43);
              reg272 = (+wire265);
              reg273 = (reg178[(5'h16):(5'h12)] >= $signed($signed(($signed(reg97) >>> {reg95,
                  reg139,
                  reg139}))));
              reg274 <= $signed(reg206);
            end
          else
            begin
              reg268 <= wire233;
              reg270 <= $unsigned(($signed($signed(reg211)) > ({wire233[(3'h6):(3'h4)],
                      $unsigned((7'h50))} ?
                  reg88[(3'h7):(2'h2)] : ($signed(reg136) - $signed(reg178)))));
              reg271 = reg191[(5'h13):(3'h6)];
              reg274 <= $signed($signed(reg202));
              reg275 <= $unsigned($signed(((((8'had) ? reg142 : reg162) ?
                  $unsigned((8'ha3)) : $unsigned(reg174)) >= $signed((reg149 * reg213)))));
              reg276 = (~^$signed(reg164[(5'h14):(4'he)]));
            end
          reg277 <= ({$signed(reg254),
              $signed($signed(((8'hac) >>> reg178))),
              $unsigned(($signed(reg124) != reg84))} | (+reg219[(1'h0):(1'h0)]));
          reg278 = {$unsigned(wire83)};
          reg279 <= reg202[(4'h9):(1'h0)];
        end
      reg280 <= (reg136 ?
          (reg125[(4'h9):(3'h6)] ?
              reg148[(1'h0):(1'h0)] : reg255) : (&($unsigned((^reg134)) ?
              reg249 : $signed(reg175))));
      if ($signed($signed((&$unsigned((8'ha9))))))
        begin
          reg281 <= (^((^$signed({reg107, reg95, reg178})) ?
              ($unsigned(reg205[(3'h7):(2'h3)]) >= (~^$unsigned(reg227))) : $unsigned(reg272)));
          reg282 = (((-{((7'h58) <<< reg232),
                  (reg84 <= (7'h55)),
                  reg153}) * reg229[(1'h0):(1'h0)]) ?
              (~((!(reg139 ?
                  reg269 : (7'h41))) == $signed((&reg224)))) : ((($signed(reg136) ?
                  reg162 : ((7'h40) ?
                      reg211 : reg262)) || (!(reg136 >= reg164))) <= reg262));
          reg283 = $signed($unsigned(reg236));
          reg284 <= reg203;
          reg285 <= $signed($signed(reg271[(3'h6):(3'h4)]));
        end
      else
        begin
          reg281 <= (^$unsigned({reg277[(4'h8):(3'h7)]}));
          reg284 <= $signed(reg278);
          for (forvar285 = (1'h0); (forvar285 < (3'h6)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg286 <= $signed((&$signed(reg250[(4'h8):(2'h3)])));
              reg287 = $signed((+reg175));
              reg288 <= ({reg175[(1'h0):(1'h0)],
                  reg258} <= ((reg216 && reg269[(4'h8):(2'h2)]) ?
                  $signed(((^reg162) >> reg157[(1'h0):(1'h0)])) : reg202));
            end
          if (({reg208[(1'h0):(1'h0)],
                  $unsigned($signed(reg166[(1'h1):(1'h0)])),
                  $unsigned($signed(reg283[(1'h1):(1'h0)]))} ?
              (!(reg205[(3'h6):(1'h0)] ?
                  (~&((7'h46) ^ reg142)) : $signed((~^(8'h9f))))) : $unsigned(({$signed(wire82),
                  (reg226 + reg105),
                  (reg148 ? reg208 : reg208)} <= ({reg97,
                  reg279} != (8'haf))))))
            begin
              reg289 <= $signed((-(7'h4b)));
              reg290 = (reg218 ?
                  {$unsigned((reg156[(3'h4):(1'h1)] ?
                          $unsigned((7'h4d)) : (!wire78))),
                      ($unsigned((reg148 & reg186)) >= ((reg264 ?
                          reg139 : (7'h58)) <= reg97[(1'h1):(1'h1)]))} : (7'h47));
              reg291 <= reg215[(2'h3):(1'h1)];
              reg292 = reg254[(4'he):(3'h7)];
              reg293 <= reg271;
              reg294 <= $signed(($unsigned($signed($signed(wire80))) * $signed((7'h42))));
            end
          else
            begin
              reg289 <= {$signed($signed(reg128)),
                  reg125,
                  $unsigned(reg92[(2'h2):(1'h0)])};
              reg291 <= (&($signed(wire121) << reg150));
              reg292 = ((($unsigned((reg189 ? wire82 : reg232)) ?
                      $signed(reg254) : $unsigned({reg142,
                          forvar285})) != (reg293 || ($unsigned(reg134) ?
                      reg148[(1'h1):(1'h1)] : (^(7'h4c))))) ?
                  (({forvar267, reg232, reg290[(1'h1):(1'h0)]} ?
                      (reg287[(2'h3):(2'h3)] ?
                          (|reg175) : {reg279,
                              reg280,
                              reg270}) : ($unsigned(reg164) ?
                          reg293[(4'hf):(4'hc)] : reg119[(4'hf):(4'ha)])) == $unsigned(($signed((7'h43)) == reg268))) : $signed(reg229[(3'h5):(3'h4)]));
              reg293 <= {(&reg278)};
              reg294 <= $unsigned($signed((reg284[(5'h13):(1'h0)] ?
                  (!(+reg84)) : $unsigned((reg162 ? reg251 : reg215)))));
            end
          for (forvar295 = (1'h0); (forvar295 < (3'h4)); forvar295 = (forvar295 + (1'h1)))
            begin
              reg296 = (wire121 ?
                  $signed($signed({(reg150 ? (7'h4c) : reg166),
                      reg262[(4'h9):(3'h7)],
                      (~^(7'h50))})) : (7'h4c));
            end
          if ($signed(reg178[(5'h14):(3'h4)]))
            begin
              reg297 = (reg290 * reg287);
            end
          else
            begin
              reg298 <= ({wire80,
                  reg178,
                  $unsigned(((reg174 ?
                      reg97 : reg128) || $signed(reg281)))} == reg273[(4'hf):(4'h9)]);
              reg299 = (reg281 ? reg164 : $unsigned(reg96[(3'h7):(3'h4)]));
            end
        end
      for (forvar300 = (1'h0); (forvar300 < (3'h6)); forvar300 = (forvar300 + (1'h1)))
        begin
          if ($signed($unsigned((reg299[(3'h7):(3'h5)] ?
              {{reg270, forvar295, (8'hb5)}} : $signed({(7'h58)})))))
            begin
              reg301 = (7'h42);
              reg302 = (reg149 ?
                  $unsigned($unsigned(reg239)) : (^$unsigned({reg297[(2'h3):(2'h2)],
                      $signed(reg279),
                      (|reg298)})));
            end
          else
            begin
              reg301 = $unsigned(($unsigned($signed((^~reg255))) ?
                  (reg215[(3'h5):(1'h1)] ?
                      (~(^reg174)) : ((&reg269) ?
                          (reg226 ? reg250 : reg272) : {wire121,
                              reg291})) : $signed(reg114)));
              reg302 = (-$unsigned(reg280[(2'h2):(1'h1)]));
              reg303 = ((((7'h57) == wire265[(3'h7):(2'h3)]) ?
                  ($unsigned((reg284 < reg276)) ?
                      $signed(reg294) : $signed(reg202[(5'h17):(5'h15)])) : $signed($unsigned(reg142[(1'h0):(1'h0)]))) <<< ($signed($unsigned($unsigned(reg97))) ?
                  $signed(($unsigned(reg192) ?
                      (reg149 ?
                          reg232 : reg260) : reg271[(3'h4):(2'h2)])) : reg191[(3'h7):(3'h7)]));
              reg304 = $unsigned((^~$signed(reg241)));
            end
          for (forvar305 = (1'h0); (forvar305 < (3'h5)); forvar305 = (forvar305 + (1'h1)))
            begin
              reg306 = ($unsigned(((^~(reg251 ^ reg167)) ?
                      $unsigned((reg280 ?
                          wire82 : reg88)) : (~reg134[(3'h7):(1'h1)]))) ?
                  $signed({((forvar300 ? reg85 : reg212) ?
                          reg215[(5'h14):(4'hc)] : (-reg210))}) : (~reg128[(2'h2):(2'h2)]));
              reg307 <= {$signed($unsigned(reg303[(5'h12):(4'h8)])),
                  $signed($signed(reg241)),
                  ($unsigned((~&(-(8'h9e)))) ?
                      $unsigned({{reg148,
                              (7'h50)}}) : (+((reg92 < reg272) + (|reg134))))};
              reg308 = (&$signed((reg298[(4'hb):(2'h2)] | (reg232 ?
                  (reg290 < reg92) : $unsigned(reg218)))));
              reg309 <= (!$signed($unsigned(reg87)));
              reg310 = (reg270[(3'h4):(2'h3)] ?
                  (~(~|(!reg212))) : reg239[(5'h11):(4'hc)]);
            end
          reg311 <= wire266[(5'h10):(5'h10)];
          reg312 = ($unsigned(reg95[(3'h4):(1'h1)]) ?
              (-reg211[(4'hd):(3'h5)]) : ((($unsigned(reg202) && $signed(reg105)) ?
                      (-$unsigned(reg286)) : reg175[(2'h2):(1'h0)]) ?
                  ($unsigned(reg146) != {(wire233 ? reg226 : (8'hba)),
                      reg275[(3'h4):(1'h1)]}) : reg280[(1'h1):(1'h0)]));
        end
    end
  always
    @(posedge clk) begin
      reg313 <= ((^~(~|((~&reg298) ?
              (reg124 << reg249) : reg157[(3'h4):(2'h3)]))) ?
          wire80 : wire83[(1'h0):(1'h0)]);
      reg314 = reg275;
      reg315 = (reg213[(2'h2):(1'h1)] + reg252);
      reg316 = reg274[(5'h18):(5'h13)];
      reg317 <= (~^(reg316[(4'hd):(1'h0)] ?
          reg236[(2'h2):(1'h0)] : {wire79, ((-reg268) ^ reg85)}));
      if ((reg218[(5'h11):(3'h5)] ?
          $unsigned((~$unsigned(((8'ha5) ? reg143 : reg202)))) : (7'h40)))
        begin
          if ($signed(reg205[(4'hb):(1'h1)]))
            begin
              reg318 <= reg203;
              reg319 = reg274[(4'hf):(4'hc)];
              reg320 <= $signed(reg174);
              reg321 <= (reg120[(5'h1d):(5'h18)] ?
                  {reg87[(4'hb):(3'h7)]} : $unsigned(reg182[(4'hb):(3'h6)]));
              reg322 <= (~^$signed(($unsigned($unsigned(wire80)) << reg236[(5'h15):(4'h9)])));
              reg323 = (reg281[(4'ha):(2'h3)] != {wire78[(3'h6):(3'h5)],
                  $signed(reg128)});
              reg324 <= (~|$unsigned((reg119[(5'h10):(4'hc)] < $unsigned($signed((8'hb6))))));
            end
          else
            begin
              reg318 <= (~reg166[(4'h9):(4'h9)]);
              reg320 <= $signed((^(reg262[(5'h1b):(4'h8)] > reg311[(5'h14):(5'h11)])));
              reg323 = (8'hbd);
              reg325 = $signed($unsigned($signed(reg274)));
              reg326 = $signed(($unsigned($unsigned((^~reg139))) ?
                  $unsigned(reg224[(4'h8):(2'h2)]) : (~reg250)));
            end
          for (forvar327 = (1'h0); (forvar327 < (3'h4)); forvar327 = (forvar327 + (1'h1)))
            begin
              reg328 <= ($unsigned($signed(reg277)) >= (reg250 & ((~reg124) ?
                  (reg213[(4'h8):(2'h2)] ?
                      $unsigned(reg264) : reg258[(3'h7):(3'h6)]) : reg218[(4'hc):(2'h2)])));
              reg329 <= $unsigned($unsigned(reg280));
              reg330 <= {(((reg114[(4'hc):(3'h4)] ?
                              (-reg156) : {reg211, reg178, wire121}) ?
                          $signed($signed(reg329)) : $signed($signed(wire82))) ?
                      (reg136[(4'h8):(1'h1)] ~^ reg218[(5'h12):(3'h7)]) : ($unsigned((^reg157)) + (reg274[(1'h1):(1'h0)] ^~ {reg182,
                          reg321,
                          reg150}))),
                  $signed(($unsigned((~reg101)) == (~|$unsigned(wire81))))};
              reg331 = (-reg250);
              reg332 <= (~&$unsigned($signed($signed({reg136,
                  reg284,
                  reg321}))));
              reg333 = $signed($signed($signed((7'h4d))));
            end
          for (forvar334 = (1'h0); (forvar334 < (3'h5)); forvar334 = (forvar334 + (1'h1)))
            begin
              reg335 = $unsigned({reg250[(4'h8):(3'h4)],
                  ($signed(reg127) ^~ ((reg187 >>> reg105) <<< (!reg191)))});
              reg336 <= (~&reg218);
              reg337 = $signed(reg166);
            end
          for (forvar338 = (1'h0); (forvar338 < (3'h4)); forvar338 = (forvar338 + (1'h1)))
            begin
              reg339 <= ($unsigned($signed((&reg212[(1'h0):(1'h0)]))) ?
                  reg229 : (8'hbf));
            end
          for (forvar340 = (1'h0); (forvar340 < (3'h6)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 = reg260[(4'h9):(4'h8)];
              reg342 <= (~&(reg192 != $signed(((reg339 ? reg119 : reg178) ?
                  (reg216 ? reg122 : reg114) : (reg127 >= reg84)))));
              reg343 <= ($unsigned(((((7'h47) > reg311) < {reg293,
                  (8'ha5)}) != $signed((reg210 << reg139)))) <<< (reg212 ?
                  ((^(~reg329)) ?
                      (^reg215) : (|$signed(reg317))) : $signed((7'h49))));
            end
        end
      else
        begin
          for (forvar318 = (1'h0); (forvar318 < (2'h3)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg320 <= reg186;
              reg321 <= reg182[(4'hd):(4'h9)];
              reg323 = reg205[(1'h0):(1'h0)];
              reg325 = ($unsigned((~$unsigned(((7'h43) * reg206)))) ?
                  (!(~&{wire121,
                      (reg280 * wire233)})) : $unsigned(reg162[(3'h5):(3'h5)]));
            end
          reg326 = (($unsigned({$signed((8'hbe)), (wire82 ? reg288 : reg148)}) ?
                  ($unsigned(reg275) ?
                      reg337 : $unsigned($unsigned(reg313))) : (^~$unsigned(wire233))) ?
              forvar327 : (reg249 ?
                  $signed($signed(reg205[(3'h4):(3'h4)])) : $unsigned($signed({(7'h4b),
                      reg258}))));
        end
    end
  assign wire344 = (-{reg270[(3'h5):(2'h2)]});
  always
    @(posedge clk) begin
      for (forvar345 = (1'h0); (forvar345 < (3'h5)); forvar345 = (forvar345 + (1'h1)))
        begin
          if ($unsigned((8'hb7)))
            begin
              reg346 <= ((8'ha0) == $signed(reg219[(4'h8):(2'h3)]));
              reg347 <= (forvar345[(3'h4):(1'h1)] == (({forvar345} ?
                      $signed((reg330 ?
                          (7'h44) : reg156)) : (reg262[(4'h8):(1'h0)] <= reg270)) ?
                  reg157[(2'h2):(1'h0)] : reg293[(3'h4):(1'h0)]));
            end
          else
            begin
              reg348 = reg347[(4'hb):(1'h0)];
              reg349 = ((|{(-(reg87 ? (7'h4b) : reg92))}) ?
                  wire78 : $unsigned((((wire81 ?
                      reg317 : reg343) > ((7'h46) <= reg124)) || (|reg227))));
              reg350 = $unsigned(({reg349} < {($unsigned(reg349) ?
                      reg239[(4'hd):(4'hc)] : ((7'h56) ? reg119 : (8'ha4))),
                  reg279,
                  reg346[(2'h2):(1'h0)]}));
              reg351 = reg136[(3'h5):(1'h1)];
              reg352 <= reg213;
              reg353 <= $signed(reg351);
              reg354 <= $signed(($unsigned(reg174[(4'hc):(4'ha)]) >> (~&reg339[(5'h1d):(5'h1a)])));
            end
          reg355 <= reg219[(4'h9):(4'h9)];
          reg356 = $signed((reg105[(5'h15):(4'h8)] <= $signed((reg255[(3'h4):(2'h3)] ?
              reg227 : reg309[(5'h16):(3'h4)]))));
          if ({$unsigned(reg186), reg279[(1'h1):(1'h0)]})
            begin
              reg357 = reg286;
              reg358 = $signed(({reg288[(4'hd):(1'h0)]} ?
                  $unsigned(((reg330 < wire83) << wire344[(2'h2):(2'h2)])) : (reg293[(5'h14):(1'h0)] >>> reg262)));
              reg359 <= wire233;
              reg360 = ({reg97,
                      ((^(reg250 ? (7'h57) : reg329)) && $unsigned(reg329)),
                      wire79[(4'h8):(2'h3)]} ?
                  $signed((~&reg275[(3'h7):(3'h5)])) : $unsigned(reg182[(2'h3):(2'h2)]));
              reg361 <= ((8'hb5) << $unsigned($unsigned($unsigned(reg178[(4'hd):(4'hd)]))));
            end
          else
            begin
              reg357 = (|(($unsigned($signed(reg311)) ?
                  reg317[(3'h4):(2'h2)] : reg346) < $unsigned($signed(reg328))));
              reg358 = (~((~^reg125[(3'h7):(1'h0)]) | $signed((~|$unsigned(reg153)))));
              reg359 <= ((wire78 << {$signed((+reg258))}) * reg208[(4'ha):(1'h0)]);
              reg360 = (reg349[(3'h4):(1'h0)] ?
                  ((({reg125,
                      reg143} >>> reg260[(3'h4):(3'h4)]) - $signed(reg293)) ^~ $unsigned(reg128[(4'h8):(3'h6)])) : (reg224[(4'he):(2'h3)] >= ({$unsigned(reg224),
                      (reg356 ? reg353 : reg294),
                      $signed(reg313)} <<< (~(~|reg288)))));
              reg361 <= (reg332 && (^~(8'hbc)));
              reg362 <= $unsigned(reg96);
            end
          reg363 <= reg258[(4'ha):(4'h9)];
          for (forvar364 = (1'h0); (forvar364 < (3'h5)); forvar364 = (forvar364 + (1'h1)))
            begin
              reg365 = {(8'hbe)};
              reg366 = $unsigned(($unsigned($signed((reg157 >> reg97))) ?
                  {reg92[(5'h19):(5'h18)],
                      ((reg249 * reg291) <<< reg293[(5'h15):(4'h9)]),
                      ((reg275 != reg122) >= {reg157})} : reg281));
            end
          if ((7'h56))
            begin
              reg367 <= (((($unsigned(reg274) > $signed(reg355)) && {reg288[(4'he):(1'h0)]}) ?
                      reg352[(3'h6):(1'h0)] : (reg211 <<< (!reg142))) ?
                  reg191[(1'h1):(1'h0)] : {$signed((reg226[(5'h13):(3'h5)] << reg175[(3'h4):(2'h2)])),
                      ((|(+reg175)) ?
                          {(~^reg294),
                              ((8'hab) ?
                                  reg260 : reg84)} : ((reg219 >= reg353) & ((8'ha6) ?
                              reg87 : reg154))),
                      reg246});
              reg368 = reg293[(5'h13):(4'ha)];
              reg369 <= reg187;
              reg370 <= ((({(reg250 ? reg156 : reg270),
                      {reg95, reg291},
                      (wire266 ? reg270 : reg99)} ?
                  (!reg318[(1'h1):(1'h0)]) : ({reg281,
                      reg357} != reg254[(1'h0):(1'h0)])) << $signed($unsigned({reg175}))) ~^ $unsigned(reg357[(3'h5):(3'h4)]));
              reg371 <= ($unsigned((+(reg270[(1'h0):(1'h0)] ?
                  (&(7'h4c)) : {forvar345,
                      reg360,
                      (8'hbd)}))) == (+reg95[(2'h3):(1'h1)]));
              reg372 = reg206;
              reg373 = $unsigned(reg286[(4'h9):(2'h3)]);
            end
          else
            begin
              reg367 <= $signed($unsigned(((8'h9d) ?
                  (reg156[(4'hd):(1'h0)] ?
                      ((8'hba) >= reg361) : (reg373 * reg371)) : (reg346 ?
                      $signed(reg355) : (reg343 > (8'hb4))))));
              reg369 <= (8'haa);
              reg370 <= (|(reg236 << $unsigned((wire233 < (8'hbf)))));
            end
        end
      if ((~&(reg281[(3'h7):(1'h1)] ?
          (~&(reg320 ?
              $unsigned(reg361) : (!reg361))) : $unsigned(reg203[(3'h6):(2'h2)]))))
        begin
          reg374 = $unsigned(reg270);
          reg375 = (|$signed((|$unsigned((reg128 ? reg114 : reg275)))));
          for (forvar376 = (1'h0); (forvar376 < (2'h3)); forvar376 = (forvar376 + (1'h1)))
            begin
              reg377 = reg350;
              reg378 = reg167[(1'h1):(1'h1)];
              reg379 = (wire233 ^~ reg251);
            end
        end
      else
        begin
          for (forvar374 = (1'h0); (forvar374 < (2'h2)); forvar374 = (forvar374 + (1'h1)))
            begin
              reg376 <= $unsigned({$signed((8'ha9))});
              reg377 = {$signed(wire121[(5'h14):(4'ha)])};
              reg378 = ((reg377[(4'hc):(3'h6)] == reg213[(1'h0):(1'h0)]) ?
                  $signed(reg154[(3'h5):(3'h4)]) : ($unsigned((|reg374)) ^~ $unsigned(($unsigned(reg286) ?
                      $signed(reg191) : (~^reg288)))));
            end
          if (($unsigned(reg239) | (~|(|(reg182 ?
              $unsigned(forvar345) : (reg260 ? reg182 : reg352))))))
            begin
              reg379 = reg286[(2'h3):(2'h2)];
              reg380 <= reg288;
              reg381 <= (~^{reg351[(3'h7):(2'h3)]});
              reg382 <= $unsigned(reg354);
              reg383 <= $signed(((~|{(reg156 ?
                      reg250 : (8'hb0))}) < $signed($signed($signed(reg146)))));
            end
          else
            begin
              reg379 = ($unsigned({$unsigned(reg216[(2'h3):(2'h2)]),
                  ($signed(forvar345) | $unsigned(reg375)),
                  ($unsigned(reg268) != $signed((7'h4b)))}) - (+{$unsigned(reg320[(1'h0):(1'h0)]),
                  {$unsigned(reg365)}}));
            end
          reg384 = (!$signed(reg329));
          reg385 = {{$unsigned((-reg239)), $signed(reg317[(4'hf):(2'h3)])},
              reg182};
          if ((-reg127))
            begin
              reg386 = $unsigned(reg362);
              reg387 <= ($unsigned($unsigned({(reg264 - reg263),
                      {reg139, reg127, reg239}})) ?
                  {reg191[(5'h1e):(5'h14)],
                      (~&reg251[(4'hb):(3'h4)])} : (&(($signed(reg330) ?
                      (reg258 <<< reg249) : (&reg352)) ^ reg127[(2'h3):(1'h0)])));
              reg388 = (reg148[(1'h1):(1'h0)] ?
                  $signed((|($unsigned(forvar376) ?
                      (reg384 ?
                          reg192 : reg211) : (&reg134)))) : {$unsigned($signed((reg367 >>> reg328)))});
              reg389 = wire82;
              reg390 = ($unsigned((($signed(reg352) ?
                      (forvar364 <<< reg191) : ((7'h50) ?
                          reg99 : reg291)) && {reg227[(2'h2):(1'h0)],
                      $unsigned(reg351),
                      {reg208, reg348}})) ?
                  (reg95[(3'h6):(1'h1)] >> $signed(reg313[(1'h0):(1'h0)])) : reg363);
              reg391 = ((!reg279) << (((-wire78) ?
                      $signed((~^(7'h54))) : $unsigned((reg125 * reg348))) ?
                  (reg357[(1'h1):(1'h0)] >= {(wire81 ^~ (7'h46)),
                      (reg263 ? reg218 : reg120),
                      reg189[(4'hb):(3'h7)]}) : ((+reg128[(5'h19):(4'he)]) != $unsigned((~reg232)))));
            end
          else
            begin
              reg386 = $signed($signed((7'h47)));
              reg387 <= {(|(reg383[(3'h5):(3'h4)] || (~|$signed((8'hb3)))))};
              reg392 <= (reg381 ? $unsigned((+reg218)) : reg388);
              reg393 <= (&($signed($signed(reg213)) | ($signed((reg215 ?
                      reg380 : reg307)) ?
                  $unsigned(reg275) : reg124)));
              reg394 <= ($unsigned($unsigned((reg289 ~^ (^~reg329)))) ?
                  reg343[(4'hc):(4'hb)] : ((reg347[(3'h6):(3'h6)] > reg239[(3'h6):(3'h4)]) < $unsigned({wire79[(1'h0):(1'h0)]})));
              reg395 <= {$signed((reg351 <<< $unsigned((!reg384))))};
              reg396 <= reg318;
            end
        end
      reg397 = ($unsigned(wire344) & $unsigned(((-reg268) ?
          $signed(reg317[(3'h6):(3'h6)]) : reg392[(3'h4):(2'h3)])));
      if (reg280[(1'h0):(1'h0)])
        begin
          reg398 <= $signed($signed(reg227));
          for (forvar399 = (1'h0); (forvar399 < (2'h3)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg400 <= $unsigned(($unsigned($signed(reg380)) << reg313[(4'h8):(3'h6)]));
              reg401 = $unsigned(reg167[(3'h4):(3'h4)]);
              reg402 <= ({(((reg250 + (8'hb0)) ?
                          (reg215 ? reg361 : reg114) : (reg154 ?
                              reg384 : reg174)) ^~ ({reg376,
                          reg390} <<< ((8'hb3) ? reg216 : reg369))),
                      reg329,
                      (8'hb4)} ?
                  (($unsigned({reg366, reg258}) ?
                      reg369 : reg397[(5'h12):(2'h3)]) >>> reg347[(5'h15):(4'h9)]) : reg84[(5'h17):(4'hc)]);
              reg403 = reg203[(2'h2):(2'h2)];
              reg404 <= (reg218 >= reg378[(5'h1a):(5'h15)]);
              reg405 = (reg156 ?
                  reg241 : {($unsigned(((8'hb4) ? (7'h49) : reg149)) ?
                          reg359 : $signed($unsigned(reg142)))});
              reg406 <= {reg226, (^~reg187[(3'h7):(3'h7)])};
            end
        end
      else
        begin
          reg399 = reg203[(1'h1):(1'h0)];
          reg401 = (~&$unsigned(((-(8'had)) < ((reg216 - reg398) ?
              reg212 : (reg208 < (8'ha5))))));
        end
      if ($signed({$signed(($signed(reg128) * (|reg362))),
          $signed($unsigned($unsigned((8'ha0)))),
          ((~&$signed(reg114)) * reg393[(2'h2):(1'h0)])}))
        begin
          if ((reg148 ? reg92 : reg354))
            begin
              reg407 = reg359[(3'h6):(3'h6)];
              reg408 <= $unsigned(reg372[(3'h4):(3'h4)]);
              reg409 <= $signed((($signed((~reg148)) * ((reg348 ?
                          forvar399 : reg87) ?
                      {reg277, reg156, reg370} : (reg174 ? reg219 : reg88))) ?
                  $signed($signed((!(7'h52)))) : $signed($signed((reg264 << wire78)))));
              reg410 <= (reg357[(3'h7):(3'h4)] | $unsigned($signed(reg320)));
              reg411 = $unsigned($unsigned((^(+(wire121 ? reg356 : reg153)))));
              reg412 <= (^(wire78 ?
                  $unsigned($unsigned((reg205 ?
                      reg281 : reg386))) : (^$unsigned((reg324 < (7'h49))))));
            end
          else
            begin
              reg407 = $signed({$unsigned($signed((reg313 || reg358)))});
              reg408 <= (((+(((7'h42) ? reg353 : reg134) > {reg139,
                  reg372})) & (reg357 & $unsigned((~^wire265)))) || (&(|((|reg206) ?
                  $unsigned(reg313) : (^~reg227)))));
              reg409 <= $signed((reg400[(2'h2):(1'h0)] || (((!reg394) && reg401) <<< $unsigned((reg84 ?
                  reg206 : reg346)))));
              reg411 = reg354[(3'h4):(2'h2)];
              reg413 = (7'h49);
            end
          reg414 = (^~(&(reg142 ?
              reg249[(5'h11):(3'h7)] : reg88[(4'h8):(1'h0)])));
          reg415 = $unsigned(($unsigned(((!(8'h9e)) && $signed(reg85))) + $signed($signed((reg352 ?
              reg203 : (8'hbe))))));
          if ((reg275[(3'h4):(2'h3)] && ((~$unsigned((reg389 ?
              (8'hb0) : wire79))) != {$unsigned((reg127 ? (7'h4e) : reg148))})))
            begin
              reg416 = $unsigned({$unsigned(reg120),
                  $signed((&(8'ha9))),
                  $signed(reg232)});
              reg417 = $unsigned(((+$unsigned(reg246[(4'hb):(4'ha)])) ?
                  ((reg387 < (reg411 ~^ reg404)) << (~(reg236 ^ reg404))) : $signed($unsigned((reg374 > reg255)))));
              reg418 <= ((^~((8'hbe) ?
                  (^~(!reg150)) : ((reg149 - reg289) ?
                      (-forvar345) : $unsigned((8'hba))))) ^~ $unsigned($signed($signed(reg311))));
              reg419 <= {reg361[(4'hd):(4'hd)],
                  reg375[(3'h4):(2'h3)],
                  $unsigned(reg376[(5'h15):(4'hb)])};
              reg420 = forvar345[(3'h5):(3'h5)];
              reg421 <= (reg342[(3'h5):(3'h5)] ?
                  (({(~&reg420), (reg150 ~^ reg192)} ?
                          reg388[(5'h12):(2'h3)] : (reg363[(5'h10):(4'hd)] ?
                              reg213 : reg378[(4'he):(4'h8)])) ?
                      (($signed(reg239) != (reg415 ?
                          reg396 : reg387)) - ((reg293 > reg157) || reg241)) : $signed((^reg403))) : (~|{($unsigned(reg330) ?
                          reg416[(1'h1):(1'h1)] : $unsigned((7'h42))),
                      reg219,
                      (^~(reg349 ? reg373 : reg153))}));
            end
          else
            begin
              reg418 <= ((~^(^~reg146[(3'h5):(3'h5)])) ?
                  $unsigned($unsigned((~|((7'h4e) * reg85)))) : $signed((reg218[(4'hc):(1'h1)] ~^ (reg124[(2'h3):(1'h1)] ?
                      (reg128 | wire78) : {reg407, reg210}))));
              reg420 = (8'hac);
            end
        end
      else
        begin
          for (forvar407 = (1'h0); (forvar407 < (1'h0)); forvar407 = (forvar407 + (1'h1)))
            begin
              reg408 <= reg218[(3'h6):(1'h1)];
              reg409 <= (~^($signed({{reg402, reg162}}) ?
                  reg139 : (^~(~^reg241[(4'ha):(3'h6)]))));
              reg411 = ($unsigned(reg381[(1'h1):(1'h1)]) == ($unsigned((^~$signed(reg294))) >>> (~&((~reg239) ^ $signed(reg122)))));
              reg412 <= ($unsigned($unsigned($signed($signed(reg391)))) ?
                  (reg216[(1'h0):(1'h0)] ?
                      $signed($signed((~^reg311))) : reg361[(5'h11):(2'h3)]) : ((~^(reg336[(3'h7):(3'h4)] ?
                          reg343 : $unsigned(reg328))) ?
                      $signed(reg400) : (&($signed(reg356) - $signed(reg150)))));
              reg413 = reg182;
              reg418 <= {{(8'hbc),
                      reg167[(1'h1):(1'h0)],
                      ($signed(reg399) != (~^$unsigned((8'had))))},
                  reg354};
            end
          reg420 = ($signed(reg274[(4'hf):(4'hf)]) ?
              wire83[(5'h11):(3'h6)] : (7'h54));
          for (forvar421 = (1'h0); (forvar421 < (3'h5)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg422 <= $signed(reg380[(5'h1a):(4'hf)]);
              reg423 = $unsigned((|reg279[(1'h0):(1'h0)]));
              reg424 <= (~$signed($signed($signed({reg189}))));
              reg425 = $unsigned((~&(reg255 ~^ {(reg351 ? (8'hab) : (7'h58)),
                  reg395,
                  reg408})));
              reg426 <= (+{reg362[(1'h1):(1'h1)],
                  ((&(forvar421 ? reg361 : reg224)) >> reg369[(1'h1):(1'h0)]),
                  {{((7'h4d) ^~ reg374)}}});
            end
          reg427 <= ({{((wire265 ? wire83 : reg139) ? (~&reg401) : reg336)},
                  reg329[(5'h15):(2'h3)]} ?
              $signed($signed({(reg270 - reg142),
                  (reg85 < (7'h45)),
                  reg401})) : reg347);
          for (forvar428 = (1'h0); (forvar428 < (1'h0)); forvar428 = (forvar428 + (1'h1)))
            begin
              reg429 = (reg394[(2'h3):(2'h2)] >>> (((~^$unsigned(reg352)) & {$unsigned(reg349),
                      ((8'hac) ? reg385 : wire344)}) ?
                  reg311 : (reg97 ?
                      ((reg395 ?
                          forvar376 : reg427) ^~ reg210[(3'h5):(1'h1)]) : $unsigned((reg229 ?
                          reg377 : reg386)))));
              reg430 = reg134[(1'h0):(1'h0)];
              reg431 <= ((~^$signed(wire344)) ?
                  (reg328 ?
                      ({(8'had), reg157} ?
                          (-(reg361 ^~ reg157)) : $unsigned((reg397 ?
                              reg365 : reg367))) : reg249[(3'h4):(1'h0)]) : $signed(({reg311,
                      reg355,
                      (^(7'h46))} > wire83[(4'ha):(2'h3)])));
              reg432 = (8'ha8);
            end
        end
      if ((((reg313[(4'hc):(3'h7)] ?
          reg291[(1'h0):(1'h0)] : ($signed(reg408) ?
              {reg210,
                  (7'h4a),
                  reg406} : $unsigned(reg392))) < reg320[(1'h0):(1'h0)]) ^ reg124))
        begin
          for (forvar433 = (1'h0); (forvar433 < (2'h2)); forvar433 = (forvar433 + (1'h1)))
            begin
              reg434 <= (+($signed({reg95[(3'h5):(3'h5)], $signed(reg182)}) ?
                  ($unsigned((&(8'ha0))) ^~ wire80[(1'h1):(1'h1)]) : reg88));
              reg435 <= $unsigned(reg370);
              reg436 = ($unsigned({($unsigned((8'ha2)) ?
                      $signed(reg99) : reg401)}) == $unsigned($signed(reg429)));
            end
          for (forvar437 = (1'h0); (forvar437 < (1'h0)); forvar437 = (forvar437 + (1'h1)))
            begin
              reg438 <= $unsigned(reg105);
              reg439 = (8'hb0);
            end
        end
      else
        begin
          reg433 = ($signed({(reg324 ? (8'hb7) : reg307)}) ?
              (($unsigned($signed(reg408)) ?
                  {reg224,
                      (&forvar399)} : (^$unsigned((7'h4e)))) ^~ $unsigned((~&reg95[(3'h6):(3'h5)]))) : $signed((~^reg393)));
          reg434 <= reg260;
          if ({(~|reg402[(5'h10):(4'he)]),
              (&(forvar399 ? (^{reg255, (8'haa)}) : $unsigned(reg400))),
              ((~reg324) ?
                  {((reg285 ? forvar428 : wire265) ~^ (reg264 || reg332)),
                      (8'hbe)} : (reg189 & (!(reg289 >= (8'haa)))))})
            begin
              reg436 = reg409;
              reg437 <= {$signed((reg150[(1'h0):(1'h0)] != $signed((reg124 && reg381)))),
                  $signed($unsigned(reg251[(5'h11):(2'h3)])),
                  $signed(reg400[(2'h3):(1'h1)])};
              reg439 = (!$signed(reg154[(2'h2):(1'h0)]));
              reg440 <= (~&((~($signed(reg202) + $unsigned(reg397))) ?
                  {{(~^reg388)}} : (reg164 || reg390)));
            end
          else
            begin
              reg435 <= {reg320};
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed($unsigned(reg318[(3'h7):(3'h5)])))
        begin
          reg441 <= (~^(-({((7'h51) ? reg251 : reg128),
              reg167,
              $signed(reg329)} >= ($unsigned(reg115) & (+reg134)))));
          reg442 = $unsigned((-$unsigned(reg162[(2'h3):(2'h3)])));
          reg443 <= reg427[(4'ha):(1'h0)];
          if ((reg321[(2'h3):(1'h0)] + $unsigned(($signed((wire265 * reg270)) ?
              {$signed(reg153),
                  reg321[(2'h3):(2'h3)]} : reg362[(3'h5):(2'h3)]))))
            begin
              reg444 = {reg268[(1'h1):(1'h1)],
                  ((((&reg376) ?
                      reg330[(1'h0):(1'h0)] : reg226[(1'h1):(1'h0)]) ^ ((7'h51) ?
                      reg119[(5'h14):(3'h6)] : $unsigned(reg400))) + {(7'h4c),
                      reg410[(3'h6):(3'h4)]})};
              reg445 = $unsigned((|$unsigned(reg254)));
              reg446 <= $signed(reg270);
              reg447 = ($unsigned($unsigned(reg438[(2'h2):(1'h1)])) ^ $signed((~^$signed((reg216 ?
                  reg142 : reg255)))));
              reg448 <= (-(reg396 ?
                  $unsigned(($signed(reg205) <= wire344)) : $unsigned(reg354[(3'h6):(3'h4)])));
              reg449 <= $unsigned(reg336[(4'hd):(4'hd)]);
              reg450 = {$signed(((-$unsigned(reg422)) ?
                      ((reg119 ? reg409 : reg260) ^ (reg166 ?
                          reg355 : (8'hb7))) : reg394))};
            end
          else
            begin
              reg446 <= reg435;
              reg448 <= (~^$signed((reg354[(3'h6):(3'h6)] ?
                  (-(reg164 - reg307)) : (&(wire344 & reg236)))));
              reg450 = $signed({(~&((reg328 <= reg371) & {wire78,
                      reg361,
                      reg96})),
                  $signed($signed($signed(reg125))),
                  (8'hac)});
              reg451 <= (reg191 == reg434[(1'h0):(1'h0)]);
            end
          if ((8'h9e))
            begin
              reg452 = {$unsigned(reg189),
                  {$unsigned(reg254[(4'hd):(4'ha)]),
                      (wire121[(4'hc):(4'ha)] ?
                          $signed($signed(reg128)) : (8'ha5)),
                      {((reg298 ? reg143 : reg320) ?
                              (reg387 ? reg156 : (7'h46)) : {(8'hb6), reg174}),
                          reg359,
                          reg107}}};
              reg453 <= {($unsigned((reg329 ?
                      reg249 : (wire82 || reg178))) + (~|((~|reg246) & (~&reg400)))),
                  $unsigned((|$signed($signed(reg342))))};
              reg454 = (reg162 ?
                  {$unsigned($signed(reg219)),
                      (~(&(~|reg150))),
                      $unsigned(reg219)} : (({reg280,
                          (reg148 ? reg174 : reg451),
                          (reg284 ? reg410 : reg383)} ?
                      reg166[(2'h2):(1'h1)] : ((8'hbd) ?
                          (+reg362) : ((7'h4f) != (7'h56)))) >> ((~^$signed((8'hb2))) | (reg153 ?
                      {reg426} : (reg127 >> reg419)))));
              reg455 = {reg336,
                  $unsigned(((+(reg382 ?
                      reg409 : (8'hac))) == ($unsigned(reg101) != (reg434 ?
                      reg398 : reg263)))),
                  ($signed((~^(reg211 ^ reg277))) ~^ reg143[(4'h8):(3'h7)])};
              reg456 <= $signed((~^(~^reg321[(2'h3):(1'h1)])));
              reg457 = (&reg412);
            end
          else
            begin
              reg453 <= {$signed(reg178)};
              reg456 <= $signed(({reg154,
                      $unsigned(reg408),
                      $signed(reg241[(3'h5):(2'h3)])} ?
                  $unsigned(reg226) : $signed(reg452[(5'h1a):(4'hb)])));
              reg458 <= reg191;
              reg459 = $signed(reg236);
            end
          for (forvar460 = (1'h0); (forvar460 < (1'h1)); forvar460 = (forvar460 + (1'h1)))
            begin
              reg461 <= reg157[(1'h0):(1'h0)];
              reg462 <= $signed(reg307);
              reg463 <= $signed(wire266);
              reg464 <= $unsigned($unsigned($unsigned({$signed((7'h47))})));
              reg465 <= $unsigned((7'h56));
              reg466 <= reg88;
            end
        end
      else
        begin
          for (forvar441 = (1'h0); (forvar441 < (2'h2)); forvar441 = (forvar441 + (1'h1)))
            begin
              reg442 = reg167[(2'h2):(2'h2)];
              reg444 = ($unsigned(reg444[(5'h11):(4'hc)]) >> $unsigned(($unsigned((^(8'hbc))) ?
                  ($unsigned((8'ha8)) ?
                      (~|wire83) : (reg343 << reg107)) : reg298)));
              reg446 <= (reg449 ?
                  $unsigned($signed(reg309)) : $unsigned(((~&(wire233 & wire121)) < ($signed(reg294) ^ $signed(reg122)))));
              reg447 = reg127;
            end
          for (forvar448 = (1'h0); (forvar448 < (3'h4)); forvar448 = (forvar448 + (1'h1)))
            begin
              reg450 = (+$signed($signed(reg353)));
              reg451 <= (|(({(reg451 & reg427),
                      {reg192}} >>> (!(reg241 ~^ (7'h40)))) ?
                  ((|$signed(reg127)) ? reg210 : reg443) : {{(|reg453),
                          (7'h55),
                          (reg211 ? reg442 : reg275)},
                      $unsigned($signed(reg122)),
                      ($signed(reg418) ?
                          $unsigned(reg216) : reg285[(3'h4):(2'h3)])}));
              reg453 <= (reg206 == $signed((|((reg412 ? (8'hbf) : reg359) ?
                  reg450 : reg362[(4'h9):(3'h7)]))));
              reg454 = wire233;
            end
          for (forvar455 = (1'h0); (forvar455 < (3'h4)); forvar455 = (forvar455 + (1'h1)))
            begin
              reg457 = (~^reg313);
              reg458 <= $signed({((~^(reg263 ^ reg249)) ? reg442 : reg216)});
            end
          reg459 = (({reg453} * (((8'ha0) <= $unsigned(reg330)) ?
                  (reg454[(1'h1):(1'h0)] ?
                      reg462[(5'h15):(4'h9)] : (reg410 ?
                          reg438 : (8'ha0))) : ((reg260 << reg396) >>> {reg318,
                      reg452,
                      reg402}))) ?
              (+(reg437[(5'h14):(4'h9)] ^ {(reg270 > (7'h46)),
                  reg313,
                  (reg189 <<< reg241)})) : $signed(($signed((reg249 ?
                      reg146 : reg148)) ?
                  $unsigned((|reg408)) : (((7'h46) ? reg293 : reg139) ?
                      $signed(reg255) : (|(8'hac))))));
        end
    end
  assign wire467 = ((wire121 > {reg343[(3'h4):(2'h2)]}) ?
                       (reg134 || (((reg329 ? reg254 : (7'h41)) | {reg107,
                           (8'hbd)}) - $signed({reg346,
                           reg363}))) : reg321[(1'h1):(1'h1)]);
  assign wire468 = (~^{$signed($unsigned({reg381, wire233})),
                       $signed(wire266),
                       reg398});
  assign wire469 = reg127[(4'hd):(3'h6)];
  assign wire470 = $signed(reg258);
  assign wire471 = ((reg449[(2'h3):(2'h3)] ?
                           $unsigned(({reg322, reg241, reg134} ?
                               ((8'h9e) | reg369) : (8'ha7))) : ((^~$signed(reg187)) ?
                               {$signed((8'ha4)),
                                   (reg246 || reg322),
                                   (reg252 != reg139)} : ((!reg264) ?
                                   ((7'h40) <= reg270) : ((8'hb1) | reg260)))) ?
                       reg258 : ((~(8'ha7)) ?
                           $signed((-(^~reg440))) : (($signed(reg189) && (reg174 > (7'h47))) <<< $signed({reg342}))));
  always
    @(posedge clk) begin
      for (forvar472 = (1'h0); (forvar472 < (1'h1)); forvar472 = (forvar472 + (1'h1)))
        begin
          reg473 <= reg270;
          if ($signed(reg317[(4'h8):(2'h3)]))
            begin
              reg474 = ($unsigned((!reg167)) ?
                  wire469[(3'h4):(1'h1)] : $unsigned($unsigned($unsigned($signed(reg134)))));
              reg475 = (^~wire344[(3'h4):(2'h3)]);
              reg476 <= (($unsigned(($signed(reg288) ?
                      {reg149} : wire83[(4'ha):(2'h3)])) | reg466[(3'h6):(1'h0)]) ?
                  reg149 : $unsigned(reg320[(1'h1):(1'h0)]));
              reg477 <= reg213[(4'hf):(4'he)];
            end
          else
            begin
              reg476 <= reg97[(1'h1):(1'h1)];
              reg478 = (8'h9d);
            end
          reg479 = (~&reg291);
          reg480 = $unsigned({($signed(reg330) ?
                  reg150[(2'h2):(1'h1)] : ($unsigned((8'ha6)) ^ (~&reg473))),
              reg96[(3'h6):(3'h4)]});
          reg481 <= wire78[(3'h7):(3'h4)];
          reg482 = reg114;
          reg483 <= reg477[(2'h3):(1'h0)];
        end
      for (forvar484 = (1'h0); (forvar484 < (3'h4)); forvar484 = (forvar484 + (1'h1)))
        begin
          reg485 = {$signed($unsigned(($signed(reg462) >> (reg284 <= reg218)))),
              $signed($unsigned(reg424[(4'hb):(4'h8)]))};
          reg486 <= reg361;
          for (forvar487 = (1'h0); (forvar487 < (1'h1)); forvar487 = (forvar487 + (1'h1)))
            begin
              reg488 = $signed($signed((~reg434)));
              reg489 = {(((~&$signed(reg258)) + $signed($signed(wire78))) ?
                      $unsigned($signed($unsigned(reg298))) : reg352[(5'h11):(4'hd)]),
                  ($signed({{(8'hbf), reg120},
                      $unsigned(reg146)}) && (~^(+{(8'haf), reg393})))};
              reg490 = (~&((&reg157[(3'h4):(1'h1)]) ?
                  {reg157,
                      ((reg96 >= (8'hb6)) <<< $unsigned(reg239)),
                      wire81} : reg419));
            end
          for (forvar491 = (1'h0); (forvar491 < (1'h1)); forvar491 = (forvar491 + (1'h1)))
            begin
              reg492 <= $unsigned((reg409[(2'h3):(1'h1)] ?
                  $signed(reg394) : ((~reg250) ?
                      reg119[(5'h19):(4'he)] : ({reg392, reg150} ?
                          (reg435 ? reg298 : reg371) : {reg410,
                              reg166,
                              reg241}))));
              reg493 <= $unsigned($signed(($unsigned(reg480[(3'h5):(2'h3)]) ?
                  $unsigned($unsigned((7'h4e))) : (reg419 < (reg367 && reg346)))));
              reg494 <= reg182;
              reg495 = reg434[(4'h9):(3'h6)];
              reg496 <= (($signed({(+reg96), $unsigned(reg219), reg456}) ?
                      (7'h41) : reg270[(2'h2):(2'h2)]) ?
                  (8'hba) : $signed((|{(reg120 ? wire467 : reg318)})));
            end
        end
      for (forvar497 = (1'h0); (forvar497 < (1'h1)); forvar497 = (forvar497 + (1'h1)))
        begin
          if (((reg321 > reg480[(2'h2):(1'h0)]) && reg149))
            begin
              reg498 = $signed(reg494[(3'h5):(2'h2)]);
              reg499 <= wire471;
              reg500 = reg202;
              reg501 = (8'h9c);
              reg502 <= (8'hb3);
              reg503 = (^reg387[(5'h15):(3'h7)]);
            end
          else
            begin
              reg499 <= reg313[(2'h3):(2'h2)];
              reg502 <= reg329[(5'h1e):(5'h13)];
              reg504 <= reg438[(2'h2):(1'h0)];
            end
          reg505 <= $signed(wire470);
          reg506 <= (8'ha0);
          for (forvar507 = (1'h0); (forvar507 < (3'h5)); forvar507 = (forvar507 + (1'h1)))
            begin
              reg508 = $signed(reg404[(2'h3):(1'h0)]);
              reg509 = reg424[(4'h8):(3'h6)];
            end
          reg510 <= reg246[(2'h2):(2'h2)];
        end
    end
  assign wire511 = ($unsigned((+$signed(reg355))) >> (wire121 || {reg321,
                       wire78[(4'hb):(3'h7)]}));
  always
    @(posedge clk) begin
      reg512 = {{(reg150[(2'h3):(1'h0)] & wire470[(4'hc):(4'h8)]),
              (+(!(wire82 ? (8'haa) : (8'h9f)))),
              wire78[(4'h9):(4'h8)]},
          $unsigned(reg437[(5'h1f):(5'h13)])};
      reg513 <= {(reg322[(2'h3):(1'h1)] >> (~(+(reg270 ? reg275 : (8'hb5))))),
          wire80[(5'h11):(5'h10)],
          $unsigned($signed(reg448[(4'hc):(2'h3)]))};
      for (forvar514 = (1'h0); (forvar514 < (2'h3)); forvar514 = (forvar514 + (1'h1)))
        begin
          reg515 = $unsigned($unsigned(({(reg477 ^~ (7'h41)),
              reg212,
              reg139[(2'h3):(1'h1)]} - ($unsigned(reg343) ?
              $signed(reg275) : (reg227 == reg355)))));
          if (reg441[(2'h2):(1'h0)])
            begin
              reg516 <= reg355;
              reg517 <= ($unsigned(($signed($signed(wire81)) ^~ reg192)) ?
                  ($unsigned($signed((reg453 ?
                      (7'h52) : (7'h44)))) <= reg84[(5'h16):(5'h15)]) : reg505);
            end
          else
            begin
              reg518 = (reg95[(1'h1):(1'h1)] ^ $unsigned({(-(reg513 ?
                      (8'haf) : reg499)),
                  $signed({reg216, reg456}),
                  reg309}));
              reg519 = {$signed(((((7'h4a) ? reg466 : reg517) ?
                          reg382[(4'hd):(4'hb)] : (reg289 ^~ reg419)) ?
                      $unsigned($unsigned(reg254)) : ({(8'hb6),
                              reg451,
                              reg434} ?
                          reg101[(2'h3):(1'h0)] : wire511[(4'ha):(2'h2)]))),
                  (^{{$unsigned(reg189), reg178},
                      ($signed(reg120) != (~&reg274))})};
              reg520 = $unsigned(reg449);
            end
          reg521 <= (reg394 != $unsigned((|reg264)));
        end
      for (forvar522 = (1'h0); (forvar522 < (2'h3)); forvar522 = (forvar522 + (1'h1)))
        begin
          reg523 = ($unsigned((forvar522 ?
                  reg262 : $unsigned((reg87 ~^ reg361)))) ?
              $signed(($signed(reg330) >> $signed($unsigned(reg150)))) : (($signed({(8'haa),
                  reg275,
                  reg506}) + (reg250 ~^ $signed(reg458))) || ((|$signed(wire266)) ?
                  (reg435[(4'hf):(2'h3)] ?
                      (reg178 ?
                          reg332 : reg396) : $signed(reg203)) : $signed($signed(reg499)))));
          reg524 = (((($signed(reg404) ? $unsigned(reg513) : $signed((8'h9e))) ?
                  $signed((reg431 ? reg252 : reg406)) : {$signed(reg150),
                      (|reg260)}) - $unsigned($signed((reg150 <= reg252)))) ?
              reg449[(4'he):(4'hd)] : (!(~|({reg139, reg215, reg216} >> {reg362,
                  reg263}))));
        end
    end
  assign wire525 = ((!$unsigned((+reg370))) ?
                       {($unsigned($signed(reg241)) != ($unsigned(reg120) <= (reg400 | reg521))),
                           (|($unsigned(reg254) ?
                               reg521[(4'hc):(3'h6)] : (8'hbc)))} : ((($signed(wire344) ^ reg483) ?
                               wire80[(1'h1):(1'h1)] : (^~reg404[(4'ha):(2'h3)])) ?
                           $signed({$signed(reg336)}) : {(&$signed(reg317))}));
  always
    @(posedge clk) begin
      for (forvar526 = (1'h0); (forvar526 < (3'h6)); forvar526 = (forvar526 + (1'h1)))
        begin
          if (reg517[(1'h1):(1'h1)])
            begin
              reg527 = reg483[(2'h2):(1'h0)];
              reg528 <= $signed($signed($unsigned(((reg182 + reg227) ?
                  (reg451 ? reg343 : reg521) : reg294))));
              reg529 = ($unsigned((($signed(reg149) ?
                      reg124[(2'h2):(2'h2)] : {(7'h4e)}) << $unsigned(reg502))) ?
                  ((7'h53) << (~$signed(wire78))) : reg115);
            end
          else
            begin
              reg528 <= $unsigned($signed(($signed($signed(reg187)) ~^ (|{reg309}))));
              reg529 = reg288;
              reg530 = $signed((^~(({reg167, reg205, (8'ha2)} ?
                  $signed((7'h54)) : ((8'h9e) ?
                      reg462 : reg97)) != $unsigned(reg492[(1'h1):(1'h1)]))));
            end
          for (forvar531 = (1'h0); (forvar531 < (1'h0)); forvar531 = (forvar531 + (1'h1)))
            begin
              reg532 <= ((-((^~(reg275 >= reg322)) >> $unsigned($unsigned(reg270)))) ?
                  (7'h43) : $unsigned(reg128[(5'h12):(5'h10)]));
              reg533 <= reg473;
              reg534 = (!$signed($signed((!{reg380, reg210, reg354}))));
              reg535 <= reg394;
            end
          if ($unsigned(((|((&(8'ha2)) ?
              (~(8'hb0)) : (!reg369))) <= $unsigned($signed((reg258 ?
              reg262 : reg383))))))
            begin
              reg536 <= $unsigned(reg270);
              reg537 <= (reg115 - {((~&$unsigned(reg284)) ?
                      $signed(((8'hb7) ?
                          reg328 : reg157)) : ((reg492 == reg419) > reg499)),
                  {$signed($unsigned(reg210))},
                  $unsigned(($unsigned((7'h57)) ?
                      {(8'hae), reg418} : reg210[(2'h2):(2'h2)]))});
              reg538 <= ($signed(($unsigned((~reg451)) + reg402)) ?
                  (($unsigned((!wire470)) ?
                          (reg174 && (reg157 >>> reg354)) : $unsigned((wire467 ?
                              reg371 : (7'h40)))) ?
                      $unsigned((+$unsigned((7'h41)))) : (($unsigned(reg268) ?
                              (reg504 ?
                                  reg127 : reg529) : reg87[(4'h9):(2'h3)]) ?
                          reg154[(4'h8):(2'h3)] : (8'ha9))) : reg431[(2'h3):(2'h3)]);
              reg539 = $unsigned(((^~$signed((reg174 ? reg434 : reg164))) ?
                  (~$signed({(8'haa)})) : reg352));
              reg540 = reg529[(2'h3):(1'h1)];
              reg541 = $signed(($signed(reg449) == (reg317 ?
                  $unsigned($signed(reg268)) : reg281[(2'h2):(1'h1)])));
              reg542 = $unsigned(reg189);
            end
          else
            begin
              reg539 = ($unsigned($unsigned((reg212 ?
                      (-reg346) : $signed(wire265)))) ?
                  (($unsigned({wire80, reg394}) ?
                          (|reg142[(1'h0):(1'h0)]) : reg205) ?
                      reg506[(5'h1a):(5'h16)] : $signed((reg537[(5'h16):(3'h7)] ~^ (~|reg540)))) : $signed((reg203[(3'h7):(1'h0)] ?
                      $unsigned((reg215 - reg381)) : $unsigned((^~reg187)))));
            end
          for (forvar543 = (1'h0); (forvar543 < (1'h1)); forvar543 = (forvar543 + (1'h1)))
            begin
              reg544 <= $signed(($unsigned($unsigned(reg216)) ?
                  $unsigned($unsigned({reg354, reg361})) : (7'h4e)));
              reg545 <= ((reg504[(2'h3):(1'h1)] != ((wire82 ?
                      wire470[(4'h8):(1'h1)] : reg441) - reg530)) ?
                  {(|{(reg537 > (8'hba)), $signed(reg154), (~^reg293)}),
                      $unsigned((((7'h44) >>> (8'haf)) ?
                          (reg422 + reg317) : (reg437 > reg164))),
                      reg84[(1'h0):(1'h0)]} : $unsigned(reg250[(4'h8):(2'h3)]));
              reg546 <= (|(8'hb7));
              reg547 <= $unsigned(((wire525[(2'h2):(1'h0)] ?
                  ($signed(reg435) & (reg510 ~^ reg410)) : ((reg251 ?
                          reg255 : reg154) ?
                      ((8'h9d) > reg329) : $signed((8'hb3)))) | (($unsigned(reg463) <= {reg92,
                  (8'h9c),
                  reg449}) ^ (-reg506[(1'h0):(1'h0)]))));
              reg548 = reg359;
            end
        end
      reg549 <= ((&reg229) ? reg539 : (wire80[(4'ha):(2'h2)] == reg251));
      for (forvar550 = (1'h0); (forvar550 < (3'h4)); forvar550 = (forvar550 + (1'h1)))
        begin
          for (forvar551 = (1'h0); (forvar551 < (3'h4)); forvar551 = (forvar551 + (1'h1)))
            begin
              reg552 <= (reg499 ?
                  $signed((~&($signed(reg263) ^~ reg387))) : ({$unsigned({reg418}),
                          (-(reg186 && reg533)),
                          $signed((-reg285))} ?
                      (reg418 ?
                          {(reg342 ? wire511 : (7'h49)),
                              (wire470 ?
                                  reg437 : reg339)} : reg232[(4'he):(1'h0)]) : ($signed($unsigned(wire80)) > $unsigned(wire83))));
              reg553 <= (^$unsigned(reg254));
              reg554 = reg213[(4'hb):(4'h8)];
            end
          reg555 <= $signed(reg548[(4'ha):(3'h7)]);
          if ((($signed($unsigned($unsigned(reg281))) ?
              $signed($unsigned(reg249)) : reg530) | ($signed({(reg426 - reg409),
              (!wire79),
              (-forvar551)}) ~^ reg481)))
            begin
              reg556 <= (reg548 ^~ reg435[(4'hf):(4'hb)]);
              reg557 <= $unsigned(((8'hb7) ?
                  reg537 : ($unsigned($unsigned(reg232)) != ((reg380 <= reg538) * (!reg134)))));
              reg558 <= $signed($unsigned(reg270));
              reg559 = ((({(reg343 && reg421),
                      (~|reg542),
                      (reg419 ?
                          (7'h52) : reg92)} >= wire471[(4'ha):(4'ha)]) || reg434[(4'hb):(4'h9)]) ?
                  $unsigned(($unsigned($unsigned(reg291)) ?
                      $signed(reg232[(1'h0):(1'h0)]) : {(8'ha6),
                          {reg191, reg418},
                          $unsigned(reg262)})) : {$unsigned($signed((+reg496))),
                      (~&reg437)});
            end
          else
            begin
              reg556 <= ($unsigned($unsigned($unsigned((^~reg206)))) ?
                  {$unsigned((reg254[(4'hc):(1'h0)] >= (-(8'hb1))))} : (reg371[(2'h2):(1'h1)] >= $signed(reg392[(3'h4):(2'h2)])));
            end
          reg560 = $signed((({reg289[(1'h1):(1'h0)]} - $signed(reg125)) ^ ((8'ha8) ?
              (reg435[(4'hf):(4'hd)] || reg506) : (+$unsigned(reg277)))));
          if ($signed((^(!$unsigned({(7'h42)})))))
            begin
              reg561 = {$signed(($unsigned({reg343,
                      reg293}) > reg318[(5'h13):(3'h6)])),
                  reg175[(2'h2):(1'h1)]};
            end
          else
            begin
              reg562 <= (reg339[(5'h17):(2'h3)] ?
                  ({(reg381[(3'h7):(1'h1)] & $signed(reg156)),
                      reg88[(3'h6):(3'h5)]} || (reg307[(1'h0):(1'h0)] ?
                      reg120 : (~reg453[(3'h5):(2'h3)]))) : {reg461,
                      {reg453, reg546[(2'h2):(1'h1)]},
                      reg249[(4'ha):(1'h1)]});
              reg563 = ($signed($signed(((|reg167) ?
                  (&(7'h56)) : reg343[(4'hf):(4'hd)]))) | wire80);
              reg564 = (({({reg332, reg367} ?
                      $signed(reg320) : reg426[(1'h1):(1'h0)]),
                  (7'h46),
                  reg535[(5'h19):(5'h11)]} << (8'ha1)) | (^{reg311,
                  (((7'h40) - reg494) > reg547[(1'h1):(1'h1)])}));
              reg565 <= ((reg260 ?
                      {$signed($signed(reg535)),
                          reg481,
                          reg398[(3'h7):(1'h1)]} : (~|wire344[(1'h1):(1'h0)])) ?
                  $unsigned(($unsigned((^(7'h46))) ~^ $unsigned(reg535[(5'h16):(4'h9)]))) : $signed(reg182[(2'h3):(2'h3)]));
              reg566 <= $unsigned((((~^((8'hb4) == reg191)) - wire80) <<< reg324[(5'h18):(5'h15)]));
              reg567 <= (-(7'h44));
            end
          if ($unsigned(reg355[(3'h7):(2'h3)]))
            begin
              reg568 = {($signed(($signed(reg557) ?
                      {reg492,
                          reg541,
                          (8'haf)} : reg412[(3'h5):(2'h2)])) < $unsigned(reg128)),
                  ({$signed(reg532[(5'h14):(2'h3)])} ?
                      reg215[(2'h2):(2'h2)] : ($unsigned(wire468[(4'h8):(1'h0)]) ?
                          ($signed((7'h4b)) - (reg307 < wire525)) : $unsigned(reg382))),
                  reg88[(1'h1):(1'h1)]};
            end
          else
            begin
              reg568 = $signed((reg246[(1'h1):(1'h1)] ?
                  (~(forvar550[(1'h0):(1'h0)] && (reg361 << reg150))) : reg192[(3'h5):(1'h1)]));
              reg569 = reg293[(3'h4):(1'h1)];
              reg570 = reg559;
              reg571 = ((~&$unsigned((8'hbf))) ?
                  {reg370,
                      reg453[(4'hb):(3'h4)]} : $signed($unsigned({(7'h47)})));
              reg572 = (|$unsigned((((reg224 ^ (8'hb0)) ?
                  (reg298 == (7'h45)) : wire121) + $unsigned((reg408 * reg438)))));
              reg573 = {reg164[(5'h1d):(5'h14)],
                  ((|(~|reg263)) ?
                      (reg354 ?
                          (^$unsigned(reg437)) : reg398[(3'h4):(1'h0)]) : reg167[(1'h1):(1'h0)])};
              reg574 <= (7'h51);
            end
          if ({$unsigned((&reg208)),
              reg175[(2'h2):(1'h1)],
              $signed($unsigned(reg318))})
            begin
              reg575 = reg473;
              reg576 = reg355[(4'he):(3'h5)];
              reg577 <= reg548[(4'h9):(3'h5)];
              reg578 = reg542[(4'hb):(4'h8)];
              reg579 = (^($unsigned($signed((-(7'h4a)))) ^~ ((|$unsigned(reg174)) <<< ($unsigned(reg264) - (|reg227)))));
              reg580 <= $signed((reg87 ^ reg419[(2'h3):(1'h1)]));
              reg581 <= $signed(((^$unsigned($signed((8'had)))) >>> $signed($signed($unsigned(reg127)))));
            end
          else
            begin
              reg575 = (reg167[(1'h0):(1'h0)] >>> $unsigned(((((7'h57) >>> reg570) ^ wire467[(3'h4):(1'h1)]) ~^ $unsigned($unsigned(reg362)))));
              reg576 = (reg441 ^~ ((^~reg285) ^ (~&$unsigned({(7'h57)}))));
              reg577 <= reg427[(1'h0):(1'h0)];
              reg578 = ($signed((((reg275 >>> reg567) ? forvar551 : wire81) ?
                  (~reg566[(3'h6):(3'h4)]) : (8'hbd))) > reg381[(1'h0):(1'h0)]);
              reg580 <= ($unsigned(reg124) ?
                  (reg506[(3'h6):(1'h1)] ?
                      {$unsigned((7'h4d)),
                          $signed((reg547 ^ wire233)),
                          reg313[(4'ha):(4'h9)]} : $signed(((forvar550 ?
                          reg309 : (8'hac)) << (reg532 ?
                          reg418 : (8'hbe))))) : ((~&reg328) ?
                      (&reg164[(4'h8):(1'h1)]) : (reg438 ?
                          $signed((reg434 ? reg560 : reg410)) : (~&((8'h9e) ?
                              reg219 : wire467)))));
              reg582 = reg465[(3'h7):(3'h6)];
            end
        end
      reg583 <= reg264;
      if ((reg434 ?
          $unsigned((reg274 ~^ $signed($unsigned(reg382)))) : ({(reg120 * reg380[(5'h13):(5'h12)]),
                  reg572} ?
              (reg280[(1'h1):(1'h1)] ?
                  ((reg376 ?
                      reg398 : reg362) > $unsigned(reg219)) : reg127) : (reg232[(4'hd):(4'hc)] <<< reg367[(3'h4):(1'h0)]))))
        begin
          reg584 = (!(-reg577[(2'h3):(1'h1)]));
        end
      else
        begin
          for (forvar584 = (1'h0); (forvar584 < (1'h1)); forvar584 = (forvar584 + (1'h1)))
            begin
              reg585 <= reg189[(4'he):(4'hb)];
            end
          for (forvar586 = (1'h0); (forvar586 < (3'h6)); forvar586 = (forvar586 + (1'h1)))
            begin
              reg587 = $signed($unsigned(reg494[(4'h9):(3'h6)]));
              reg588 <= $unsigned(((((reg435 || reg208) >>> reg87) ^ reg206) ?
                  reg250[(4'ha):(4'ha)] : ({$unsigned(forvar584)} ?
                      wire266 : ({reg268, reg219, reg279} ?
                          wire78 : (|reg120)))));
              reg589 = {(reg167 ?
                      ($signed((reg251 != (8'hb6))) ?
                          $unsigned((wire344 ?
                              (7'h44) : (7'h50))) : $signed((~|reg328))) : reg186)};
            end
          reg590 <= $unsigned(({(8'ha5),
                  ((reg410 <<< reg150) ?
                      reg202[(5'h15):(2'h3)] : $unsigned(reg202)),
                  $signed((reg336 ? reg226 : reg557))} ?
              $signed(wire82) : reg277[(3'h5):(1'h0)]));
          for (forvar591 = (1'h0); (forvar591 < (3'h5)); forvar591 = (forvar591 + (1'h1)))
            begin
              reg592 = reg421[(2'h3):(2'h2)];
              reg593 = ((8'hac) ?
                  ((~({reg406} ?
                      $signed(reg210) : (reg587 & reg453))) & ($unsigned((reg255 ?
                      reg422 : reg446)) > reg275[(4'h8):(4'h8)])) : reg533[(2'h3):(2'h3)]);
              reg594 <= $signed(($signed((reg545[(1'h1):(1'h0)] ?
                      (reg162 ? reg461 : reg182) : reg362)) ?
                  {($signed(forvar584) >> (&reg464))} : ($unsigned($signed(reg313)) ?
                      (^~reg592) : (~|(reg483 <<< (7'h44))))));
              reg595 <= reg107;
              reg596 <= (reg229[(3'h4):(1'h1)] ?
                  $signed(reg541[(3'h6):(1'h0)]) : ((wire83[(2'h3):(2'h2)] > $unsigned($unsigned(reg254))) * (^(reg561 ?
                      $unsigned(reg584) : $signed(reg329)))));
            end
          for (forvar597 = (1'h0); (forvar597 < (3'h4)); forvar597 = (forvar597 + (1'h1)))
            begin
              reg598 = reg483;
              reg599 = $signed(reg492);
              reg600 <= reg431;
              reg601 = $signed($signed(($unsigned((reg552 ^ reg175)) << reg309)));
              reg602 = (((((reg205 * reg595) || (reg538 >> reg572)) & ((reg203 >= reg205) == (reg486 ?
                  reg187 : reg527))) == ($signed(reg143) ?
                  {reg97[(1'h1):(1'h0)],
                      reg595[(4'hb):(3'h5)],
                      (reg208 ~^ wire467)} : ((&wire469) || $unsigned(reg202)))) - (&$signed((reg336[(4'ha):(2'h3)] * ((8'hbd) << reg125)))));
              reg603 = (reg218 ~^ (^$unsigned(($signed(reg321) ?
                  $signed(reg441) : $signed(reg367)))));
            end
          reg604 <= ({$unsigned(reg426),
              $signed(((reg596 - wire469) ^ reg534[(4'hf):(4'h9)]))} | reg410[(3'h5):(3'h5)]);
          for (forvar605 = (1'h0); (forvar605 < (1'h1)); forvar605 = (forvar605 + (1'h1)))
            begin
              reg606 = reg294[(2'h3):(2'h3)];
              reg607 <= $signed(reg156);
              reg608 <= ((reg122 ~^ ($signed({reg309, reg566, reg202}) ?
                      ($signed(reg361) ?
                          $signed(reg578) : wire469[(4'h9):(2'h2)]) : (reg587[(2'h2):(2'h2)] ?
                          (~|reg441) : (reg328 && reg211)))) ?
                  reg481 : ((~$unsigned(reg548[(1'h0):(1'h0)])) ?
                      (!reg595[(3'h5):(3'h4)]) : (8'h9f)));
              reg609 <= {$unsigned($signed(reg280))};
              reg610 = (~|$signed(((reg232[(4'hb):(1'h0)] ^~ reg496[(4'ha):(2'h3)]) < $unsigned(reg189))));
            end
        end
      for (forvar611 = (1'h0); (forvar611 < (1'h0)); forvar611 = (forvar611 + (1'h1)))
        begin
          for (forvar612 = (1'h0); (forvar612 < (1'h0)); forvar612 = (forvar612 + (1'h1)))
            begin
              reg613 = $signed(($signed($signed($signed(reg424))) | (+$unsigned(wire511[(4'h9):(3'h4)]))));
              reg614 <= (^((-$signed($unsigned(reg293))) ?
                  (reg298[(4'hd):(1'h1)] >> (|reg530[(4'hd):(2'h3)])) : $signed(reg456)));
              reg615 = (+$signed(($unsigned($signed(reg219)) ?
                  $unsigned((!(8'hae))) : $signed($signed(reg451)))));
              reg616 <= {(~$signed($signed({(8'ha1), reg216}))),
                  reg359[(3'h6):(3'h6)],
                  (7'h54)};
            end
        end
    end
  assign wire617 = (&$unsigned((~&$unsigned($unsigned(reg502)))));
endmodule