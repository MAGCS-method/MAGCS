(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h9ee):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire3;
  input wire [(5'h10):(1'h0)] wire2;
  input wire signed [(5'h11):(1'h0)] wire1;
  input wire signed [(5'h18):(1'h0)] wire0;
  wire [(5'h13):(1'h0)] wire1769;
  wire signed [(5'h15):(1'h0)] wire1707;
  wire signed [(4'h9):(1'h0)] wire1631;
  wire [(5'h10):(1'h0)] wire337;
  wire signed [(5'h10):(1'h0)] wire24;
  wire [(5'h18):(1'h0)] wire1690;
  wire signed [(5'h11):(1'h0)] wire1691;
  wire [(3'h5):(1'h0)] wire1693;
  wire signed [(4'he):(1'h0)] wire1694;
  reg signed [(5'h18):(1'h0)] reg1783 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1781 = (1'h0);
  reg [(5'h16):(1'h0)] reg1779 = (1'h0);
  reg [(3'h5):(1'h0)] reg1778 = (1'h0);
  reg [(4'ha):(1'h0)] reg1774 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1773 = (1'h0);
  reg [(4'hf):(1'h0)] reg1770 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1766 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1764 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1761 = (1'h0);
  reg [(3'h6):(1'h0)] reg1760 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1759 = (1'h0);
  reg [(5'h13):(1'h0)] reg1757 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1756 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1755 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1751 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1750 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1748 = (1'h0);
  reg [(4'hd):(1'h0)] reg1747 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1744 = (1'h0);
  reg [(3'h7):(1'h0)] reg1743 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1742 = (1'h0);
  reg [(4'hd):(1'h0)] reg1738 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1736 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1731 = (1'h0);
  reg [(5'h15):(1'h0)] reg1730 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1729 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1728 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1726 = (1'h0);
  reg [(4'hb):(1'h0)] reg1725 = (1'h0);
  reg [(4'h8):(1'h0)] reg1720 = (1'h0);
  reg [(5'h18):(1'h0)] reg1718 = (1'h0);
  reg [(2'h2):(1'h0)] reg1716 = (1'h0);
  reg [(5'h16):(1'h0)] reg1714 = (1'h0);
  reg [(4'h9):(1'h0)] reg1704 = (1'h0);
  reg [(5'h10):(1'h0)] reg1703 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1698 = (1'h0);
  reg [(4'he):(1'h0)] reg1701 = (1'h0);
  reg [(5'h14):(1'h0)] reg1699 = (1'h0);
  reg [(4'hd):(1'h0)] reg1697 = (1'h0);
  reg signed [(4'he):(1'h0)] reg356 = (1'h0);
  reg [(3'h4):(1'h0)] reg353 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg350 = (1'h0);
  reg [(5'h14):(1'h0)] reg349 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg347 = (1'h0);
  reg signed [(4'he):(1'h0)] reg344 = (1'h0);
  reg [(5'h15):(1'h0)] reg340 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg21 = (1'h0);
  reg [(5'h13):(1'h0)] reg18 = (1'h0);
  reg [(5'h11):(1'h0)] reg15 = (1'h0);
  reg [(2'h3):(1'h0)] reg12 = (1'h0);
  reg [(2'h2):(1'h0)] reg5 = (1'h0);
  reg [(5'h18):(1'h0)] reg1633 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1636 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1637 = (1'h0);
  reg [(5'h11):(1'h0)] reg1640 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1641 = (1'h0);
  reg [(5'h10):(1'h0)] reg1642 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1647 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1649 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1654 = (1'h0);
  reg [(3'h5):(1'h0)] reg1657 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1658 = (1'h0);
  reg [(4'hd):(1'h0)] reg1655 = (1'h0);
  reg [(5'h10):(1'h0)] reg1661 = (1'h0);
  reg [(4'h8):(1'h0)] reg1662 = (1'h0);
  reg [(4'he):(1'h0)] reg1663 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1665 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1667 = (1'h0);
  reg [(5'h13):(1'h0)] reg1668 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1672 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1673 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1674 = (1'h0);
  reg [(5'h18):(1'h0)] reg1676 = (1'h0);
  reg [(4'hd):(1'h0)] reg1681 = (1'h0);
  reg [(4'hf):(1'h0)] reg1682 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1683 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1687 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1688 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1689 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1782 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1780 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1777 = (1'h0);
  reg [(4'hd):(1'h0)] reg1776 = (1'h0);
  reg [(3'h5):(1'h0)] reg1775 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1772 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1771 = (1'h0);
  reg [(4'he):(1'h0)] reg1768 = (1'h0);
  reg [(2'h3):(1'h0)] reg1767 = (1'h0);
  reg [(4'h8):(1'h0)] reg1765 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1763 = (1'h0);
  reg [(4'h8):(1'h0)] reg1762 = (1'h0);
  reg [(3'h6):(1'h0)] reg1758 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1749 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1754 = (1'h0);
  reg [(5'h17):(1'h0)] reg1753 = (1'h0);
  reg [(5'h15):(1'h0)] reg1752 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1749 = (1'h0);
  reg [(4'hb):(1'h0)] reg1746 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1745 = (1'h0);
  reg [(4'hb):(1'h0)] reg1741 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1740 = (1'h0);
  reg [(4'he):(1'h0)] reg1739 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1737 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1735 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1734 = (1'h0);
  reg [(2'h2):(1'h0)] reg1733 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1732 = (1'h0);
  reg [(4'he):(1'h0)] reg1721 = (1'h0);
  reg [(4'h8):(1'h0)] reg1727 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1726 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1724 = (1'h0);
  reg [(2'h3):(1'h0)] reg1723 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1722 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1721 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1719 = (1'h0);
  reg [(2'h2):(1'h0)] reg1717 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1715 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1713 = (1'h0);
  reg [(4'hb):(1'h0)] reg1712 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1711 = (1'h0);
  reg [(4'ha):(1'h0)] reg1710 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1709 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1708 = (1'h0);
  reg [(4'hd):(1'h0)] reg1706 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1705 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1700 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1702 = (1'h0);
  reg [(4'h8):(1'h0)] reg1700 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1698 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1696 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1686 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1685 = (1'h0);
  reg [(4'h8):(1'h0)] reg1684 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1671 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1680 = (1'h0);
  reg [(4'hc):(1'h0)] reg1679 = (1'h0);
  reg [(4'he):(1'h0)] reg1678 = (1'h0);
  reg [(4'h8):(1'h0)] reg1677 = (1'h0);
  reg [(5'h16):(1'h0)] reg1675 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1671 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1670 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1669 = (1'h0);
  reg [(5'h14):(1'h0)] reg1666 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1664 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1660 = (1'h0);
  reg [(5'h15):(1'h0)] reg1659 = (1'h0);
  reg [(5'h14):(1'h0)] reg1656 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1655 = (1'h0);
  reg [(5'h16):(1'h0)] reg1653 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1652 = (1'h0);
  reg [(2'h3):(1'h0)] reg1651 = (1'h0);
  reg [(5'h11):(1'h0)] reg1650 = (1'h0);
  reg [(4'hf):(1'h0)] reg1648 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1646 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1645 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1644 = (1'h0);
  reg [(5'h15):(1'h0)] reg1643 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1639 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1638 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1635 = (1'h0);
  reg [(3'h5):(1'h0)] reg1634 = (1'h0);
  reg [(2'h2):(1'h0)] reg355 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg354 = (1'h0);
  reg [(3'h4):(1'h0)] reg352 = (1'h0);
  reg [(2'h3):(1'h0)] reg351 = (1'h0);
  reg [(5'h13):(1'h0)] forvar348 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg348 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg346 = (1'h0);
  reg [(2'h2):(1'h0)] reg345 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg343 = (1'h0);
  reg [(4'h8):(1'h0)] reg342 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg339 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg22 = (1'h0);
  reg [(5'h18):(1'h0)] forvar20 = (1'h0);
  reg [(4'h8):(1'h0)] forvar19 = (1'h0);
  reg [(4'ha):(1'h0)] reg17 = (1'h0);
  reg [(4'he):(1'h0)] reg16 = (1'h0);
  reg [(2'h2):(1'h0)] reg14 = (1'h0);
  reg [(3'h6):(1'h0)] reg13 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg11 = (1'h0);
  reg [(2'h3):(1'h0)] reg10 = (1'h0);
  reg [(3'h4):(1'h0)] reg9 = (1'h0);
  reg [(3'h7):(1'h0)] reg8 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg6 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4 = (1'h0);
  assign y = {wire1769,
                 wire1707,
                 wire1631,
                 wire337,
                 wire24,
                 wire1690,
                 wire1691,
                 wire1693,
                 wire1694,
                 reg1783,
                 reg1781,
                 reg1779,
                 reg1778,
                 reg1774,
                 reg1773,
                 reg1770,
                 reg1766,
                 reg1764,
                 reg1761,
                 reg1760,
                 reg1759,
                 reg1757,
                 reg1756,
                 reg1755,
                 reg1751,
                 reg1750,
                 reg1748,
                 reg1747,
                 reg1744,
                 reg1743,
                 reg1742,
                 reg1738,
                 reg1736,
                 reg1731,
                 reg1730,
                 reg1729,
                 reg1728,
                 reg1726,
                 reg1725,
                 reg1720,
                 reg1718,
                 reg1716,
                 reg1714,
                 reg1704,
                 reg1703,
                 reg1698,
                 reg1701,
                 reg1699,
                 reg1697,
                 reg356,
                 reg353,
                 reg350,
                 reg349,
                 reg347,
                 reg344,
                 reg340,
                 reg23,
                 reg21,
                 reg18,
                 reg15,
                 reg12,
                 reg5,
                 reg1633,
                 reg1636,
                 reg1637,
                 reg1640,
                 reg1641,
                 reg1642,
                 reg1647,
                 reg1649,
                 reg1654,
                 reg1657,
                 reg1658,
                 reg1655,
                 reg1661,
                 reg1662,
                 reg1663,
                 reg1665,
                 reg1667,
                 reg1668,
                 reg1672,
                 reg1673,
                 reg1674,
                 reg1676,
                 reg1681,
                 reg1682,
                 reg1683,
                 reg1687,
                 reg1688,
                 reg1689,
                 reg1782,
                 reg1780,
                 reg1777,
                 reg1776,
                 reg1775,
                 forvar1772,
                 reg1771,
                 reg1768,
                 reg1767,
                 reg1765,
                 reg1763,
                 reg1762,
                 reg1758,
                 reg1749,
                 reg1754,
                 reg1753,
                 reg1752,
                 forvar1749,
                 reg1746,
                 reg1745,
                 reg1741,
                 reg1740,
                 reg1739,
                 reg1737,
                 reg1735,
                 forvar1734,
                 reg1733,
                 reg1732,
                 reg1721,
                 reg1727,
                 forvar1726,
                 reg1724,
                 reg1723,
                 reg1722,
                 forvar1721,
                 reg1719,
                 reg1717,
                 reg1715,
                 reg1713,
                 reg1712,
                 forvar1711,
                 reg1710,
                 reg1709,
                 reg1708,
                 reg1706,
                 reg1705,
                 forvar1700,
                 reg1702,
                 reg1700,
                 forvar1698,
                 forvar1696,
                 forvar1686,
                 forvar1685,
                 reg1684,
                 forvar1671,
                 reg1680,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1675,
                 reg1671,
                 reg1670,
                 reg1669,
                 reg1666,
                 forvar1664,
                 reg1660,
                 reg1659,
                 reg1656,
                 forvar1655,
                 reg1653,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1648,
                 forvar1646,
                 reg1645,
                 reg1644,
                 reg1643,
                 forvar1639,
                 forvar1638,
                 reg1635,
                 reg1634,
                 reg355,
                 reg354,
                 reg352,
                 reg351,
                 forvar348,
                 reg348,
                 reg346,
                 reg345,
                 reg343,
                 reg342,
                 reg341,
                 reg339,
                 reg22,
                 forvar20,
                 forvar19,
                 reg17,
                 reg16,
                 reg14,
                 reg13,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 forvar7,
                 reg6,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (2'h2)); forvar4 = (forvar4 + (1'h1)))
        begin
          reg5 <= wire0;
          reg6 = {$unsigned((!{(~|wire0)})),
              ((wire3 ?
                  $signed($unsigned(wire1)) : (((8'ha1) ? wire3 : wire3) ?
                      wire1 : $unsigned(wire2))) > ($signed(reg5[(1'h0):(1'h0)]) ?
                  wire2[(4'he):(1'h0)] : (wire0 ?
                      (^(8'hb1)) : $unsigned(wire0))))};
          for (forvar7 = (1'h0); (forvar7 < (3'h4)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg8 = (~$signed(wire2[(3'h6):(1'h1)]));
              reg9 = wire3[(3'h7):(2'h3)];
              reg10 = forvar4[(4'h8):(1'h1)];
            end
          if (($unsigned((~reg10)) ?
              reg10[(2'h2):(2'h2)] : reg9[(2'h3):(1'h1)]))
            begin
              reg11 = ((wire2[(4'hc):(3'h6)] >> ({(^~forvar7)} ?
                      (7'h43) : $signed(((8'h9f) ? forvar4 : wire0)))) ?
                  $signed($signed(({wire3, (8'haf)} ?
                      (wire2 ?
                          wire2 : reg5) : (+forvar7)))) : $unsigned({(((7'h46) ?
                          forvar4 : reg10) || reg6),
                      {$unsigned(forvar7), forvar4}}));
            end
          else
            begin
              reg12 <= $unsigned(reg10[(2'h3):(1'h0)]);
              reg13 = (reg6[(4'he):(2'h3)] ?
                  (~&(reg5 != reg11[(1'h0):(1'h0)])) : reg11[(1'h1):(1'h1)]);
              reg14 = (~|$signed(({wire1[(1'h1):(1'h0)]} ?
                  {$signed(reg9),
                      (~wire1)} : (reg11[(2'h2):(1'h1)] ~^ (reg6 > wire0)))));
              reg15 <= wire2;
              reg16 = $unsigned($signed({reg13[(2'h3):(2'h2)]}));
            end
        end
      reg17 = (!$unsigned(((reg8 ? (reg8 && (7'h44)) : {wire3}) ?
          $unsigned($signed(reg14)) : (~|$unsigned(reg15)))));
      reg18 <= {$unsigned(((((8'hbc) ? (8'haf) : (8'hae)) ?
              (reg6 ? reg8 : reg16) : (reg17 ? reg8 : reg17)) <<< {{(7'h41),
                  wire1}})),
          $unsigned({{(forvar7 ? reg11 : wire1)}, $signed((^reg8))})};
      for (forvar19 = (1'h0); (forvar19 < (1'h0)); forvar19 = (forvar19 + (1'h1)))
        begin
          for (forvar20 = (1'h0); (forvar20 < (1'h0)); forvar20 = (forvar20 + (1'h1)))
            begin
              reg21 <= (wire1 ?
                  forvar4 : ($signed($unsigned(reg6)) ?
                      reg17[(3'h5):(2'h2)] : (~^$signed(forvar7))));
              reg22 = (-wire0[(4'hf):(1'h1)]);
            end
          reg23 <= reg15;
        end
    end
  assign wire24 = $unsigned($signed($signed($unsigned({reg12}))));
  module25 #() modinst338 (wire337, clk, reg23, wire0, wire1, reg21);
  always
    @(posedge clk) begin
      if (wire2[(2'h3):(1'h1)])
        begin
          reg339 = ((($unsigned($unsigned(reg23)) ?
                  $signed(reg18[(3'h7):(1'h0)]) : ($signed((8'hbc)) ^ (reg23 ?
                      reg12 : wire2))) ^ {$unsigned((reg12 >>> wire337))}) ?
              ((~|({wire337} ^ $unsigned(wire337))) ?
                  $unsigned({$unsigned(wire337)}) : (-(!{wire0}))) : (&$signed({wire24[(4'hd):(2'h2)],
                  reg12})));
        end
      else
        begin
          if ($signed(($signed(wire3[(4'he):(3'h5)]) || ((~&(reg15 != reg339)) << ($signed((8'hac)) && (wire1 >= (8'ha4)))))))
            begin
              reg340 <= (reg23 > wire2[(4'hd):(3'h6)]);
            end
          else
            begin
              reg339 = ($signed($signed(((&reg21) == reg5))) ?
                  wire1[(4'ha):(3'h7)] : (~wire24));
              reg340 <= $unsigned(wire1);
              reg341 = ((8'h9d) <= {{reg12, wire337[(1'h1):(1'h0)]},
                  (!(^~(reg5 >= (8'hb8))))});
              reg342 = (~|($unsigned(($signed(wire2) ~^ $unsigned(reg5))) ?
                  (|wire3[(4'h8):(3'h7)]) : $unsigned($unsigned({reg18}))));
            end
          reg343 = (reg340[(1'h1):(1'h0)] * $unsigned(($unsigned({reg340,
              reg12}) && $unsigned({wire0}))));
          reg344 <= $unsigned((^~({(wire24 ?
                  wire3 : reg339)} >= (~$unsigned(reg342)))));
        end
      reg345 = (reg21[(4'h9):(3'h7)] ~^ (8'h9d));
    end
  always
    @(posedge clk) begin
      reg346 = reg15[(4'hb):(4'ha)];
      if (reg344[(4'he):(2'h3)])
        begin
          if (wire24[(2'h2):(2'h2)])
            begin
              reg347 <= {{{(((8'hb4) < reg340) ? (-wire3) : $unsigned(reg5))},
                      wire3}};
              reg348 = $unsigned(($unsigned(($signed(wire1) || (reg347 <<< wire1))) ?
                  reg344[(4'hb):(4'hb)] : (wire2[(4'hb):(3'h6)] + ((&wire0) << wire3))));
            end
          else
            begin
              reg348 = {(+({wire3} ?
                      $unsigned(reg5[(2'h2):(1'h1)]) : (^((7'h42) <= reg346)))),
                  $unsigned(reg344)};
              reg349 <= {wire24[(4'hd):(3'h6)]};
            end
        end
      else
        begin
          reg347 <= ($signed((((wire24 + reg18) * (^~(8'h9c))) ~^ reg21)) >= wire1[(2'h2):(1'h0)]);
          for (forvar348 = (1'h0); (forvar348 < (2'h3)); forvar348 = (forvar348 + (1'h1)))
            begin
              reg349 <= (~wire3[(2'h3):(2'h2)]);
              reg350 <= ($signed($unsigned({((8'ha7) || wire24)})) ^~ $unsigned($signed((wire337 || (-reg346)))));
              reg351 = reg340[(2'h2):(2'h2)];
              reg352 = (((8'hb8) | ({$unsigned(wire0)} ?
                      $unsigned($signed(reg344)) : wire1[(3'h4):(1'h1)])) ?
                  reg350 : (({{reg350, wire1}} ?
                          ({reg348} ?
                              $unsigned((8'hbc)) : (reg348 ?
                                  reg349 : reg21)) : wire24[(1'h1):(1'h0)]) ?
                      {((forvar348 ?
                              (7'h44) : wire24) > $unsigned(reg348))} : {$signed((+reg12)),
                          (^$signed(reg21))}));
            end
        end
    end
  always
    @(posedge clk) begin
      reg353 <= {wire337[(4'h8):(3'h6)], (8'ha9)};
      reg354 = (+reg353[(1'h0):(1'h0)]);
      reg355 = $signed((8'hb6));
      reg356 <= reg18[(4'hd):(3'h4)];
    end
  module357 #() modinst1632 (wire1631, clk, wire1, reg23, reg344, reg349);
  always
    @(posedge clk) begin
      reg1633 <= wire0;
      reg1634 = wire24;
      reg1635 = $signed($signed($signed((^~$unsigned(wire3)))));
    end
  always
    @(posedge clk) begin
      reg1636 <= (!wire2);
      reg1637 <= wire24;
    end
  always
    @(posedge clk) begin
      for (forvar1638 = (1'h0); (forvar1638 < (1'h0)); forvar1638 = (forvar1638 + (1'h1)))
        begin
          for (forvar1639 = (1'h0); (forvar1639 < (2'h2)); forvar1639 = (forvar1639 + (1'h1)))
            begin
              reg1640 <= $signed(reg347[(2'h3):(1'h1)]);
              reg1641 <= ((reg350[(4'h8):(3'h5)] ?
                  (&{$signed((8'h9e))}) : wire1[(3'h4):(2'h3)]) >> (&{$unsigned((+reg340))}));
              reg1642 <= $signed($signed($unsigned(((wire0 > reg353) >>> (&reg18)))));
            end
          reg1643 = wire24;
          reg1644 = {(wire3[(5'h11):(4'hb)] >> ((&(wire3 ? wire24 : wire24)) ?
                  wire1 : $unsigned($unsigned(reg1641)))),
              $signed(reg1642[(4'he):(4'ha)])};
          reg1645 = reg349[(5'h11):(5'h11)];
          for (forvar1646 = (1'h0); (forvar1646 < (1'h1)); forvar1646 = (forvar1646 + (1'h1)))
            begin
              reg1647 <= $unsigned((reg15[(4'hb):(3'h7)] ?
                  reg353 : $unsigned(((reg349 ? reg5 : reg349) ?
                      {reg21, forvar1639} : (reg350 ? reg1642 : reg23)))));
              reg1648 = $unsigned($unsigned($unsigned(reg1633[(5'h16):(4'hf)])));
              reg1649 <= ((8'hb2) != {{$signed(forvar1646),
                      {forvar1646[(3'h5):(2'h2)]}},
                  $unsigned(reg1633[(2'h2):(1'h0)])});
              reg1650 = wire2[(2'h2):(2'h2)];
              reg1651 = $unsigned($signed($signed(forvar1639)));
            end
        end
      if ((reg344 | {(((reg1650 ^ reg1642) ?
              $signed(wire2) : $signed(wire3)) & ($unsigned(reg1647) ?
              (reg349 ? wire337 : reg356) : {wire24})),
          $signed($signed(((8'ha1) ? reg1648 : wire337)))}))
        begin
          reg1652 = $signed($unsigned(forvar1639[(4'hb):(4'ha)]));
          reg1653 = {($unsigned(((reg356 > wire3) ?
                      $unsigned(reg15) : (&reg1652))) ?
                  reg344[(1'h1):(1'h1)] : reg12[(1'h0):(1'h0)])};
          reg1654 <= reg1645[(3'h4):(1'h1)];
          for (forvar1655 = (1'h0); (forvar1655 < (3'h4)); forvar1655 = (forvar1655 + (1'h1)))
            begin
              reg1656 = reg1645;
              reg1657 <= forvar1646[(5'h11):(4'h8)];
              reg1658 <= reg1647[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg1654 <= (8'ha1);
          if ($signed($unsigned($unsigned(((8'ha4) + wire2)))))
            begin
              reg1655 <= (~($unsigned($signed(reg5)) <<< reg353[(1'h0):(1'h0)]));
              reg1657 <= $signed((wire24 ?
                  ({$unsigned(wire2), {reg1637, forvar1638}} ?
                      ((reg1647 >= (7'h4a)) ?
                          $unsigned(forvar1638) : $signed((8'hb8))) : $signed((reg340 ?
                          wire24 : (7'h45)))) : $signed(wire337[(1'h0):(1'h0)])));
            end
          else
            begin
              reg1655 <= reg350;
              reg1656 = $signed(forvar1638);
              reg1659 = $unsigned({($signed($signed((7'h42))) + ($unsigned((8'hb2)) || reg1652))});
            end
          if ((7'h44))
            begin
              reg1660 = (($unsigned(forvar1646) ?
                      $unsigned(((~(8'ha1)) * (reg1652 ?
                          (8'hb7) : reg1650))) : $signed(reg23[(3'h7):(3'h6)])) ?
                  $signed({((~wire3) <= reg340[(4'he):(4'he)])}) : reg1643);
            end
          else
            begin
              reg1660 = {($signed($signed($signed(reg5))) ?
                      reg347[(2'h2):(2'h2)] : {$signed(reg1642[(5'h10):(3'h7)]),
                          $signed(reg1633)})};
              reg1661 <= reg1652[(4'hf):(4'h9)];
              reg1662 <= (&({(reg350[(3'h7):(3'h4)] || ((8'ha8) < reg1644)),
                  reg1653[(4'h8):(3'h4)]} ^~ {$signed($unsigned(reg1655))}));
              reg1663 <= $signed($unsigned($unsigned($unsigned($unsigned(reg356)))));
            end
          for (forvar1664 = (1'h0); (forvar1664 < (1'h1)); forvar1664 = (forvar1664 + (1'h1)))
            begin
              reg1665 <= ((~|(($signed((8'hb1)) ?
                      (!forvar1638) : reg1655[(1'h1):(1'h1)]) ?
                  reg1648 : reg353)) < reg1644);
              reg1666 = (&reg350);
              reg1667 <= ({(~{(reg347 + reg23), (wire24 >> reg1666)})} ?
                  reg356[(4'h9):(4'h9)] : ((reg1652[(1'h0):(1'h0)] <= wire2[(4'hd):(1'h0)]) | $signed({reg1633})));
              reg1668 <= reg1659;
            end
        end
      if ($signed(($signed($unsigned($unsigned(forvar1664))) > $unsigned(forvar1638[(1'h1):(1'h1)]))))
        begin
          if ((reg1658 == (~|reg1658[(2'h2):(2'h2)])))
            begin
              reg1669 = (&(!$unsigned($signed(reg1658[(4'ha):(3'h7)]))));
              reg1670 = $signed($signed((((wire337 ? reg1654 : reg1640) ?
                      $unsigned(reg12) : reg1663[(2'h2):(1'h1)]) ?
                  {$signed(reg1667)} : (forvar1664 * $unsigned(forvar1655)))));
              reg1671 = $signed(reg1656);
              reg1672 <= $unsigned({reg21,
                  (|((reg1655 ? (8'ha8) : wire0) << reg1642))});
            end
          else
            begin
              reg1672 <= (~|reg1669[(2'h2):(1'h1)]);
            end
          if ((~$signed($signed(($signed(reg349) ?
              reg1650[(4'h9):(4'h9)] : $unsigned(reg1644))))))
            begin
              reg1673 <= (reg1670[(2'h3):(1'h0)] ?
                  {reg1667[(2'h2):(1'h1)],
                      $signed(forvar1638)} : $unsigned((~&(!((8'ha6) ?
                      reg353 : reg1652)))));
            end
          else
            begin
              reg1673 <= (($unsigned(($signed(reg1666) ?
                          wire1631[(3'h7):(2'h3)] : (&reg1640))) ?
                      $unsigned($signed((reg1665 < reg1651))) : (forvar1639[(3'h4):(1'h1)] ?
                          $unsigned(reg1650) : ((reg1663 ?
                              reg18 : reg1670) << reg1648))) ?
                  (reg12[(2'h2):(1'h0)] ?
                      reg1662 : $signed((reg1644[(4'hc):(3'h4)] ?
                          (~^(8'hb3)) : (&(7'h48))))) : forvar1638);
              reg1674 <= reg353[(1'h0):(1'h0)];
            end
          reg1675 = (reg1668 & reg349);
          if ({({$unsigned(reg1647[(3'h6):(3'h4)])} ?
                  (((reg1660 * reg1653) ? reg1643 : (-wire1631)) ?
                      (!(^~forvar1655)) : (^{reg349})) : $unsigned((~|(~(8'hbf)))))})
            begin
              reg1676 <= reg344;
            end
          else
            begin
              reg1677 = {($signed($unsigned(wire24[(4'he):(1'h0)])) < ($unsigned($signed((8'h9d))) * $signed({(8'h9e),
                      reg1652})))};
            end
          if ($signed($signed(reg349)))
            begin
              reg1678 = reg1669[(2'h3):(1'h1)];
              reg1679 = reg350;
              reg1680 = reg1675[(4'he):(3'h5)];
            end
          else
            begin
              reg1678 = (~((+$unsigned((8'h9e))) ? reg349 : {(~(^~reg1674))}));
              reg1679 = $unsigned(reg1662[(1'h1):(1'h0)]);
            end
        end
      else
        begin
          reg1669 = (&reg1653[(5'h10):(4'he)]);
          reg1670 = reg350[(3'h4):(1'h0)];
          for (forvar1671 = (1'h0); (forvar1671 < (3'h4)); forvar1671 = (forvar1671 + (1'h1)))
            begin
              reg1675 = (reg1655[(3'h5):(1'h1)] ?
                  $signed(((8'ha0) ~^ (+reg1674[(5'h12):(4'ha)]))) : ((~|$unsigned((reg1672 != reg1666))) ^~ $signed(reg1653)));
              reg1676 <= (&(((reg1658[(4'he):(1'h1)] ?
                          $unsigned(forvar1646) : $unsigned(reg356)) ?
                      (reg1680 ^~ $unsigned(reg21)) : {(reg15 ?
                              (8'ha9) : reg356)}) ?
                  (~^reg1645) : reg1645));
              reg1681 <= $unsigned(reg1654);
              reg1682 <= (((~|reg1669) ?
                  {reg350[(4'ha):(4'ha)],
                      ({(8'hbc)} ?
                          $signed(reg344) : (reg1663 ?
                              reg1665 : wire24))} : reg1671[(1'h1):(1'h0)]) ^ $signed({$unsigned((forvar1664 ?
                      reg1671 : reg344))}));
              reg1683 <= (~((!reg1671) ?
                  ($signed(wire1631[(2'h2):(1'h1)]) ?
                      {((8'hab) ?
                              reg1663 : reg1682)} : {(+(8'ha9))}) : (((~^reg1659) ?
                      ((8'ha7) ? (7'h4a) : reg340) : (reg1637 ?
                          reg12 : reg1675)) >> reg1671[(3'h7):(3'h5)])));
            end
          reg1684 = (((8'ha8) ?
              $unsigned(($signed(forvar1638) ?
                  $unsigned(reg356) : (~forvar1639))) : forvar1655[(2'h3):(1'h0)]) >>> $signed((~|wire24)));
        end
      for (forvar1685 = (1'h0); (forvar1685 < (1'h1)); forvar1685 = (forvar1685 + (1'h1)))
        begin
          for (forvar1686 = (1'h0); (forvar1686 < (2'h3)); forvar1686 = (forvar1686 + (1'h1)))
            begin
              reg1687 <= (+(((~^reg1645) ?
                  reg344[(3'h7):(3'h6)] : $unsigned($signed(forvar1685))) - (~$unsigned((reg1640 ~^ (7'h46))))));
              reg1688 <= (~&(~&(8'ha9)));
              reg1689 <= {$signed({{{forvar1639}, $signed(reg12)}})};
            end
        end
    end
  assign wire1690 = ($unsigned((reg1674[(5'h14):(1'h0)] >>> $unsigned($signed(reg1674)))) ?
                        (&$signed(reg1663[(1'h1):(1'h1)])) : reg356[(1'h0):(1'h0)]);
  module25 #() modinst1692 (wire1691, clk, reg23, reg18, reg1667, reg1640);
  assign wire1693 = $unsigned((8'ha5));
  module25 #() modinst1695 (.wire28(reg1662), .clk(clk), .wire27(reg15), .y(wire1694), .wire26(wire337), .wire29(reg1655));
  always
    @(posedge clk) begin
      for (forvar1696 = (1'h0); (forvar1696 < (2'h3)); forvar1696 = (forvar1696 + (1'h1)))
        begin
          reg1697 <= {(~&$signed($unsigned((^reg1673)))),
              $unsigned(reg18[(1'h1):(1'h0)])};
        end
      if ((reg350 ? reg1640 : $unsigned($unsigned({wire1, $signed(reg1640)}))))
        begin
          for (forvar1698 = (1'h0); (forvar1698 < (1'h1)); forvar1698 = (forvar1698 + (1'h1)))
            begin
              reg1699 <= reg1640[(4'h8):(1'h0)];
              reg1700 = (|reg23);
              reg1701 <= $signed((~^(!wire337)));
            end
          reg1702 = {(8'ha9)};
        end
      else
        begin
          reg1698 <= reg347[(2'h2):(1'h1)];
          reg1699 <= (~|reg350[(3'h4):(3'h4)]);
          for (forvar1700 = (1'h0); (forvar1700 < (2'h2)); forvar1700 = (forvar1700 + (1'h1)))
            begin
              reg1701 <= $unsigned(reg1665[(1'h1):(1'h0)]);
              reg1702 = ($unsigned(wire24[(4'ha):(4'ha)]) & $signed($unsigned((^~$signed(wire3)))));
              reg1703 <= $unsigned($signed(reg18[(1'h0):(1'h0)]));
              reg1704 <= $signed(($signed((^~reg5)) != $signed((-wire1))));
              reg1705 = reg349[(4'hb):(4'h8)];
            end
        end
      reg1706 = reg1688[(2'h2):(1'h0)];
    end
  assign wire1707 = $unsigned(reg1667);
  always
    @(posedge clk) begin
      if ($signed($unsigned($unsigned((^~reg1688)))))
        begin
          reg1708 = $unsigned($signed($unsigned($signed(reg1633[(4'he):(3'h4)]))));
          reg1709 = ((({$signed(reg1667), ((7'h41) ? wire3 : (8'ha9))} ?
                  $unsigned(reg1704[(1'h1):(1'h1)]) : ((+reg1637) ?
                      ((7'h43) + reg356) : $signed(reg1668))) ?
              (($unsigned(wire2) ? wire1690 : (8'h9d)) && ((~reg1683) ?
                  {reg1708} : (reg1687 ?
                      wire1631 : wire3))) : (({reg1688} > (^reg1647)) * $signed(reg1663[(4'ha):(3'h4)]))) + $signed(reg1633));
        end
      else
        begin
          reg1708 = (reg356[(3'h4):(2'h3)] <= $signed((((reg1676 + reg1655) * (~^reg1640)) ?
              $unsigned((reg1683 * reg344)) : reg12)));
        end
      reg1710 = $signed($unsigned((-$signed($unsigned(wire0)))));
      if (reg1673)
        begin
          for (forvar1711 = (1'h0); (forvar1711 < (2'h2)); forvar1711 = (forvar1711 + (1'h1)))
            begin
              reg1712 = (^reg1662);
              reg1713 = $unsigned(reg21[(3'h4):(2'h2)]);
              reg1714 <= reg1704[(3'h5):(2'h3)];
            end
          if ((~&reg1657))
            begin
              reg1715 = $signed({(($unsigned(reg1682) ?
                      $unsigned((7'h4a)) : {reg1672}) >>> reg356[(3'h4):(1'h1)])});
            end
          else
            begin
              reg1716 <= reg1714[(4'h8):(2'h3)];
              reg1717 = reg1701[(1'h0):(1'h0)];
              reg1718 <= (((-{(reg1713 ? (8'ha5) : reg1640),
                          (reg1699 ? reg340 : reg350)}) ?
                      reg1699[(4'he):(4'he)] : reg15[(4'hb):(3'h5)]) ?
                  $unsigned(($unsigned(reg1709[(4'hb):(4'ha)]) ?
                      reg1636 : reg1683)) : (($signed($unsigned(reg350)) || wire1693[(2'h2):(1'h1)]) > ((reg15[(4'hb):(4'ha)] ?
                      wire1[(4'hf):(3'h6)] : ((8'ha3) < reg1698)) ^ $unsigned(reg1676))));
              reg1719 = (~&(((^(-reg1637)) + {$unsigned(reg1718)}) || reg12));
              reg1720 <= reg1716[(1'h0):(1'h0)];
            end
          for (forvar1721 = (1'h0); (forvar1721 < (1'h0)); forvar1721 = (forvar1721 + (1'h1)))
            begin
              reg1722 = ($unsigned({$signed({reg1714})}) <= reg1703[(1'h0):(1'h0)]);
              reg1723 = ((wire1694[(1'h0):(1'h0)] & ($signed(reg1662[(3'h6):(3'h4)]) ?
                  ((8'hbe) & (wire24 ?
                      reg18 : reg1708)) : $signed($signed(reg353)))) != ((($unsigned(wire3) > (wire0 != reg1682)) ?
                      ((~reg23) >>> (reg1683 ?
                          reg1672 : reg1717)) : {reg1719[(4'hd):(4'hd)],
                          reg1720[(3'h5):(2'h2)]}) ?
                  {$unsigned((8'ha2)),
                      (&(reg21 && reg1683))} : (|(reg1701[(4'ha):(4'h8)] ?
                      {reg1658} : (reg1687 ? wire1691 : (8'hb2))))));
              reg1724 = ($signed($unsigned((!reg1636))) ?
                  $signed({reg23[(5'h17):(3'h7)],
                      {reg1641[(1'h1):(1'h1)]}}) : $unsigned(wire1[(4'hf):(4'hf)]));
            end
          reg1725 <= {$unsigned($signed(((wire1690 ?
                  reg1665 : reg1682) * reg1657)))};
          for (forvar1726 = (1'h0); (forvar1726 < (1'h1)); forvar1726 = (forvar1726 + (1'h1)))
            begin
              reg1727 = (~$unsigned((reg1724 ?
                  reg350[(2'h2):(1'h1)] : (reg1658 ?
                      $unsigned(wire1693) : $unsigned(reg1688)))));
            end
        end
      else
        begin
          for (forvar1711 = (1'h0); (forvar1711 < (2'h3)); forvar1711 = (forvar1711 + (1'h1)))
            begin
              reg1714 <= reg1717[(2'h2):(1'h0)];
            end
          if ((8'had))
            begin
              reg1715 = (wire1693 ?
                  $unsigned(wire24[(4'hf):(4'hc)]) : (~&reg12[(2'h2):(2'h2)]));
            end
          else
            begin
              reg1716 <= $signed((^((~|(reg1682 ^ reg1718)) >> (wire2[(4'hd):(4'h9)] ?
                  $signed(reg1709) : {wire1694}))));
              reg1717 = reg1688[(3'h4):(3'h4)];
              reg1719 = ($signed((wire1690[(1'h1):(1'h1)] ?
                  $signed((reg356 ?
                      reg1674 : reg1715)) : $signed($unsigned(reg353)))) >= reg350);
              reg1721 = {reg1682[(4'ha):(2'h3)]};
              reg1722 = reg1640[(4'hd):(1'h0)];
            end
          if ((reg1667 ? reg1658 : (~|$signed((^(reg1637 != reg349))))))
            begin
              reg1725 <= ((($unsigned((wire1694 ?
                          reg1668 : reg1676)) >= ((wire2 >> reg1661) ?
                          {reg15} : (~reg1708))) ?
                      $unsigned({reg1676,
                          (reg349 << forvar1721)}) : (~&(reg1655 ?
                          {reg1667} : (^wire1693)))) ?
                  wire0[(4'hb):(4'hb)] : (($unsigned((8'ha6)) == (~|$signed(reg353))) ?
                      wire3[(4'he):(4'hc)] : $signed($signed(((7'h44) << reg356)))));
            end
          else
            begin
              reg1725 <= {((~|(-$unsigned(reg1719))) || (~(reg1654 ?
                      {reg1636} : (reg1698 << reg1636))))};
              reg1726 <= {reg1709};
            end
          if ((^((+(((8'ha1) ? reg18 : reg344) ?
                  $signed(reg1676) : ((8'hb9) ? reg1641 : reg1721))) ?
              reg1703 : (reg1665[(1'h0):(1'h0)] ?
                  ((reg1641 ^ (8'ha6)) ?
                      (reg1641 < reg1712) : $unsigned(reg1718)) : $signed($signed(reg1641))))))
            begin
              reg1727 = {reg1713,
                  ($unsigned({(7'h46), ((8'hbe) <<< forvar1726)}) ?
                      (((wire337 ? reg1703 : (8'ha8)) ?
                              $signed(reg1699) : {wire1694, reg15}) ?
                          reg1717 : reg1674[(3'h4):(3'h4)]) : (8'hb7))};
              reg1728 <= (~&((($unsigned(reg353) ^ wire2) || ((^reg1665) ?
                  (~wire2) : wire1690)) && ((~^wire337) ?
                  ((8'ha7) < $signed(reg1688)) : {{reg1662, reg1681}})));
              reg1729 <= ({(7'h49)} & reg1674[(4'hc):(1'h1)]);
              reg1730 <= reg1729[(5'h12):(4'he)];
              reg1731 <= reg1661[(3'h6):(3'h6)];
            end
          else
            begin
              reg1728 <= (({(~&reg1665[(2'h3):(1'h1)]), reg1704} ?
                  {{$unsigned(reg1687), (!reg1723)},
                      $signed((8'ha2))} : reg1730[(3'h7):(3'h7)]) >= {$unsigned(((reg1647 <= reg1701) ?
                      reg1672 : reg1720[(1'h0):(1'h0)])),
                  reg1699});
              reg1729 <= {reg1730[(4'h9):(3'h4)], reg1637};
              reg1732 = {$unsigned($signed(($unsigned((8'hb0)) <<< wire0[(4'hc):(4'h9)]))),
                  reg1697[(3'h7):(1'h1)]};
              reg1733 = reg1640;
            end
        end
      for (forvar1734 = (1'h0); (forvar1734 < (1'h1)); forvar1734 = (forvar1734 + (1'h1)))
        begin
          if (($unsigned((^~({(8'hb7),
              reg1729} && reg1637))) && $unsigned({(+reg1715)})))
            begin
              reg1735 = (7'h42);
            end
          else
            begin
              reg1736 <= ($unsigned((!($unsigned(reg1713) >>> (8'ha8)))) < wire2);
              reg1737 = (^~reg1712[(1'h1):(1'h1)]);
              reg1738 <= $unsigned(($unsigned($unsigned(forvar1711[(3'h5):(2'h2)])) ?
                  (&(reg1720 ?
                      reg1715[(2'h2):(1'h0)] : (reg353 != reg1720))) : ($unsigned(((8'hac) ?
                      reg23 : reg1718)) != ($signed(reg1720) ?
                      $signed(wire0) : wire1691[(2'h3):(1'h0)]))));
              reg1739 = {{(|(^~((8'ha4) ? reg1699 : reg1712))),
                      (~^(reg1642[(1'h0):(1'h0)] ?
                          reg1735[(5'h10):(4'h8)] : (reg1709 ^ reg1641)))}};
            end
          if (($signed(wire1) >>> (+$signed(($signed(reg23) ?
              (8'ha7) : reg12)))))
            begin
              reg1740 = (~&reg1736[(2'h2):(1'h1)]);
              reg1741 = wire24[(4'h8):(4'h8)];
              reg1742 <= {{reg349[(5'h10):(4'h8)]},
                  $signed(($signed(reg5[(2'h2):(1'h0)]) ?
                      ($unsigned(reg1722) ?
                          $signed(reg1716) : reg1725[(3'h6):(3'h5)]) : {(reg1725 <= reg1661),
                          reg1663}))};
              reg1743 <= ((~$signed((reg347[(2'h2):(1'h0)] >> reg347))) ?
                  (~^reg15[(1'h0):(1'h0)]) : {(reg1726 & ((reg1717 >= (8'haf)) - reg1724[(2'h2):(1'h1)]))});
            end
          else
            begin
              reg1740 = (($signed((8'hbc)) ?
                      (~&((reg1703 ?
                          reg1703 : wire1690) << reg15[(4'h9):(3'h6)])) : $unsigned((+(7'h42)))) ?
                  (~&(~|reg1683[(5'h11):(2'h2)])) : forvar1711[(1'h1):(1'h1)]);
            end
          if (reg1641[(2'h2):(1'h1)])
            begin
              reg1744 <= (+reg1661[(1'h0):(1'h0)]);
            end
          else
            begin
              reg1745 = ({(+$unsigned(reg353[(3'h4):(1'h0)])),
                  reg1701[(1'h0):(1'h0)]} == reg1654);
              reg1746 = (~^($signed(((reg1709 ? forvar1721 : reg1640) ?
                  {reg1726} : reg1715)) || (reg1703 ?
                  (reg1742[(1'h1):(1'h1)] ?
                      reg1663[(3'h6):(1'h0)] : reg1661) : $signed(wire1690[(4'h8):(2'h2)]))));
              reg1747 <= (^~$unsigned(({(reg1719 ? reg12 : wire1690),
                  (^reg1730)} > $signed(reg1729[(5'h10):(4'h8)]))));
              reg1748 <= $unsigned($unsigned((8'ha3)));
            end
        end
      if ((((&(~(reg1654 ? reg350 : reg21))) ?
          $signed(((reg1657 + reg1719) ?
              {reg1647,
                  reg1748} : reg1733)) : {$signed(reg349[(4'hb):(3'h6)])}) != ($unsigned($signed($signed(reg1739))) * reg1640[(4'hb):(3'h6)])))
        begin
          for (forvar1749 = (1'h0); (forvar1749 < (2'h3)); forvar1749 = (forvar1749 + (1'h1)))
            begin
              reg1750 <= (((^$unsigned((|(8'h9d)))) ?
                  (~&(^~$signed((8'ha9)))) : (+$signed($signed((8'hae))))) * (!$unsigned($signed((reg1714 ?
                  (8'hb0) : reg1728)))));
              reg1751 <= (reg1697 ?
                  (~|(&($unsigned(reg1640) << (~^reg1716)))) : ($signed($unsigned({(8'hb3)})) ?
                      forvar1749 : reg1747));
              reg1752 = (reg1731 ?
                  $unsigned({(!(^reg1715)),
                      wire1631}) : (reg1703[(3'h4):(1'h0)] ?
                      $unsigned({(wire24 ? reg1688 : reg1662),
                          (^wire1691)}) : ({(^~reg1640)} ?
                          reg21[(4'hf):(1'h1)] : reg1724[(1'h1):(1'h0)])));
              reg1753 = $unsigned((((8'h9e) ^ (reg1715[(1'h0):(1'h0)] && $unsigned(forvar1749))) ^ reg1738));
            end
          if ((7'h42))
            begin
              reg1754 = (~&reg1633[(3'h6):(1'h0)]);
            end
          else
            begin
              reg1755 <= reg1649;
            end
          reg1756 <= reg356[(4'hb):(2'h3)];
        end
      else
        begin
          reg1749 = {{$signed($signed($signed(reg356)))}};
          if ((reg1640 ? $unsigned(reg15) : reg1673))
            begin
              reg1750 <= reg1731[(3'h4):(2'h3)];
            end
          else
            begin
              reg1750 <= reg1673;
              reg1752 = forvar1721;
              reg1755 <= {reg1732[(3'h6):(1'h0)]};
              reg1756 <= (~(reg18 ?
                  (&forvar1711) : $signed((reg1733 ?
                      {reg1682} : (forvar1721 ? (7'h46) : reg1713)))));
            end
          reg1757 <= $signed({((+(+reg1730)) ?
                  ((^~(8'hb8)) ?
                      $unsigned(reg1721) : $signed(reg1723)) : $unsigned((+reg1725))),
              reg1728});
          if (wire1[(3'h6):(3'h5)])
            begin
              reg1758 = wire1693[(3'h4):(3'h4)];
              reg1759 <= {(reg23 << reg349[(4'hc):(1'h0)]),
                  $unsigned($signed((~&$signed(reg1722))))};
              reg1760 <= reg1735[(4'hf):(4'hd)];
              reg1761 <= (|$unsigned({{reg356}}));
            end
          else
            begin
              reg1759 <= $signed({reg1699});
              reg1762 = ($unsigned({((&reg1744) <<< (reg1642 ?
                          reg1752 : reg1743)),
                      (-$unsigned(reg1714))}) ?
                  {reg1753[(5'h14):(4'h9)]} : {reg1753, wire1694});
              reg1763 = reg1688[(4'h9):(3'h6)];
            end
          if ((-(+(~&((-reg1658) ? (reg1718 + reg1708) : forvar1711)))))
            begin
              reg1764 <= reg1676[(3'h6):(3'h5)];
              reg1765 = ((reg1763 << ((8'hab) ?
                      ((~&reg1641) ?
                          (reg1683 ?
                              (8'hbf) : reg15) : (reg1758 || (7'h48))) : reg1732[(3'h6):(2'h2)])) ?
                  {reg1712[(1'h0):(1'h0)]} : $unsigned($unsigned($unsigned($unsigned(wire3)))));
              reg1766 <= $unsigned(((8'hbd) ?
                  (({reg1717, reg1640} ?
                      reg1756 : (+reg1688)) << ((^reg1753) ^ (reg1654 ?
                      reg1754 : reg1665))) : (reg1736 ~^ $unsigned(((8'had) ?
                      reg1699 : reg1744)))));
            end
          else
            begin
              reg1765 = (reg1747 ?
                  (8'hb9) : ($unsigned(reg1654[(3'h5):(3'h4)]) ?
                      (reg1739 == $signed((reg1719 < reg1756))) : (((reg1724 || forvar1734) ?
                          $unsigned(reg1709) : {reg1723,
                              (7'h40)}) ^~ reg1654)));
              reg1767 = ($unsigned(reg1688) ?
                  $unsigned((~|reg1724)) : $unsigned((7'h46)));
              reg1768 = (!(~&$unsigned($unsigned(forvar1726))));
            end
        end
    end
  assign wire1769 = $unsigned({(~^reg1668[(5'h11):(5'h10)]),
                        (((reg1676 ? reg1636 : reg1654) ?
                                {reg1729, wire1694} : $unsigned((8'ha9))) ?
                            wire24 : (-reg1688[(2'h3):(1'h1)]))});
  always
    @(posedge clk) begin
      reg1770 <= reg1757;
      reg1771 = (^~{($unsigned((^~reg1657)) <<< reg1756)});
      for (forvar1772 = (1'h0); (forvar1772 < (2'h3)); forvar1772 = (forvar1772 + (1'h1)))
        begin
          reg1773 <= (!$signed($signed($signed($unsigned(wire1)))));
          reg1774 <= (reg1742[(3'h7):(3'h5)] - (~reg1661));
          reg1775 = ({$unsigned($unsigned((^~reg1736))),
                  $unsigned((&$unsigned(reg1744)))} ?
              $signed((-($signed(reg1731) != (reg1674 | reg1738)))) : {((^~(&reg340)) != (^(reg340 ?
                      wire2 : (8'hba)))),
                  ((-(reg1665 ~^ reg1756)) ?
                      {(reg1774 ? reg1682 : reg1636)} : ((~&reg1654) ?
                          reg1665[(3'h7):(3'h4)] : (reg1714 + reg1703)))});
          if (reg1663)
            begin
              reg1776 = $unsigned($unsigned({(~|(reg1738 - reg344))}));
              reg1777 = ($unsigned(reg1703[(2'h2):(1'h1)]) ?
                  reg1776 : (reg1775[(1'h1):(1'h0)] <= ($signed($signed(wire1690)) != reg1663[(4'h8):(4'h8)])));
              reg1778 <= (&($signed($signed(reg344[(4'ha):(2'h2)])) ?
                  (~^(((8'h9c) ?
                      reg1689 : (8'hb2)) * reg340)) : reg12[(1'h0):(1'h0)]));
              reg1779 <= (($signed({wire2,
                      reg1744}) == $unsigned($unsigned(wire1694[(4'ha):(4'ha)]))) ?
                  ((8'ha8) * reg1668) : ({(8'ha1), {{wire1691}, (~reg349)}} ?
                      ($signed(reg1672[(2'h2):(2'h2)]) ?
                          $signed($unsigned(reg1689)) : ((reg1657 >= reg1673) ?
                              (-reg1676) : (reg1738 && reg1718))) : (|(8'h9f))));
            end
          else
            begin
              reg1776 = $unsigned(reg1776[(3'h5):(1'h1)]);
              reg1777 = reg1743[(3'h6):(3'h4)];
              reg1778 <= $signed($signed(reg1668));
              reg1780 = ({($unsigned(((8'hbd) ? wire0 : (8'h9f))) ?
                      reg1731 : wire1),
                  (((wire0 ?
                      reg1759 : wire24) + $signed(reg353)) <= (~|(~reg1714)))} >> $unsigned((^{(&reg1761),
                  reg1718})));
            end
          reg1781 <= $signed($signed({$signed((reg1699 - (8'hb1)))}));
        end
      reg1782 = ((|$signed((|(+wire1)))) ?
          ($signed($unsigned((forvar1772 ?
              reg1720 : reg347))) >= {forvar1772[(2'h2):(1'h1)],
              reg1778[(2'h2):(1'h0)]}) : (reg1770[(4'he):(2'h2)] ^~ (($signed(reg1756) ?
              reg1698 : (-wire1)) == reg1697)));
      reg1783 <= (8'hb0);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module357
#(parameter param1629 = (+((|{((7'h46) ? (8'hb1) : (8'had))}) ? ((((8'hba) < (7'h45)) | ((8'ha6) ? (8'hba) : (7'h49))) > ((!(8'h9d)) * ((8'ha9) ? (8'ha3) : (7'h49)))) : ((-(8'ha2)) >> (((8'ha1) | (7'h4a)) < (7'h45))))), 
parameter param1630 = param1629)
(y, clk, wire358, wire359, wire360, wire361);
  output wire [(32'h976):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire358;
  input wire [(5'h18):(1'h0)] wire359;
  input wire signed [(3'h4):(1'h0)] wire360;
  input wire signed [(5'h14):(1'h0)] wire361;
  wire signed [(2'h2):(1'h0)] wire1628;
  wire [(3'h7):(1'h0)] wire1597;
  wire [(5'h12):(1'h0)] wire1596;
  wire [(3'h4):(1'h0)] wire1594;
  wire signed [(4'hb):(1'h0)] wire810;
  wire signed [(2'h2):(1'h0)] wire806;
  wire signed [(5'h14):(1'h0)] wire805;
  wire [(5'h13):(1'h0)] wire724;
  wire [(5'h13):(1'h0)] wire719;
  reg [(3'h5):(1'h0)] reg1626 = (1'h0);
  reg [(4'hc):(1'h0)] reg1625 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1612 = (1'h0);
  reg [(5'h14):(1'h0)] reg1610 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1606 = (1'h0);
  reg [(5'h13):(1'h0)] reg1622 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1621 = (1'h0);
  reg [(5'h18):(1'h0)] reg1620 = (1'h0);
  reg [(4'ha):(1'h0)] reg1616 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1615 = (1'h0);
  reg [(3'h7):(1'h0)] reg1611 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1609 = (1'h0);
  reg [(3'h7):(1'h0)] reg1608 = (1'h0);
  reg [(3'h6):(1'h0)] reg1607 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1603 = (1'h0);
  reg [(4'h8):(1'h0)] reg1600 = (1'h0);
  reg [(4'h8):(1'h0)] reg1599 = (1'h0);
  reg [(5'h17):(1'h0)] reg1598 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg851 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg844 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg850 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg849 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg848 = (1'h0);
  reg [(4'hf):(1'h0)] reg847 = (1'h0);
  reg [(2'h2):(1'h0)] reg843 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg841 = (1'h0);
  reg [(2'h3):(1'h0)] reg839 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg837 = (1'h0);
  reg [(5'h17):(1'h0)] reg834 = (1'h0);
  reg [(5'h15):(1'h0)] reg832 = (1'h0);
  reg [(4'h9):(1'h0)] reg831 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg826 = (1'h0);
  reg [(5'h13):(1'h0)] reg825 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg824 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg823 = (1'h0);
  reg [(3'h6):(1'h0)] reg821 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg820 = (1'h0);
  reg [(4'h9):(1'h0)] reg819 = (1'h0);
  reg [(3'h6):(1'h0)] reg818 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg817 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg816 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg813 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg809 = (1'h0);
  reg [(5'h15):(1'h0)] reg800 = (1'h0);
  reg [(5'h18):(1'h0)] reg796 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg804 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg803 = (1'h0);
  reg [(2'h3):(1'h0)] reg802 = (1'h0);
  reg [(4'hc):(1'h0)] reg801 = (1'h0);
  reg [(2'h2):(1'h0)] reg797 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg795 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg793 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg790 = (1'h0);
  reg [(5'h16):(1'h0)] reg788 = (1'h0);
  reg [(3'h6):(1'h0)] reg787 = (1'h0);
  reg [(5'h12):(1'h0)] reg786 = (1'h0);
  reg [(4'hc):(1'h0)] reg784 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg782 = (1'h0);
  reg [(4'hb):(1'h0)] reg778 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg774 = (1'h0);
  reg [(4'hc):(1'h0)] reg773 = (1'h0);
  reg [(5'h15):(1'h0)] reg772 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg771 = (1'h0);
  reg [(4'hf):(1'h0)] reg768 = (1'h0);
  reg [(5'h16):(1'h0)] reg767 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg763 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg762 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg760 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg758 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg757 = (1'h0);
  reg [(5'h18):(1'h0)] reg756 = (1'h0);
  reg [(4'hb):(1'h0)] reg754 = (1'h0);
  reg [(4'hd):(1'h0)] reg750 = (1'h0);
  reg [(5'h13):(1'h0)] reg749 = (1'h0);
  reg [(5'h16):(1'h0)] reg745 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg738 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg732 = (1'h0);
  reg [(5'h17):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg730 = (1'h0);
  reg [(4'h8):(1'h0)] reg728 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg723 = (1'h0);
  reg [(5'h11):(1'h0)] reg722 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg375 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg373 = (1'h0);
  reg [(4'h9):(1'h0)] reg371 = (1'h0);
  reg [(4'ha):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg366 = (1'h0);
  reg [(5'h10):(1'h0)] reg363 = (1'h0);
  reg [(4'hf):(1'h0)] reg1627 = (1'h0);
  reg [(5'h12):(1'h0)] reg1624 = (1'h0);
  reg [(2'h3):(1'h0)] reg1623 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1609 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1599 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1619 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1618 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1617 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1614 = (1'h0);
  reg [(4'h9):(1'h0)] reg1613 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1612 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1610 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1606 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1605 = (1'h0);
  reg [(4'hd):(1'h0)] reg1604 = (1'h0);
  reg [(5'h14):(1'h0)] reg1602 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1601 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar839 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg846 = (1'h0);
  reg [(5'h11):(1'h0)] reg845 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar844 = (1'h0);
  reg [(2'h2):(1'h0)] reg842 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg838 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg836 = (1'h0);
  reg [(4'h8):(1'h0)] reg835 = (1'h0);
  reg [(5'h18):(1'h0)] forvar833 = (1'h0);
  reg [(4'hc):(1'h0)] forvar827 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar830 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg829 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg828 = (1'h0);
  reg [(5'h11):(1'h0)] reg827 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar822 = (1'h0);
  reg [(2'h2):(1'h0)] reg815 = (1'h0);
  reg signed [(4'he):(1'h0)] reg814 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar812 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar811 = (1'h0);
  reg [(5'h18):(1'h0)] reg808 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg807 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar787 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar800 = (1'h0);
  reg [(4'hf):(1'h0)] reg799 = (1'h0);
  reg [(5'h14):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar796 = (1'h0);
  reg [(5'h18):(1'h0)] reg794 = (1'h0);
  reg [(5'h12):(1'h0)] reg792 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg791 = (1'h0);
  reg [(5'h18):(1'h0)] reg789 = (1'h0);
  reg [(4'hd):(1'h0)] reg785 = (1'h0);
  reg [(3'h6):(1'h0)] forvar783 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg781 = (1'h0);
  reg [(4'ha):(1'h0)] forvar780 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg779 = (1'h0);
  reg [(4'ha):(1'h0)] reg777 = (1'h0);
  reg [(2'h2):(1'h0)] forvar776 = (1'h0);
  reg [(4'ha):(1'h0)] reg775 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg770 = (1'h0);
  reg [(5'h15):(1'h0)] reg769 = (1'h0);
  reg [(5'h18):(1'h0)] forvar766 = (1'h0);
  reg [(3'h4):(1'h0)] reg765 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg764 = (1'h0);
  reg [(3'h7):(1'h0)] reg761 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar759 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg755 = (1'h0);
  reg [(3'h5):(1'h0)] forvar753 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg752 = (1'h0);
  reg [(3'h4):(1'h0)] reg751 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg748 = (1'h0);
  reg [(3'h6):(1'h0)] reg747 = (1'h0);
  reg [(3'h6):(1'h0)] reg746 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar744 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar743 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg742 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg741 = (1'h0);
  reg [(3'h7):(1'h0)] reg740 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar739 = (1'h0);
  reg [(2'h2):(1'h0)] reg737 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg736 = (1'h0);
  reg [(3'h5):(1'h0)] reg735 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg734 = (1'h0);
  reg [(2'h3):(1'h0)] reg733 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg729 = (1'h0);
  reg [(4'h8):(1'h0)] reg727 = (1'h0);
  reg [(5'h15):(1'h0)] forvar726 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar725 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg721 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg372 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg369 = (1'h0);
  reg signed [(4'he):(1'h0)] reg367 = (1'h0);
  reg [(4'ha):(1'h0)] forvar365 = (1'h0);
  reg [(4'hb):(1'h0)] reg364 = (1'h0);
  reg [(5'h14):(1'h0)] reg362 = (1'h0);
  assign y = {wire1628,
                 wire1597,
                 wire1596,
                 wire1594,
                 wire810,
                 wire806,
                 wire805,
                 wire724,
                 wire719,
                 reg1626,
                 reg1625,
                 reg1612,
                 reg1610,
                 reg1606,
                 reg1622,
                 reg1621,
                 reg1620,
                 reg1616,
                 reg1615,
                 reg1611,
                 reg1609,
                 reg1608,
                 reg1607,
                 reg1603,
                 reg1600,
                 reg1599,
                 reg1598,
                 reg851,
                 reg844,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 reg843,
                 reg841,
                 reg839,
                 reg837,
                 reg834,
                 reg832,
                 reg831,
                 reg826,
                 reg825,
                 reg824,
                 reg823,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 reg817,
                 reg816,
                 reg813,
                 reg809,
                 reg800,
                 reg796,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg797,
                 reg795,
                 reg793,
                 reg790,
                 reg788,
                 reg787,
                 reg786,
                 reg784,
                 reg782,
                 reg778,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg768,
                 reg767,
                 reg763,
                 reg762,
                 reg760,
                 reg758,
                 reg757,
                 reg756,
                 reg754,
                 reg750,
                 reg749,
                 reg745,
                 reg738,
                 reg732,
                 reg731,
                 reg730,
                 reg728,
                 reg723,
                 reg722,
                 reg375,
                 reg373,
                 reg371,
                 reg368,
                 reg366,
                 reg363,
                 reg1627,
                 reg1624,
                 reg1623,
                 forvar1609,
                 forvar1599,
                 reg1619,
                 reg1618,
                 reg1617,
                 reg1614,
                 reg1613,
                 forvar1612,
                 forvar1610,
                 forvar1606,
                 reg1605,
                 reg1604,
                 reg1602,
                 reg1601,
                 forvar839,
                 reg846,
                 reg845,
                 forvar844,
                 reg842,
                 reg840,
                 reg838,
                 reg836,
                 reg835,
                 forvar833,
                 forvar827,
                 forvar830,
                 reg829,
                 reg828,
                 reg827,
                 forvar822,
                 reg815,
                 reg814,
                 forvar812,
                 forvar811,
                 reg808,
                 reg807,
                 forvar787,
                 forvar800,
                 reg799,
                 reg798,
                 forvar796,
                 reg794,
                 reg792,
                 reg791,
                 reg789,
                 reg785,
                 forvar783,
                 reg781,
                 forvar780,
                 reg779,
                 reg777,
                 forvar776,
                 reg775,
                 reg770,
                 reg769,
                 forvar766,
                 reg765,
                 reg764,
                 reg761,
                 forvar759,
                 reg755,
                 forvar753,
                 reg752,
                 reg751,
                 reg748,
                 reg747,
                 reg746,
                 forvar744,
                 forvar743,
                 reg742,
                 reg741,
                 reg740,
                 forvar739,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg729,
                 reg727,
                 forvar726,
                 forvar725,
                 reg721,
                 reg374,
                 reg372,
                 reg370,
                 reg369,
                 reg367,
                 forvar365,
                 reg364,
                 reg362,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg362 = {(wire358[(2'h3):(1'h0)] ?
              ($unsigned({wire358}) || wire359) : (($unsigned(wire359) - wire359[(4'h8):(2'h3)]) || (~wire359[(3'h5):(3'h4)])))};
      reg363 <= (reg362[(5'h14):(5'h14)] <<< ((8'ha6) != wire360));
      reg364 = $unsigned((~(wire360[(2'h2):(1'h1)] ?
          (!((8'h9e) ~^ (8'h9d))) : reg362[(4'h8):(3'h6)])));
      for (forvar365 = (1'h0); (forvar365 < (1'h0)); forvar365 = (forvar365 + (1'h1)))
        begin
          reg366 <= wire358;
          if (((($signed(wire358[(4'ha):(4'h9)]) || $signed(reg363)) >>> (($unsigned(reg362) ?
                      forvar365 : wire361) ?
                  reg366 : (^(reg362 <= wire360)))) ?
              (reg362[(5'h12):(4'h9)] - reg364) : (8'hbb)))
            begin
              reg367 = reg362;
              reg368 <= reg366[(2'h2):(1'h0)];
              reg369 = wire358[(2'h3):(1'h0)];
              reg370 = ($signed((~^$unsigned(reg367[(2'h2):(2'h2)]))) ?
                  (((^$unsigned(reg362)) << {(wire358 ? reg363 : reg366),
                      (&reg368)}) * reg367[(1'h1):(1'h0)]) : wire361[(4'hb):(2'h3)]);
              reg371 <= {{($signed({(8'hae)}) - (|wire359))},
                  (|reg370[(4'hc):(2'h2)])};
            end
          else
            begin
              reg367 = $unsigned((!((+(reg370 < reg364)) | reg368[(2'h3):(1'h1)])));
              reg369 = reg363[(5'h10):(3'h6)];
              reg371 <= $unsigned(reg371[(1'h1):(1'h1)]);
              reg372 = {{((forvar365[(4'h8):(4'h8)] < reg369[(4'hd):(3'h4)]) != $signed((wire360 ?
                          reg371 : reg368)))},
                  ((8'ha3) * reg367)};
              reg373 <= ({reg368[(3'h6):(2'h3)]} ^ ($signed(reg367[(4'h8):(3'h7)]) <<< wire359[(4'h8):(1'h0)]));
            end
          reg374 = $unsigned($unsigned((-wire361)));
          reg375 <= (|(8'ha6));
        end
    end
  module376 #() modinst720 (.wire380(wire361), .y(wire719), .clk(clk), .wire381(reg363), .wire379(wire358), .wire377(wire359), .wire378(reg366));
  always
    @(posedge clk) begin
      reg721 = reg366[(4'he):(4'h9)];
      reg722 <= $unsigned({$signed(($unsigned(reg363) ?
              (reg721 >>> wire719) : (~&(7'h44)))),
          (~|(+$signed(wire359)))});
      reg723 <= reg721[(3'h4):(2'h2)];
    end
  assign wire724 = $signed($signed(wire358[(4'ha):(4'h9)]));
  always
    @(posedge clk) begin
      for (forvar725 = (1'h0); (forvar725 < (1'h1)); forvar725 = (forvar725 + (1'h1)))
        begin
          for (forvar726 = (1'h0); (forvar726 < (2'h2)); forvar726 = (forvar726 + (1'h1)))
            begin
              reg727 = forvar726;
            end
          if ((-(forvar725 ?
              ($unsigned(wire358[(3'h7):(3'h5)]) ?
                  $signed((+forvar726)) : ($unsigned(reg375) >= {(8'hbe)})) : reg366[(5'h13):(4'hc)])))
            begin
              reg728 <= {((7'h47) ?
                      reg722 : $unsigned(((reg366 ?
                          wire358 : reg363) >>> (reg723 + reg366)))),
                  $signed((8'hb9))};
            end
          else
            begin
              reg728 <= reg375;
            end
          reg729 = ($unsigned(({(8'ha0)} >= (8'ha8))) + reg727);
        end
      if ((~$unsigned(reg722)))
        begin
          if (($unsigned({wire358[(3'h4):(2'h2)], $unsigned((-reg375))}) ?
              reg375 : {((&(wire359 ? (8'hb6) : (8'hbc))) ?
                      (forvar725 >>> (reg371 ~^ reg366)) : ($signed(reg363) ?
                          (reg368 != wire359) : (reg722 == (8'hb7)))),
                  $signed(($signed(reg727) ? {reg373} : $unsigned(reg368)))}))
            begin
              reg730 <= ($unsigned(forvar726) ?
                  $unsigned({reg723}) : $unsigned((($signed(wire719) ?
                      {reg722} : $unsigned((8'ha0))) != reg366)));
              reg731 <= {(reg371 ^~ (&wire360)),
                  ($signed($unsigned(((8'hb4) ?
                      reg373 : (8'had)))) <= (&((~&reg722) ?
                      (reg371 < wire358) : {reg729})))};
              reg732 <= reg371[(1'h0):(1'h0)];
            end
          else
            begin
              reg733 = ((-$signed((!$signed((7'h48))))) ?
                  $signed($unsigned((((7'h46) << reg363) >= (reg731 - wire359)))) : reg731);
              reg734 = reg730;
              reg735 = {($signed(((reg731 ?
                      forvar725 : (8'hbc)) ~^ {wire359})) & (((~^wire359) ?
                      $signed(reg727) : $unsigned(wire724)) > reg366[(2'h3):(2'h2)])),
                  (reg368 ? reg731[(1'h0):(1'h0)] : reg371)};
              reg736 = (reg375 + $signed($unsigned($signed((reg729 + (8'hb2))))));
              reg737 = reg735;
            end
          reg738 <= wire719[(1'h0):(1'h0)];
          for (forvar739 = (1'h0); (forvar739 < (1'h0)); forvar739 = (forvar739 + (1'h1)))
            begin
              reg740 = (^~(!$unsigned(((8'hba) ?
                  $signed(reg737) : $unsigned(reg731)))));
              reg741 = (~|{(~$unsigned(wire360[(1'h0):(1'h0)]))});
              reg742 = reg732;
            end
        end
      else
        begin
          reg730 <= reg373;
          if ((reg729[(4'h9):(3'h5)] ? reg729 : reg722))
            begin
              reg731 <= wire360[(1'h1):(1'h0)];
              reg733 = (-$signed((&reg730[(3'h4):(2'h2)])));
              reg734 = ($unsigned($unsigned(($unsigned(reg371) * $unsigned(wire359)))) ?
                  ((forvar739 <= $unsigned($signed(reg368))) <= (^reg368[(2'h2):(1'h0)])) : (wire358[(4'hd):(1'h0)] <= ($signed($unsigned(reg729)) ?
                      (^reg373) : (~|(~&reg731)))));
            end
          else
            begin
              reg733 = (!(!$signed($signed($signed(wire724)))));
              reg734 = (&reg373[(4'h9):(2'h2)]);
            end
        end
      for (forvar743 = (1'h0); (forvar743 < (1'h0)); forvar743 = (forvar743 + (1'h1)))
        begin
          for (forvar744 = (1'h0); (forvar744 < (1'h1)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 <= $signed((|reg723));
              reg746 = (^~forvar726[(2'h3):(2'h3)]);
              reg747 = (^~wire719[(4'hb):(3'h5)]);
            end
          if ($signed((~^$signed(reg737[(2'h2):(2'h2)]))))
            begin
              reg748 = $unsigned(((!$unsigned($signed(reg738))) ~^ (({(8'hba),
                  reg728} | $unsigned(reg741)) ^~ $unsigned((reg375 ?
                  forvar725 : forvar726)))));
            end
          else
            begin
              reg749 <= (-(reg366[(2'h2):(2'h2)] ?
                  reg738[(1'h1):(1'h1)] : ((^~$unsigned(reg735)) * (reg727[(4'h8):(1'h0)] ?
                      wire724 : $signed(reg730)))));
              reg750 <= (~&reg730);
              reg751 = $unsigned(reg730[(5'h13):(1'h0)]);
              reg752 = ($unsigned((forvar744 ^~ (~|$unsigned(reg723)))) ?
                  $signed(((+wire358) ?
                      {$unsigned(reg748)} : reg731)) : (reg728 + reg375));
            end
          for (forvar753 = (1'h0); (forvar753 < (3'h4)); forvar753 = (forvar753 + (1'h1)))
            begin
              reg754 <= {$signed(((^$signed((8'hba))) ?
                      ($unsigned((8'hbe)) ?
                          (reg732 ?
                              reg375 : reg734) : reg735[(1'h1):(1'h1)]) : {$unsigned(reg731),
                          $unsigned(reg722)}))};
            end
          reg755 = (~$unsigned($signed({(reg741 ? wire719 : reg729)})));
        end
      if ((|reg728))
        begin
          reg756 <= {((~$unsigned((~reg736))) ?
                  (~^reg742[(1'h1):(1'h0)]) : ((-wire360[(3'h4):(1'h1)]) ?
                      {(-reg732),
                          reg735} : ($unsigned(wire358) + (^~reg747))))};
        end
      else
        begin
          reg756 <= reg754[(4'hb):(3'h6)];
          reg757 <= $signed($signed({($signed(reg366) - $unsigned(reg749))}));
          reg758 <= ((-forvar726[(4'hc):(4'h8)]) ^~ reg741);
          for (forvar759 = (1'h0); (forvar759 < (2'h3)); forvar759 = (forvar759 + (1'h1)))
            begin
              reg760 <= (~&$unsigned((forvar744 >> $signed(forvar744))));
              reg761 = (&((($unsigned(forvar739) ~^ reg375) & ($unsigned(reg368) ?
                  wire359 : reg733[(2'h2):(2'h2)])) != (^~reg740[(1'h1):(1'h1)])));
              reg762 <= $signed(forvar753);
              reg763 <= reg375[(2'h3):(2'h3)];
            end
        end
      reg764 = (7'h49);
    end
  always
    @(posedge clk) begin
      reg765 = reg738[(1'h1):(1'h1)];
      for (forvar766 = (1'h0); (forvar766 < (2'h3)); forvar766 = (forvar766 + (1'h1)))
        begin
          if (({({(~^reg731), reg363} ? reg757 : (~&(reg758 << reg757))),
                  $unsigned(reg722[(1'h1):(1'h0)])} ?
              (!reg758) : reg375[(3'h6):(1'h1)]))
            begin
              reg767 <= $signed((((reg750[(3'h7):(2'h3)] ?
                          $unsigned(reg757) : $signed(reg363)) ?
                      (reg722[(4'hd):(3'h5)] != $unsigned((7'h45))) : reg730) ?
                  (reg371 == reg758[(3'h4):(2'h3)]) : (7'h48)));
              reg768 <= $unsigned(reg765[(1'h1):(1'h0)]);
              reg769 = reg757[(4'hc):(4'h9)];
              reg770 = $signed({((~^reg760[(4'hb):(1'h0)]) ?
                      ($signed(reg750) & $unsigned((8'h9e))) : (~^(~|wire719))),
                  (^{(reg723 ? reg731 : reg375), reg762[(4'h8):(4'h8)]})});
            end
          else
            begin
              reg769 = reg723[(4'ha):(4'ha)];
              reg771 <= reg730[(2'h2):(1'h1)];
              reg772 <= (7'h48);
            end
          reg773 <= reg763;
          reg774 <= ($signed((($unsigned(wire724) ?
              (~^reg770) : $signed(reg765)) < forvar766[(3'h7):(3'h7)])) <<< reg762);
          reg775 = ((wire361 ? $unsigned(reg745) : reg750[(4'hc):(4'h8)]) ?
              reg763 : wire724[(4'he):(1'h1)]);
        end
      for (forvar776 = (1'h0); (forvar776 < (1'h1)); forvar776 = (forvar776 + (1'h1)))
        begin
          reg777 = forvar776;
          if ({reg728[(3'h7):(1'h0)], reg730[(1'h1):(1'h0)]})
            begin
              reg778 <= ((^reg749) || $signed((~reg732[(1'h0):(1'h0)])));
            end
          else
            begin
              reg778 <= reg756;
              reg779 = (&reg778);
            end
          for (forvar780 = (1'h0); (forvar780 < (2'h2)); forvar780 = (forvar780 + (1'h1)))
            begin
              reg781 = $signed((reg723[(4'h8):(2'h3)] ?
                  (&$unsigned((reg723 + forvar780))) : reg732));
              reg782 <= (~&reg769);
            end
          for (forvar783 = (1'h0); (forvar783 < (2'h3)); forvar783 = (forvar783 + (1'h1)))
            begin
              reg784 <= (!(~|$signed($signed(forvar783))));
              reg785 = $unsigned((($unsigned((reg774 <<< reg750)) | (^~reg763)) ^ ($unsigned((^reg366)) ?
                  $signed(wire361[(1'h0):(1'h0)]) : ((wire724 ?
                          forvar776 : reg777) ?
                      {(8'hb9)} : $unsigned(wire361)))));
            end
          reg786 <= {(^~($unsigned((7'h40)) == (~reg728[(3'h7):(2'h2)]))),
              (((reg773[(3'h6):(2'h3)] ? {wire361} : (reg765 && reg723)) ?
                  forvar780[(2'h2):(1'h1)] : ($unsigned((8'hb7)) >= {reg760,
                      (8'ha3)})) <<< reg773[(2'h3):(1'h0)])};
        end
      if ($signed((^~reg785)))
        begin
          if (wire719[(5'h10):(4'hd)])
            begin
              reg787 <= $signed(reg738);
              reg788 <= $unsigned((~({(reg363 ? forvar766 : reg760),
                      reg722[(2'h3):(2'h3)]} ?
                  ($signed(reg371) >> reg773) : reg762)));
              reg789 = ($signed((reg785[(2'h3):(2'h2)] * $signed((reg778 ?
                      (7'h48) : reg754)))) ?
                  ({{$signed(reg732)}} ?
                      wire358 : (~&(&(reg732 ?
                          reg778 : wire719)))) : $signed(reg779));
              reg790 <= reg775[(1'h1):(1'h0)];
              reg791 = (~$unsigned($unsigned(({wire360} <<< (reg790 ?
                  reg723 : reg760)))));
            end
          else
            begin
              reg787 <= reg782[(3'h7):(3'h5)];
              reg789 = (^~wire360[(1'h1):(1'h1)]);
              reg791 = {(+(&$unsigned($signed(wire724)))),
                  (&forvar783[(1'h1):(1'h0)])};
              reg792 = reg767;
              reg793 <= reg722;
            end
          if ($signed($signed(((8'hb8) < ($unsigned(wire724) ?
              $unsigned(reg771) : reg731[(2'h2):(2'h2)])))))
            begin
              reg794 = reg373;
              reg795 <= $unsigned(((!$unsigned(reg760)) ?
                  (reg782 * $signed(((8'ha8) || reg732))) : reg790[(2'h3):(2'h2)]));
            end
          else
            begin
              reg795 <= (((8'ha2) ?
                  $unsigned(wire360) : (((^reg762) ^ (!reg795)) ?
                      reg373 : (8'ha6))) >>> (-reg773));
            end
          for (forvar796 = (1'h0); (forvar796 < (2'h2)); forvar796 = (forvar796 + (1'h1)))
            begin
              reg797 <= $unsigned(reg775);
              reg798 = ($unsigned(reg375) + reg771);
              reg799 = (-$signed({(-$signed((8'haa))),
                  ((reg789 ? reg763 : reg760) ?
                      (~reg795) : $unsigned(reg756))}));
            end
          for (forvar800 = (1'h0); (forvar800 < (2'h3)); forvar800 = (forvar800 + (1'h1)))
            begin
              reg801 <= (|((reg777[(2'h2):(1'h0)] || reg799) ?
                  ((wire719 && (forvar796 ^ (8'hb5))) ?
                      ((reg765 ~^ wire359) ?
                          (reg788 ?
                              reg771 : reg728) : $unsigned(reg767)) : reg788[(5'h15):(1'h0)]) : {(8'hb0),
                      $signed($unsigned(reg760))}));
              reg802 <= reg769[(4'hc):(4'hc)];
              reg803 <= (reg730[(4'ha):(3'h5)] ?
                  (~((reg732 - reg750) ?
                      ($signed(reg786) & {forvar776,
                          reg792}) : $unsigned((~|(8'ha3))))) : (!($unsigned($signed(reg792)) > $unsigned(wire358[(4'h9):(3'h7)]))));
              reg804 <= (reg803[(1'h0):(1'h0)] ?
                  reg794[(5'h11):(4'hf)] : {(($signed((7'h42)) + (wire724 ?
                              reg784 : reg765)) ?
                          $unsigned(wire724[(4'h9):(1'h1)]) : {(reg784 ?
                                  (8'hbd) : reg757)})});
            end
        end
      else
        begin
          for (forvar787 = (1'h0); (forvar787 < (2'h3)); forvar787 = (forvar787 + (1'h1)))
            begin
              reg789 = (+$unsigned((~&$unsigned(reg786))));
              reg791 = (8'haa);
              reg793 <= {forvar766[(5'h18):(3'h6)]};
            end
          reg795 <= (reg774 ?
              forvar780 : $unsigned((+{reg781[(1'h1):(1'h1)]})));
          if (((reg730 - $signed($unsigned(reg781[(2'h3):(2'h2)]))) ^ {{((reg771 ?
                      (7'h44) : wire724) ^ (~reg799))}}))
            begin
              reg796 <= $signed(((((8'hb2) ?
                      $signed(reg771) : reg782[(2'h2):(2'h2)]) ?
                  $unsigned({reg728,
                      wire719}) : reg368) >= forvar800[(2'h3):(1'h1)]));
              reg797 <= reg799[(3'h4):(3'h4)];
              reg798 = $unsigned(((~|(^~(reg796 ^~ (7'h40)))) ?
                  wire719[(4'h8):(1'h0)] : $signed($unsigned((reg786 ^ reg375)))));
              reg799 = reg769;
              reg800 <= $unsigned(($signed((8'ha3)) | reg790));
            end
          else
            begin
              reg796 <= reg363;
            end
        end
    end
  assign wire805 = reg773;
  assign wire806 = $signed((+($unsigned($unsigned(reg793)) ?
                       (reg363[(4'hb):(3'h7)] < $unsigned((8'hb2))) : {reg786[(4'hd):(1'h0)],
                           ((8'hbf) >>> reg801)})));
  always
    @(posedge clk) begin
      reg807 = (reg723[(4'hd):(3'h7)] | {reg750});
      reg808 = {reg375};
      reg809 <= (~&$unsigned((reg732 || $signed(((7'h40) > reg795)))));
    end
  assign wire810 = wire806;
  always
    @(posedge clk) begin
      for (forvar811 = (1'h0); (forvar811 < (2'h3)); forvar811 = (forvar811 + (1'h1)))
        begin
          for (forvar812 = (1'h0); (forvar812 < (2'h2)); forvar812 = (forvar812 + (1'h1)))
            begin
              reg813 <= $signed(reg762[(3'h4):(2'h3)]);
              reg814 = ((reg796[(4'hb):(4'ha)] != wire360[(2'h3):(1'h0)]) - ({(^~wire810),
                  reg373[(3'h5):(3'h5)]} <<< (^~(reg762 ?
                  reg757 : {(7'h48)}))));
              reg815 = (wire359[(5'h11):(4'hd)] ?
                  reg728[(1'h0):(1'h0)] : reg767[(5'h14):(3'h4)]);
              reg816 <= ({({$signed(reg772)} ?
                      reg763[(1'h1):(1'h0)] : (reg771 << reg802))} + (^~$signed(((reg756 >= wire724) ?
                  ((8'ha3) ? reg757 : reg757) : $unsigned(reg762)))));
              reg817 <= (^~(!$unsigned(reg760)));
            end
          reg818 <= $unsigned({reg368[(4'h8):(3'h6)]});
          if ($unsigned(($signed((!(wire361 | (8'hae)))) ?
              (reg375 ?
                  (+(reg778 < reg749)) : (((8'hae) ?
                      (8'h9d) : reg723) >= reg817)) : (reg788 & reg788))))
            begin
              reg819 <= reg800;
              reg820 <= reg758[(5'h16):(1'h0)];
              reg821 <= (^wire360[(3'h4):(1'h0)]);
            end
          else
            begin
              reg819 <= {((~|reg760) ?
                      {(~(+wire358)), reg732[(1'h1):(1'h1)]} : (~((forvar811 ?
                          wire361 : wire724) << $unsigned(reg818)))),
                  reg821};
              reg820 <= {reg722[(5'h11):(2'h2)],
                  (((^~(^~wire361)) && $unsigned((wire805 ~^ reg738))) ?
                      ($signed((8'ha2)) ?
                          $signed(reg813[(3'h5):(2'h3)]) : reg814) : $unsigned($unsigned(forvar811)))};
              reg821 <= $signed((~|($unsigned((~&reg802)) ^ ($signed(reg790) >> (reg790 ^~ wire361)))));
            end
          for (forvar822 = (1'h0); (forvar822 < (1'h1)); forvar822 = (forvar822 + (1'h1)))
            begin
              reg823 <= (!{reg796});
              reg824 <= $signed(($unsigned((~^(reg750 ? reg731 : reg754))) ?
                  (-((^reg778) + (!reg796))) : wire360[(1'h1):(1'h1)]));
              reg825 <= (&$signed({$signed($signed(reg772)),
                  ($signed((7'h46)) < reg772)}));
              reg826 <= (!$signed({reg371[(2'h3):(2'h3)],
                  $unsigned((reg750 + wire360))}));
            end
        end
      if (reg819)
        begin
          reg827 = (-$signed((reg793[(4'h8):(4'h8)] ~^ reg760)));
          reg828 = (wire810 ?
              reg363[(3'h6):(2'h2)] : $signed($signed(reg817[(3'h4):(1'h0)])));
          reg829 = reg787[(3'h6):(3'h4)];
          for (forvar830 = (1'h0); (forvar830 < (2'h3)); forvar830 = (forvar830 + (1'h1)))
            begin
              reg831 <= reg802;
              reg832 <= {$signed($unsigned((reg829[(3'h4):(1'h1)] & reg828[(1'h1):(1'h0)])))};
            end
        end
      else
        begin
          for (forvar827 = (1'h0); (forvar827 < (3'h4)); forvar827 = (forvar827 + (1'h1)))
            begin
              reg828 = $signed((((~reg771[(4'h8):(3'h6)]) > ((reg790 ?
                          reg363 : wire805) ?
                      $signed(reg732) : reg375[(3'h5):(3'h5)])) ?
                  ($signed((reg820 ?
                      reg782 : reg793)) <<< reg763) : $unsigned(($unsigned(reg795) >> $signed(reg821)))));
            end
          reg829 = $unsigned(wire358);
          for (forvar830 = (1'h0); (forvar830 < (2'h3)); forvar830 = (forvar830 + (1'h1)))
            begin
              reg831 <= $unsigned({(8'hbc)});
              reg832 <= ((-(reg784[(3'h5):(2'h2)] ~^ (8'hbb))) ~^ (reg778[(4'hb):(3'h6)] ?
                  $unsigned(wire719) : (reg829 ?
                      reg373 : ((~^forvar811) ?
                          (reg821 * reg754) : forvar812[(2'h2):(2'h2)]))));
            end
          for (forvar833 = (1'h0); (forvar833 < (2'h2)); forvar833 = (forvar833 + (1'h1)))
            begin
              reg834 <= (8'haf);
              reg835 = reg804;
              reg836 = {({($signed(reg804) ?
                          $signed(reg756) : $unsigned(reg366))} ^~ forvar827)};
              reg837 <= {{{(!$unsigned(reg786))}, $unsigned((!(^reg757)))}};
            end
        end
      reg838 = reg757[(4'he):(1'h0)];
    end
  always
    @(posedge clk) begin
      if ((((^$signed(reg802)) <= {reg788, (~&reg826)}) ?
          (|(reg738 * reg749[(3'h5):(1'h1)])) : reg730[(5'h13):(4'he)]))
        begin
          if ($signed($unsigned((reg750[(3'h5):(3'h4)] ~^ $signed($unsigned(reg823))))))
            begin
              reg839 <= $unsigned(reg797);
              reg840 = {{($unsigned(reg763[(2'h2):(1'h0)]) ?
                          reg738[(1'h0):(1'h0)] : ((-wire360) == (~&(8'hbd))))},
                  reg825};
              reg841 <= $signed((~&(^~(8'haf))));
              reg842 = reg793[(4'hc):(4'ha)];
            end
          else
            begin
              reg840 = (reg758 || (^($signed({reg837,
                  wire806}) ^~ $signed((+reg818)))));
            end
          reg843 <= reg772;
          for (forvar844 = (1'h0); (forvar844 < (1'h0)); forvar844 = (forvar844 + (1'h1)))
            begin
              reg845 = {(({{reg731, wire358}, ((8'ha8) ? reg731 : (8'hbe))} ?
                          (wire805[(4'he):(4'h9)] ?
                              (reg762 ?
                                  reg756 : reg839) : $signed(reg831)) : reg723[(3'h4):(2'h2)]) ?
                      reg749 : reg757)};
              reg846 = reg728;
              reg847 <= {$unsigned({$signed((reg768 ? reg800 : reg823))})};
              reg848 <= $signed((~^(8'hb0)));
            end
          reg849 <= reg797[(1'h1):(1'h1)];
          reg850 <= (((((reg837 ? (8'ha4) : reg797) ?
                      reg825[(3'h5):(2'h3)] : (reg817 == reg366)) ?
                  reg802 : ({reg757} | (reg768 ^~ reg839))) * reg749[(1'h1):(1'h1)]) ?
              ($unsigned($signed(reg796)) & $unsigned($signed((reg793 + reg371)))) : {(wire806[(1'h0):(1'h0)] - reg821)});
        end
      else
        begin
          for (forvar839 = (1'h0); (forvar839 < (1'h1)); forvar839 = (forvar839 + (1'h1)))
            begin
              reg840 = reg832;
              reg842 = {$signed({((reg788 <<< reg771) | $unsigned((8'hb9))),
                      reg738[(1'h0):(1'h0)]})};
              reg843 <= ($unsigned((({wire360, wire358} ?
                      reg831[(4'h8):(2'h3)] : (reg823 >= reg771)) || $unsigned($unsigned(reg787)))) ?
                  {reg754[(4'ha):(3'h4)],
                      ((-reg758) ~^ wire806)} : reg837[(1'h1):(1'h0)]);
              reg844 <= $signed(reg837);
              reg847 <= wire719;
            end
          reg848 <= ($unsigned($signed($signed((reg760 ^ reg758)))) >> reg793[(1'h0):(1'h0)]);
        end
      reg851 <= $signed((8'hb2));
    end
  module852 #() modinst1595 (wire1594, clk, reg788, reg824, reg731, reg837);
  assign wire1596 = ((($signed($unsigned(reg768)) ?
                            (reg732 & (reg787 + reg731)) : (~{reg790})) ?
                        (((|reg728) ?
                                ((8'hb2) ? (7'h46) : reg782) : (reg843 ?
                                    reg850 : (8'hb6))) ?
                            reg788 : (!(!reg821))) : reg824) >> (+reg749[(5'h13):(1'h0)]));
  assign wire1597 = wire805;
  always
    @(posedge clk) begin
      reg1598 <= ((!$signed($signed(reg848[(3'h4):(2'h3)]))) < {reg818[(3'h4):(1'h1)]});
    end
  always
    @(posedge clk) begin
      if (wire724)
        begin
          if (((($unsigned((reg758 ? reg804 : reg722)) + ({reg803} ?
                  (reg767 <= reg373) : (reg795 << reg760))) ?
              (~|{reg745[(3'h4):(3'h4)]}) : ((~$signed(reg809)) ^ $unsigned((~&reg768)))) <<< (8'hbe)))
            begin
              reg1599 <= ({wire805[(1'h1):(1'h0)]} ?
                  (^~((^reg722[(1'h1):(1'h1)]) < $unsigned(reg728[(2'h3):(2'h3)]))) : $signed({((wire805 < reg802) ?
                          {reg371} : {reg763})}));
              reg1600 <= (~|reg819[(3'h4):(1'h0)]);
              reg1601 = (&(8'hbe));
              reg1602 = (8'haf);
              reg1603 <= $unsigned(($signed(reg820[(5'h13):(5'h12)]) != $signed(((wire724 << reg730) ~^ reg813))));
            end
          else
            begin
              reg1601 = wire1597[(3'h6):(3'h4)];
              reg1603 <= $unsigned((|(~($signed(reg1598) ^~ (8'hbe)))));
              reg1604 = $signed(reg837);
              reg1605 = ($unsigned(((&$unsigned(reg773)) ^~ reg750)) ?
                  wire806 : (~reg731));
            end
          for (forvar1606 = (1'h0); (forvar1606 < (2'h3)); forvar1606 = (forvar1606 + (1'h1)))
            begin
              reg1607 <= reg1604[(2'h2):(1'h0)];
              reg1608 <= $unsigned(wire806[(2'h2):(1'h1)]);
              reg1609 <= $unsigned({($unsigned((reg371 - (7'h41))) ?
                      $signed((reg797 ^~ (7'h42))) : $unsigned((!reg841)))});
            end
          for (forvar1610 = (1'h0); (forvar1610 < (1'h0)); forvar1610 = (forvar1610 + (1'h1)))
            begin
              reg1611 <= ((($signed({reg1603}) <<< reg844) ?
                  (((reg786 ? reg848 : wire1597) ?
                          reg816[(1'h0):(1'h0)] : (-(8'ha4))) ?
                      reg795[(2'h2):(2'h2)] : (~^reg826[(1'h0):(1'h0)])) : wire361[(3'h6):(3'h5)]) <<< $unsigned(reg768));
            end
          for (forvar1612 = (1'h0); (forvar1612 < (2'h2)); forvar1612 = (forvar1612 + (1'h1)))
            begin
              reg1613 = reg738;
              reg1614 = $signed((~^reg826));
              reg1615 <= (+({(^(~(7'h43))),
                  $signed(reg801)} ^~ $unsigned(({(8'hbf)} ?
                  (reg1607 > reg820) : reg1605[(1'h1):(1'h0)]))));
              reg1616 <= reg793[(2'h3):(2'h3)];
              reg1617 = reg839[(1'h1):(1'h1)];
            end
          if ($unsigned((((7'h40) - $unsigned({reg760, reg848})) ?
              (reg773 << $unsigned((reg1607 ^ reg1598))) : ($signed(wire359) <= (+(reg757 - wire1596))))))
            begin
              reg1618 = forvar1612[(3'h4):(2'h2)];
              reg1619 = reg1614[(3'h6):(3'h5)];
            end
          else
            begin
              reg1620 <= ({$unsigned({reg773, $unsigned((7'h41))})} ?
                  $unsigned(((forvar1610[(3'h4):(1'h1)] ? reg1602 : wire361) ?
                      ((reg832 ^ reg774) ?
                          {reg844,
                              reg366} : (reg754 + (8'hbc))) : $signed((8'hb8)))) : ($unsigned(($unsigned(wire360) <<< (+forvar1606))) != reg774[(3'h7):(2'h3)]));
              reg1621 <= reg825;
              reg1622 <= (|{(8'hb2)});
            end
        end
      else
        begin
          for (forvar1599 = (1'h0); (forvar1599 < (2'h2)); forvar1599 = (forvar1599 + (1'h1)))
            begin
              reg1600 <= ((((reg839[(2'h2):(2'h2)] ?
                      reg768 : $unsigned(reg772)) | reg363[(5'h10):(3'h5)]) ?
                  wire1594 : ((reg851[(3'h4):(1'h0)] ?
                          $signed(reg837) : reg847) ?
                      $signed($unsigned(reg844)) : wire719[(4'ha):(1'h0)])) ~^ reg368[(3'h7):(1'h0)]);
              reg1603 <= (&reg851);
              reg1606 <= {(~|$unsigned((reg774 ?
                      reg749[(5'h13):(5'h10)] : $unsigned(reg825)))),
                  wire806[(1'h1):(1'h1)]};
              reg1607 <= reg851;
              reg1608 <= (8'hb1);
            end
          for (forvar1609 = (1'h0); (forvar1609 < (2'h3)); forvar1609 = (forvar1609 + (1'h1)))
            begin
              reg1610 <= ($signed(reg1600[(3'h7):(1'h0)]) + reg757[(1'h0):(1'h0)]);
              reg1611 <= reg1618;
              reg1612 <= {(+$unsigned(reg782))};
              reg1613 = reg820;
            end
          reg1615 <= {(8'hb8)};
          if (((~&{({(8'ha8), reg826} > {reg790, reg787}),
              (8'hb7)}) && $unsigned(($signed(wire358) ?
              reg1612 : {{reg1608}, (reg728 ? reg1618 : reg839)}))))
            begin
              reg1616 <= $unsigned((reg1598[(5'h10):(3'h4)] ?
                  $signed(reg1603) : (&(wire1596 ?
                      (reg837 <= reg1614) : $signed(reg1603)))));
            end
          else
            begin
              reg1616 <= $signed(reg821[(2'h2):(2'h2)]);
              reg1620 <= $unsigned((((+$signed(reg800)) <= ($unsigned(reg839) ?
                      (wire359 && reg821) : reg801[(3'h6):(1'h1)])) ?
                  (reg1602 > $signed($signed((8'h9d)))) : reg768[(4'h9):(4'h8)]));
            end
          if ($signed(reg723[(3'h7):(2'h2)]))
            begin
              reg1623 = reg1622[(2'h2):(1'h0)];
              reg1624 = {$unsigned(forvar1599[(4'h9):(4'h8)]),
                  $unsigned($signed((8'h9c)))};
              reg1625 <= {$signed((reg824 ^ (7'h43))), reg1608};
              reg1626 <= ({((~|reg774) ^~ $signed(reg773[(2'h3):(1'h0)]))} ?
                  reg1610[(5'h10):(4'he)] : (&{(reg790[(1'h0):(1'h0)] << (reg847 || wire805))}));
              reg1627 = $signed($signed(((!(reg1624 - (7'h41))) > ($signed(reg1598) >= $signed(reg824)))));
            end
          else
            begin
              reg1623 = (!((~^reg1603[(1'h0):(1'h0)]) <<< ($unsigned(reg824[(4'hb):(2'h2)]) >>> (!reg824))));
              reg1624 = (reg1604[(2'h3):(1'h0)] > {reg849[(4'hc):(4'h9)],
                  reg1609});
            end
        end
    end
  assign wire1628 = ($unsigned($signed((reg821[(2'h2):(2'h2)] ?
                        $unsigned((8'hba)) : $signed(reg774)))) < $unsigned(reg841));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module25
#(parameter param335 = (~^(((((8'hb0) ? (8'ha0) : (7'h49)) ? (~&(8'ha0)) : {(8'h9f), (8'ha6)}) ? (((8'ha8) & (8'ha3)) && {(8'hb6), (8'hbf)}) : (7'h41)) ? {{(-(8'had))}, (((8'h9f) ? (7'h45) : (8'h9c)) ? {(8'ha6)} : (^~(8'hba)))} : ((((8'hb1) ? (7'h40) : (7'h4a)) ? ((7'h4a) ? (8'ha9) : (8'ha2)) : ((8'ha9) ? (8'ha0) : (8'haf))) ? {(^(8'hb8)), ((8'ha5) || (8'hae))} : ((~(8'hbf)) || ((8'haa) ? (8'h9e) : (8'h9c)))))), 
parameter param336 = (!param335))
(y, clk, wire29, wire28, wire27, wire26);
  output wire [(32'hb4b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire29;
  input wire signed [(4'h8):(1'h0)] wire28;
  input wire [(4'ha):(1'h0)] wire27;
  input wire [(5'h10):(1'h0)] wire26;
  wire [(4'hc):(1'h0)] wire334;
  wire [(5'h11):(1'h0)] wire332;
  wire [(5'h10):(1'h0)] wire236;
  wire signed [(2'h2):(1'h0)] wire173;
  wire [(4'hc):(1'h0)] wire143;
  wire signed [(3'h5):(1'h0)] wire142;
  wire [(3'h5):(1'h0)] wire95;
  wire signed [(4'h9):(1'h0)] wire49;
  wire signed [(2'h3):(1'h0)] wire48;
  wire signed [(4'hb):(1'h0)] wire47;
  wire signed [(5'h16):(1'h0)] wire46;
  wire [(5'h11):(1'h0)] wire45;
  reg signed [(5'h15):(1'h0)] reg30 = (1'h0);
  reg [(5'h11):(1'h0)] reg31 = (1'h0);
  reg [(3'h4):(1'h0)] reg32 = (1'h0);
  reg [(5'h17):(1'h0)] reg37 = (1'h0);
  reg [(4'h9):(1'h0)] reg40 = (1'h0);
  reg [(4'hb):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg43 = (1'h0);
  reg [(3'h5):(1'h0)] reg44 = (1'h0);
  reg [(4'hb):(1'h0)] reg51 = (1'h0);
  reg [(3'h4):(1'h0)] reg52 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg53 = (1'h0);
  reg [(5'h12):(1'h0)] reg54 = (1'h0);
  reg [(5'h13):(1'h0)] reg55 = (1'h0);
  reg [(4'hb):(1'h0)] reg56 = (1'h0);
  reg [(5'h15):(1'h0)] reg60 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg61 = (1'h0);
  reg [(4'ha):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg68 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg70 = (1'h0);
  reg [(3'h7):(1'h0)] reg73 = (1'h0);
  reg [(4'he):(1'h0)] reg74 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg75 = (1'h0);
  reg [(5'h14):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg79 = (1'h0);
  reg [(2'h2):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg82 = (1'h0);
  reg [(5'h12):(1'h0)] reg84 = (1'h0);
  reg [(5'h11):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg94 = (1'h0);
  reg [(4'hb):(1'h0)] reg97 = (1'h0);
  reg [(2'h2):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg102 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg104 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg112 = (1'h0);
  reg [(2'h3):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg109 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg117 = (1'h0);
  reg [(5'h13):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg120 = (1'h0);
  reg [(5'h12):(1'h0)] reg121 = (1'h0);
  reg [(4'hd):(1'h0)] reg123 = (1'h0);
  reg [(4'hc):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg129 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg130 = (1'h0);
  reg [(5'h18):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg133 = (1'h0);
  reg [(5'h16):(1'h0)] reg136 = (1'h0);
  reg [(4'hf):(1'h0)] reg138 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg139 = (1'h0);
  reg [(5'h15):(1'h0)] reg147 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg158 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg163 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg167 = (1'h0);
  reg [(5'h18):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg172 = (1'h0);
  reg [(5'h14):(1'h0)] reg174 = (1'h0);
  reg [(3'h6):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg184 = (1'h0);
  reg [(2'h2):(1'h0)] reg185 = (1'h0);
  reg [(4'hd):(1'h0)] reg186 = (1'h0);
  reg [(5'h12):(1'h0)] reg187 = (1'h0);
  reg [(4'hf):(1'h0)] reg190 = (1'h0);
  reg [(3'h7):(1'h0)] reg191 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg192 = (1'h0);
  reg [(4'h9):(1'h0)] reg194 = (1'h0);
  reg [(2'h2):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg197 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg198 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg199 = (1'h0);
  reg [(3'h5):(1'h0)] reg200 = (1'h0);
  reg [(2'h2):(1'h0)] reg177 = (1'h0);
  reg [(4'hf):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg207 = (1'h0);
  reg [(4'h8):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg210 = (1'h0);
  reg [(5'h17):(1'h0)] reg212 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg213 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg215 = (1'h0);
  reg [(4'he):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg220 = (1'h0);
  reg [(4'hd):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg224 = (1'h0);
  reg [(4'he):(1'h0)] reg225 = (1'h0);
  reg [(2'h2):(1'h0)] reg233 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg235 = (1'h0);
  reg signed [(4'he):(1'h0)] reg234 = (1'h0);
  reg [(2'h3):(1'h0)] reg232 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar231 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg230 = (1'h0);
  reg [(5'h17):(1'h0)] reg229 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar228 = (1'h0);
  reg [(3'h7):(1'h0)] reg227 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg208 = (1'h0);
  reg [(5'h17):(1'h0)] forvar206 = (1'h0);
  reg [(4'h9):(1'h0)] reg218 = (1'h0);
  reg [(4'hf):(1'h0)] reg217 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg214 = (1'h0);
  reg [(3'h7):(1'h0)] reg211 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar208 = (1'h0);
  reg [(5'h15):(1'h0)] reg206 = (1'h0);
  reg [(5'h11):(1'h0)] reg205 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar204 = (1'h0);
  reg [(3'h7):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg201 = (1'h0);
  reg [(5'h13):(1'h0)] reg189 = (1'h0);
  reg [(3'h6):(1'h0)] forvar178 = (1'h0);
  reg [(3'h4):(1'h0)] reg196 = (1'h0);
  reg [(5'h14):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar189 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg188 = (1'h0);
  reg [(5'h15):(1'h0)] forvar183 = (1'h0);
  reg [(5'h10):(1'h0)] reg182 = (1'h0);
  reg [(3'h4):(1'h0)] reg180 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg178 = (1'h0);
  reg [(2'h2):(1'h0)] forvar177 = (1'h0);
  reg [(4'hb):(1'h0)] reg176 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar169 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg168 = (1'h0);
  reg [(5'h18):(1'h0)] forvar165 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg162 = (1'h0);
  reg [(5'h18):(1'h0)] reg161 = (1'h0);
  reg [(5'h12):(1'h0)] reg159 = (1'h0);
  reg [(3'h7):(1'h0)] reg157 = (1'h0);
  reg [(5'h13):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar155 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg154 = (1'h0);
  reg [(5'h18):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg151 = (1'h0);
  reg [(3'h7):(1'h0)] reg150 = (1'h0);
  reg [(4'hb):(1'h0)] reg149 = (1'h0);
  reg [(5'h13):(1'h0)] forvar148 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg146 = (1'h0);
  reg [(4'h8):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg144 = (1'h0);
  reg [(5'h18):(1'h0)] reg141 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg140 = (1'h0);
  reg [(4'h9):(1'h0)] reg137 = (1'h0);
  reg [(2'h2):(1'h0)] reg135 = (1'h0);
  reg [(2'h2):(1'h0)] forvar134 = (1'h0);
  reg [(5'h14):(1'h0)] reg132 = (1'h0);
  reg [(3'h5):(1'h0)] forvar128 = (1'h0);
  reg [(4'h9):(1'h0)] reg127 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg126 = (1'h0);
  reg [(3'h5):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg122 = (1'h0);
  reg [(5'h15):(1'h0)] reg118 = (1'h0);
  reg [(4'hb):(1'h0)] reg116 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg107 = (1'h0);
  reg [(4'hb):(1'h0)] forvar96 = (1'h0);
  reg [(3'h7):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg111 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar109 = (1'h0);
  reg [(5'h11):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar107 = (1'h0);
  reg [(5'h16):(1'h0)] reg103 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg100 = (1'h0);
  reg [(5'h10):(1'h0)] reg99 = (1'h0);
  reg [(4'hd):(1'h0)] reg98 = (1'h0);
  reg [(5'h15):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg93 = (1'h0);
  reg [(5'h13):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar89 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg88 = (1'h0);
  reg [(4'ha):(1'h0)] reg87 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg83 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg80 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg78 = (1'h0);
  reg [(4'hf):(1'h0)] reg77 = (1'h0);
  reg [(4'h9):(1'h0)] reg72 = (1'h0);
  reg [(3'h4):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar69 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg69 = (1'h0);
  reg [(5'h14):(1'h0)] reg67 = (1'h0);
  reg [(2'h2):(1'h0)] reg66 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg65 = (1'h0);
  reg signed [(4'he):(1'h0)] reg63 = (1'h0);
  reg [(2'h2):(1'h0)] reg62 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar59 = (1'h0);
  reg [(5'h14):(1'h0)] reg58 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg57 = (1'h0);
  reg [(4'hb):(1'h0)] forvar50 = (1'h0);
  reg [(5'h10):(1'h0)] forvar38 = (1'h0);
  reg [(4'hb):(1'h0)] reg42 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg39 = (1'h0);
  reg [(4'h9):(1'h0)] reg38 = (1'h0);
  reg [(5'h10):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg35 = (1'h0);
  reg [(5'h13):(1'h0)] reg34 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg33 = (1'h0);
  assign y = {wire334,
                 wire332,
                 wire236,
                 wire173,
                 wire143,
                 wire142,
                 wire95,
                 wire49,
                 wire48,
                 wire47,
                 wire46,
                 wire45,
                 reg30,
                 reg31,
                 reg32,
                 reg37,
                 reg40,
                 reg41,
                 reg43,
                 reg44,
                 reg51,
                 reg52,
                 reg53,
                 reg54,
                 reg55,
                 reg56,
                 reg60,
                 reg61,
                 reg64,
                 reg68,
                 reg70,
                 reg73,
                 reg74,
                 reg75,
                 reg76,
                 reg79,
                 reg81,
                 reg82,
                 reg84,
                 reg86,
                 reg90,
                 reg92,
                 reg94,
                 reg97,
                 reg101,
                 reg102,
                 reg104,
                 reg105,
                 reg106,
                 reg112,
                 reg113,
                 reg109,
                 reg117,
                 reg119,
                 reg120,
                 reg121,
                 reg123,
                 reg125,
                 reg129,
                 reg130,
                 reg131,
                 reg133,
                 reg136,
                 reg138,
                 reg139,
                 reg147,
                 reg152,
                 reg158,
                 reg160,
                 reg163,
                 reg166,
                 reg167,
                 reg171,
                 reg172,
                 reg174,
                 reg175,
                 reg179,
                 reg181,
                 reg184,
                 reg185,
                 reg186,
                 reg187,
                 reg190,
                 reg191,
                 reg192,
                 reg194,
                 reg195,
                 reg197,
                 reg198,
                 reg199,
                 reg200,
                 reg177,
                 reg183,
                 reg203,
                 reg207,
                 reg209,
                 reg210,
                 reg212,
                 reg213,
                 reg215,
                 reg219,
                 reg220,
                 reg222,
                 reg223,
                 reg224,
                 reg225,
                 reg233,
                 reg235,
                 reg234,
                 reg232,
                 forvar231,
                 reg230,
                 reg229,
                 forvar228,
                 reg227,
                 reg226,
                 reg221,
                 reg208,
                 forvar206,
                 reg218,
                 reg217,
                 reg216,
                 reg214,
                 reg211,
                 forvar208,
                 reg206,
                 reg205,
                 forvar204,
                 reg202,
                 reg201,
                 reg189,
                 forvar178,
                 reg196,
                 reg193,
                 forvar189,
                 reg188,
                 forvar183,
                 reg182,
                 reg180,
                 reg178,
                 forvar177,
                 reg176,
                 reg170,
                 forvar169,
                 reg168,
                 forvar165,
                 reg164,
                 reg162,
                 reg161,
                 reg159,
                 reg157,
                 reg156,
                 forvar155,
                 reg154,
                 reg153,
                 reg148,
                 reg151,
                 reg150,
                 reg149,
                 forvar148,
                 reg146,
                 reg145,
                 reg144,
                 reg141,
                 reg140,
                 reg137,
                 reg135,
                 forvar134,
                 reg132,
                 forvar128,
                 reg127,
                 reg126,
                 reg124,
                 reg122,
                 reg118,
                 reg116,
                 reg115,
                 reg107,
                 forvar96,
                 reg114,
                 reg111,
                 reg110,
                 forvar109,
                 reg108,
                 forvar107,
                 reg103,
                 reg100,
                 reg99,
                 reg98,
                 reg96,
                 reg93,
                 reg91,
                 forvar89,
                 reg88,
                 reg87,
                 reg85,
                 reg83,
                 reg80,
                 reg78,
                 reg77,
                 reg72,
                 reg71,
                 forvar69,
                 reg69,
                 reg67,
                 reg66,
                 reg65,
                 reg63,
                 reg62,
                 forvar59,
                 reg58,
                 reg57,
                 forvar50,
                 forvar38,
                 reg42,
                 reg39,
                 reg38,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned($signed(wire27[(2'h2):(1'h1)])))
        begin
          if (wire27)
            begin
              reg30 <= wire29[(4'ha):(1'h0)];
              reg31 <= (8'hbd);
            end
          else
            begin
              reg30 <= ($unsigned(($signed((wire27 >> reg30)) ?
                      $signed((~&reg31)) : ((+reg30) < {(8'ha2), (8'hb0)}))) ?
                  $signed(wire26) : $unsigned((((reg31 ?
                          wire26 : wire27) || {(8'hb6), reg30}) ?
                      $unsigned((~^wire28)) : wire27)));
              reg31 <= {reg31};
              reg32 <= ((8'haf) != $unsigned($signed(wire28[(1'h1):(1'h0)])));
              reg33 = $unsigned(reg32[(1'h1):(1'h0)]);
            end
          if (reg33[(4'hb):(3'h6)])
            begin
              reg34 = (7'h40);
              reg35 = (!{(reg31 ?
                      ($unsigned(reg31) ?
                          (wire29 ^ wire28) : reg32[(2'h3):(1'h1)]) : $unsigned((reg30 ?
                          reg31 : reg33))),
                  (&reg31[(3'h7):(3'h7)])});
              reg36 = (~{wire29[(4'h8):(2'h3)]});
            end
          else
            begin
              reg37 <= (^(+{((reg34 ? reg31 : wire29) ?
                      reg36 : (reg30 ? reg34 : wire27)),
                  $unsigned((!reg32))}));
              reg38 = ((((+(reg37 - reg34)) * reg37) || (|reg35)) ?
                  $unsigned({((~^reg36) && reg32[(1'h0):(1'h0)])}) : ((!$unsigned($unsigned(reg32))) ?
                      $signed($unsigned({reg37, reg34})) : reg37));
              reg39 = wire26;
              reg40 <= $unsigned(reg34);
              reg41 <= ({reg33[(3'h6):(1'h1)]} | $unsigned({reg30[(2'h3):(2'h3)],
                  wire29[(2'h3):(1'h1)]}));
            end
          reg42 = $signed(((reg36[(5'h10):(4'hf)] + $signed((reg36 ?
                  (8'hb2) : reg37))) ?
              reg38[(2'h3):(2'h3)] : ((&$signed(reg30)) ?
                  (8'hb0) : reg33[(5'h12):(5'h10)])));
        end
      else
        begin
          reg33 = ($unsigned(reg39) || $unsigned((^$signed(wire26))));
          reg37 <= {(^~(reg33 ?
                  $signed(reg39[(1'h0):(1'h0)]) : ((+(7'h4a)) ?
                      reg37 : (reg34 ^~ wire27))))};
          for (forvar38 = (1'h0); (forvar38 < (2'h3)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 = wire27;
            end
          reg40 <= $unsigned($signed(reg37[(5'h17):(5'h13)]));
        end
      reg43 <= (&$unsigned((^((+(8'had)) ~^ $unsigned(reg35)))));
      reg44 <= $unsigned(reg34[(5'h11):(4'hb)]);
    end
  assign wire45 = (~&{$signed(wire29[(3'h7):(3'h4)]),
                      ($unsigned($unsigned(wire26)) ?
                          ((wire28 * wire28) ? reg30 : (^~wire28)) : ((reg30 ?
                              reg37 : (8'h9e)) - (reg30 >= (8'hb6))))});
  assign wire46 = (reg40 ?
                      ($unsigned({$unsigned(wire27)}) >>> ($unsigned((!wire29)) ?
                          ((^~(7'h44)) <<< (wire45 ^ wire27)) : ($signed(reg44) <<< (wire26 & reg30)))) : ((-((~^wire26) != reg32)) < reg41));
  assign wire47 = (wire29 ?
                      {(~|wire45)} : $signed((($signed(wire26) << (8'hba)) | (8'hab))));
  assign wire48 = {$unsigned((($signed(wire46) == (reg31 & (8'h9d))) ?
                          wire46[(4'hc):(4'h8)] : $signed((wire29 == (8'ha4))))),
                      wire28[(3'h7):(2'h3)]};
  assign wire49 = $signed(reg32);
  always
    @(posedge clk) begin
      for (forvar50 = (1'h0); (forvar50 < (3'h4)); forvar50 = (forvar50 + (1'h1)))
        begin
          if (wire48[(1'h0):(1'h0)])
            begin
              reg51 <= $unsigned(($signed($unsigned(wire26[(4'he):(3'h7)])) ?
                  (($unsigned(wire26) << $signed(wire26)) ?
                      wire26 : wire49[(4'h8):(3'h4)]) : reg40[(4'h9):(3'h5)]));
              reg52 <= {$signed($unsigned(((wire28 ? wire47 : wire48) ?
                      reg40[(3'h6):(2'h2)] : (reg31 >>> forvar50))))};
            end
          else
            begin
              reg51 <= wire45[(3'h6):(1'h1)];
              reg52 <= $unsigned(((~^({(8'ha4)} ?
                      (forvar50 ^~ wire48) : (reg43 & wire47))) ?
                  ($unsigned($unsigned(reg31)) >= wire45[(4'h8):(3'h6)]) : (8'had)));
              reg53 <= wire48[(2'h2):(2'h2)];
            end
          reg54 <= forvar50[(2'h3):(1'h0)];
          reg55 <= $signed(({$unsigned(reg40)} || (^~($unsigned(wire46) >> (^wire29)))));
          reg56 <= (wire47[(2'h2):(1'h0)] || (8'haa));
        end
      reg57 = ({((!$signed(reg44)) ?
                  $signed(reg32[(2'h2):(2'h2)]) : ((reg44 ? reg52 : (8'hb6)) ?
                      {wire29, wire27} : (reg40 && reg51)))} ?
          ({(wire26 - wire28[(4'h8):(3'h5)])} ^~ $signed((-wire27))) : reg43[(3'h7):(3'h7)]);
      reg58 = {((8'hb8) | reg54[(4'hc):(3'h4)])};
      for (forvar59 = (1'h0); (forvar59 < (1'h1)); forvar59 = (forvar59 + (1'h1)))
        begin
          reg60 <= (($signed({reg55[(4'hb):(3'h7)]}) <= {(!((8'ha1) | reg52))}) >>> reg30);
          if (wire47)
            begin
              reg61 <= (reg44[(2'h3):(2'h3)] ?
                  $unsigned(($signed((wire26 ?
                      reg32 : reg40)) >> ((forvar59 < reg43) <= (reg60 ?
                      forvar50 : wire29)))) : reg37[(4'he):(4'hc)]);
              reg62 = {$unsigned((~^(|reg32[(1'h0):(1'h0)]))),
                  wire45[(4'hd):(4'h8)]};
            end
          else
            begin
              reg62 = {$unsigned((~^$unsigned(reg58[(4'hd):(4'h9)])))};
              reg63 = reg55[(5'h12):(3'h4)];
              reg64 <= {(({reg31} != ({wire45, reg40} ?
                      $signed(wire28) : ((8'hb7) ?
                          (7'h43) : (8'ha3)))) <<< (&$unsigned($unsigned(reg51))))};
              reg65 = (^reg37[(2'h2):(2'h2)]);
            end
        end
      reg66 = $unsigned($unsigned((reg31[(1'h0):(1'h0)] >> (^~(reg55 ?
          reg43 : reg64)))));
    end
  always
    @(posedge clk) begin
      reg67 = (reg32 ?
          reg51[(3'h6):(1'h0)] : $signed($unsigned($unsigned((reg54 & (8'ha0))))));
    end
  always
    @(posedge clk) begin
      reg68 <= reg64[(2'h2):(2'h2)];
    end
  always
    @(posedge clk) begin
      if ((^~($unsigned($signed((wire47 ?
          reg52 : reg40))) | (wire46[(5'h12):(5'h11)] ? wire47 : reg64))))
        begin
          reg69 = $signed((!$signed(wire29)));
        end
      else
        begin
          for (forvar69 = (1'h0); (forvar69 < (2'h2)); forvar69 = (forvar69 + (1'h1)))
            begin
              reg70 <= reg40;
              reg71 = $unsigned((^reg56));
              reg72 = ((((reg51[(3'h4):(3'h4)] ? reg55 : {reg70}) ^~ ((wire26 ?
                      wire47 : reg44) | {reg56})) ^~ $signed({$unsigned(reg71),
                      (reg41 ? forvar69 : reg52)})) ?
                  ((8'hb4) ?
                      (&{$unsigned(reg43)}) : $signed(wire28)) : (&reg70));
              reg73 <= $signed($signed(reg70[(2'h2):(2'h2)]));
            end
          if ($unsigned($unsigned((~reg73))))
            begin
              reg74 <= (~^((~|(8'hb4)) ?
                  ($unsigned(reg30) ?
                      {reg68,
                          wire27[(2'h2):(1'h0)]} : reg51) : ($unsigned(reg41) >= (-(reg53 ?
                      reg60 : reg52)))));
              reg75 <= $signed((|$signed($signed((reg72 ? reg30 : reg74)))));
              reg76 <= (~|$signed(($unsigned((reg75 ?
                  reg56 : (7'h42))) < ((reg51 ?
                  reg74 : wire48) != reg43[(5'h10):(4'hd)]))));
              reg77 = reg53[(3'h4):(3'h4)];
              reg78 = ($signed($signed(reg73[(3'h6):(1'h1)])) ?
                  (^~(|(8'hbb))) : ((+reg41[(4'h9):(2'h2)]) ?
                      $signed($unsigned({reg64})) : reg53[(2'h2):(1'h0)]));
            end
          else
            begin
              reg77 = $unsigned(reg68[(4'hc):(3'h6)]);
            end
          reg79 <= $signed(($signed($signed((reg69 >>> wire26))) <<< wire47));
          reg80 = $unsigned((reg73[(3'h6):(3'h5)] > reg78));
        end
    end
  always
    @(posedge clk) begin
      reg81 <= {reg44};
      if (reg56[(2'h2):(1'h0)])
        begin
          if ($signed({(-$unsigned($signed(wire29)))}))
            begin
              reg82 <= ({(8'hb2), (7'h47)} ?
                  (~{(reg51 ? {reg51} : {reg70, reg60}),
                      reg51[(4'h8):(1'h1)]}) : reg37);
              reg83 = ({$signed((^~((8'h9d) ? (8'h9c) : reg55))),
                  reg44[(3'h5):(2'h2)]} | reg64);
              reg84 <= {$signed(($unsigned($unsigned(reg68)) || {$unsigned((8'hbf))})),
                  {$unsigned(reg44)}};
              reg85 = $signed((+(({reg60} ?
                      $signed(reg37) : wire48[(2'h3):(2'h2)]) ?
                  ({reg41, reg41} ?
                      $unsigned(reg55) : (|reg31)) : reg79[(5'h17):(1'h1)])));
              reg86 <= (~reg53[(1'h1):(1'h1)]);
            end
          else
            begin
              reg82 <= (7'h4a);
              reg84 <= $signed((&$signed(wire45)));
              reg85 = ($unsigned($unsigned(({reg83} * (reg74 ?
                  wire46 : reg85)))) ^~ reg68[(3'h7):(1'h0)]);
            end
        end
      else
        begin
          reg83 = $unsigned(reg74);
        end
      if ($unsigned(reg64))
        begin
          reg87 = wire47[(3'h5):(1'h1)];
        end
      else
        begin
          reg87 = {($signed($signed((wire27 ?
                  reg74 : reg68))) >>> ((-reg86[(1'h1):(1'h0)]) ?
                  ($signed(reg32) ? $signed(reg83) : $signed(reg82)) : reg37)),
              $signed({wire48[(2'h2):(1'h1)], $unsigned((~(8'hb3)))})};
        end
      reg88 = reg70;
      for (forvar89 = (1'h0); (forvar89 < (1'h0)); forvar89 = (forvar89 + (1'h1)))
        begin
          if ((&wire46[(5'h13):(4'he)]))
            begin
              reg90 <= {($unsigned((~|$signed((8'ha4)))) + wire47[(2'h2):(1'h1)])};
              reg91 = (^{reg51[(4'ha):(4'h8)]});
            end
          else
            begin
              reg90 <= (~^reg82);
              reg91 = (~($unsigned(reg55) ?
                  (|{((8'hb8) ? reg64 : (8'ha4))}) : {reg32,
                      ({reg53, reg68} >> (~|reg68))}));
              reg92 <= wire49[(2'h3):(1'h1)];
              reg93 = (reg54 <<< (|reg91[(2'h3):(1'h0)]));
              reg94 <= (-(reg56 ?
                  ({(reg92 ? reg81 : reg73), $unsigned((8'hb3))} ?
                      $signed(reg60[(2'h2):(1'h0)]) : ($signed((8'ha5)) | (reg83 && (7'h46)))) : reg93[(3'h6):(1'h1)]));
            end
        end
    end
  assign wire95 = reg52;
  always
    @(posedge clk) begin
      if (((!reg76) < reg52[(3'h4):(2'h2)]))
        begin
          reg96 = $unsigned($unsigned(reg60[(2'h2):(1'h1)]));
          if (reg30)
            begin
              reg97 <= ({wire29,
                      ({reg92[(2'h3):(2'h3)], {reg92}} ?
                          reg40 : reg41[(4'h9):(2'h2)])} ?
                  $signed(reg43[(4'he):(4'he)]) : $signed((~$unsigned(reg73))));
            end
          else
            begin
              reg98 = ((^{(8'ha2)}) >> ($signed($unsigned($unsigned(reg68))) ?
                  (7'h49) : ($signed((~|(8'ha6))) <= $unsigned(reg68[(5'h11):(4'hf)]))));
              reg99 = ((^~{({reg73} ^~ reg82)}) << (&(((reg98 << reg31) ^ $unsigned(reg43)) ?
                  $unsigned({reg32}) : wire49)));
              reg100 = {(($signed((-wire47)) > reg53[(4'h8):(2'h3)]) ~^ $unsigned($signed(((7'h47) >> wire26)))),
                  (|reg37[(5'h14):(4'hd)])};
            end
          if ((~&{reg32, reg52}))
            begin
              reg101 <= $signed(((~^$unsigned($unsigned(wire27))) ?
                  (~^(+reg82)) : (reg98 ~^ ({reg73,
                      reg68} >= wire45[(2'h3):(2'h2)]))));
              reg102 <= {(($unsigned((reg54 ?
                      reg100 : reg97)) - reg53[(1'h0):(1'h0)]) < {($signed(reg86) ?
                          (reg76 ? wire45 : reg41) : (reg30 ? reg82 : wire27)),
                      $unsigned($unsigned(reg40))}),
                  $signed(((~&(&reg56)) * (7'h45)))};
            end
          else
            begin
              reg101 <= (|(~^$unsigned((|wire26))));
              reg103 = (wire95[(1'h1):(1'h0)] ?
                  $signed((({reg32} ? (|wire48) : $signed(reg74)) ?
                      (|(reg101 <= reg32)) : (^$unsigned(reg94)))) : ({$signed((&reg76)),
                          $signed($unsigned(wire26))} ?
                      reg100 : ({reg81, (7'h48)} * ((wire47 ?
                          reg75 : reg61) - {reg56, wire26}))));
              reg104 <= {reg73[(1'h0):(1'h0)],
                  (!({(wire26 ? reg64 : reg81)} >>> (7'h40)))};
              reg105 <= $unsigned($unsigned(reg53));
              reg106 <= {(reg51[(2'h3):(1'h1)] ^~ ($unsigned($signed(wire26)) ?
                      (wire46[(1'h0):(1'h0)] & (wire28 != wire49)) : {(&reg44)}))};
            end
          for (forvar107 = (1'h0); (forvar107 < (1'h0)); forvar107 = (forvar107 + (1'h1)))
            begin
              reg108 = {($signed(($signed(reg51) ?
                      wire27 : {reg43, wire26})) << (|reg81[(1'h0):(1'h0)]))};
            end
          for (forvar109 = (1'h0); (forvar109 < (1'h1)); forvar109 = (forvar109 + (1'h1)))
            begin
              reg110 = ((^$unsigned({wire29[(4'hd):(4'hd)],
                  $signed((8'hb8))})) ^ ($unsigned(((~(8'hba)) ~^ $signed(reg100))) ?
                  (reg79[(2'h2):(1'h0)] <= $unsigned((reg74 ?
                      wire49 : (7'h4a)))) : ((reg81[(1'h1):(1'h1)] ^~ (^wire49)) ?
                      reg82[(4'hc):(2'h2)] : reg37)));
              reg111 = ($signed($unsigned({reg53[(3'h6):(1'h1)]})) <<< $unsigned(((wire49[(4'h9):(3'h5)] >> reg102) ?
                  $signed((8'ha1)) : $unsigned({reg30}))));
              reg112 <= wire95[(1'h0):(1'h0)];
              reg113 <= $signed((|{{(reg99 ? (8'ha2) : (8'h9d))},
                  ((reg103 ? reg111 : (8'ha9)) ?
                      reg97[(3'h6):(3'h5)] : $signed((7'h40)))}));
              reg114 = $signed(((~&$signed($unsigned(wire49))) ?
                  reg81 : reg104));
            end
        end
      else
        begin
          for (forvar96 = (1'h0); (forvar96 < (2'h3)); forvar96 = (forvar96 + (1'h1)))
            begin
              reg97 <= ($signed($signed((8'ha6))) | reg43);
              reg101 <= (reg110[(4'hc):(2'h2)] ^ {(((reg44 >= (8'h9f)) < reg104) + $unsigned($signed(forvar96)))});
            end
          if (wire95[(2'h3):(1'h1)])
            begin
              reg102 <= reg111;
              reg103 = (reg113 ?
                  (~&{(|{(8'hac)}),
                      {(reg81 - reg75)}}) : $signed($unsigned($signed(wire48))));
              reg104 <= ((reg30[(5'h14):(2'h2)] ?
                      reg108 : ({$signed(reg103)} >= reg61)) ?
                  (((reg104 ?
                          reg111[(2'h2):(1'h0)] : $signed(reg104)) || reg73) ?
                      $unsigned(({reg56} >= reg54)) : wire27[(2'h2):(1'h0)]) : (|(-({reg92} ?
                      reg40 : $unsigned(reg92)))));
              reg105 <= ((&{$signed((+reg73))}) >> (~reg110[(3'h7):(2'h3)]));
            end
          else
            begin
              reg103 = $unsigned((~^$unsigned($unsigned($unsigned(reg64)))));
            end
          reg107 = wire45[(3'h5):(2'h3)];
          reg109 <= $signed({(reg96 ?
                  {(reg54 >>> (7'h47)),
                      $unsigned(wire49)} : (reg94 >> (!wire26))),
              (reg96[(5'h12):(2'h2)] ?
                  (reg108[(4'he):(1'h1)] ~^ (wire29 ?
                      forvar107 : reg103)) : reg60[(2'h3):(1'h0)])});
          reg112 <= reg30[(4'hb):(3'h5)];
        end
      reg115 = ($signed(reg82[(4'hc):(4'h8)]) | reg86);
      if (((-reg30) & $unsigned({$signed(reg54[(4'hc):(4'hb)]), (&reg104)})))
        begin
          reg116 = reg73[(1'h0):(1'h0)];
          if (wire28)
            begin
              reg117 <= (~&wire48[(2'h2):(1'h0)]);
              reg118 = ({$signed($signed($signed(reg79))),
                      $signed(($signed(reg74) ?
                          ((8'ha8) != reg54) : reg102[(4'hc):(4'h9)]))} ?
                  reg60[(2'h2):(1'h1)] : wire26);
              reg119 <= (reg104 + reg60[(1'h0):(1'h0)]);
              reg120 <= $unsigned(reg32[(1'h0):(1'h0)]);
            end
          else
            begin
              reg117 <= $unsigned($unsigned(reg116[(4'h9):(3'h7)]));
              reg119 <= ($unsigned(wire95[(1'h1):(1'h0)]) ^ (&wire45[(4'h9):(2'h2)]));
              reg120 <= {(^~{((wire95 ? reg53 : reg73) == reg110)}),
                  (!(($unsigned((8'hb5)) >= (reg113 ? reg96 : (8'ha6))) ?
                      (^~reg43) : reg61[(2'h2):(1'h0)]))};
              reg121 <= ((forvar109 ?
                  (reg100 ?
                      wire27[(4'h9):(3'h7)] : $unsigned($signed(reg70))) : reg44) - (reg51 <= $signed(((reg100 >> (8'ha4)) ?
                  (reg79 ? reg44 : (8'hbb)) : (reg37 > reg106)))));
              reg122 = ({($signed((7'h48)) ?
                          reg102[(4'hf):(4'hf)] : (reg110[(1'h1):(1'h0)] ?
                              ((7'h49) ? reg99 : reg74) : ((8'haa) ?
                                  reg44 : (8'ha7)))),
                      $unsigned(($unsigned((8'ha1)) != (!wire48)))} ?
                  reg97 : wire27[(2'h2):(2'h2)]);
            end
          if (reg120)
            begin
              reg123 <= (+$unsigned($unsigned(({reg74} >>> (~reg110)))));
              reg124 = reg53;
              reg125 <= (-$signed($signed($unsigned($signed(reg98)))));
              reg126 = (reg68[(5'h10):(3'h6)] ?
                  ((&reg104) <= ((((7'h46) ? reg97 : wire47) ?
                          $signed(reg103) : (~&reg117)) ?
                      $signed((reg92 ?
                          reg97 : reg86)) : $unsigned(((7'h43) >>> reg73)))) : ((-(+forvar107[(3'h7):(3'h6)])) ?
                      $unsigned(({reg70} ?
                          $unsigned(reg31) : $signed((7'h43)))) : $unsigned(({(7'h42),
                          reg104} || (reg32 ? (8'ha3) : reg60)))));
            end
          else
            begin
              reg124 = $unsigned({$signed(({wire95, reg122} ?
                      reg114[(3'h4):(1'h0)] : $signed(reg56))),
                  ({(reg86 ? reg64 : reg56), (reg98 ? reg90 : reg74)} ?
                      $signed(reg118) : $signed((|reg56)))});
              reg125 <= (+$signed(({wire28} & (~|(wire95 ? reg79 : reg105)))));
              reg126 = reg119;
              reg127 = reg82[(1'h1):(1'h1)];
            end
          for (forvar128 = (1'h0); (forvar128 < (2'h2)); forvar128 = (forvar128 + (1'h1)))
            begin
              reg129 <= reg113;
              reg130 <= (&($unsigned(((reg79 <= (8'had)) != (wire29 >> wire29))) == reg40[(3'h6):(2'h3)]));
              reg131 <= (&{((|(reg124 ? reg41 : (7'h42))) ?
                      (&(+reg115)) : reg55),
                  $signed(reg101)});
              reg132 = {((-(~|{reg41, reg101})) ?
                      reg92 : $signed((reg98 ? $unsigned(reg84) : (^reg112)))),
                  reg108[(4'hb):(1'h0)]};
            end
          reg133 <= reg40[(1'h1):(1'h0)];
        end
      else
        begin
          reg117 <= (!reg96[(3'h7):(3'h6)]);
        end
      if ($unsigned(($signed((reg96[(4'h8):(2'h2)] < $unsigned(reg31))) ?
          (^~{((8'ha7) ^~ reg123)}) : (-{reg81[(1'h0):(1'h0)], reg108}))))
        begin
          for (forvar134 = (1'h0); (forvar134 < (1'h1)); forvar134 = (forvar134 + (1'h1)))
            begin
              reg135 = $unsigned(reg105);
              reg136 <= $signed(reg99[(3'h6):(3'h4)]);
              reg137 = reg105;
              reg138 <= reg64;
            end
          reg139 <= {((^~reg117[(4'h8):(2'h2)]) ^ (!wire95[(1'h1):(1'h0)]))};
          reg140 = (($unsigned(reg138) > (^(^forvar109))) >>> $signed(reg133[(5'h14):(3'h5)]));
        end
      else
        begin
          for (forvar134 = (1'h0); (forvar134 < (2'h3)); forvar134 = (forvar134 + (1'h1)))
            begin
              reg136 <= $signed(forvar134);
              reg138 <= $signed(reg118[(5'h10):(4'hb)]);
            end
        end
      reg141 = ((($unsigned(((8'h9e) >> reg79)) << $unsigned({reg129})) || reg133[(5'h14):(4'hc)]) ?
          ((wire29 ? $unsigned((~|reg99)) : (reg132 * reg98)) ?
              ($unsigned($unsigned(reg115)) ?
                  $signed(((8'h9c) >= (8'h9c))) : {reg92[(4'hc):(3'h7)]}) : {(~|$signed(reg107))}) : {($unsigned(reg107) >> (forvar128 << reg104[(3'h5):(3'h4)])),
              reg138});
    end
  assign wire142 = {$signed($unsigned(reg40))};
  assign wire143 = reg53;
  always
    @(posedge clk) begin
      reg144 = reg55;
      reg145 = (wire48[(2'h3):(1'h1)] >> wire143);
      if (reg84)
        begin
          reg146 = reg92[(5'h14):(5'h13)];
          reg147 <= (($signed({reg44}) ?
                  (^$unsigned($signed((8'hbc)))) : reg79) ?
              (~$unsigned($unsigned($signed(reg86)))) : $unsigned($signed({$signed(reg146)})));
        end
      else
        begin
          reg147 <= reg92;
        end
      if ($unsigned($unsigned($unsigned({$signed(reg123),
          (reg121 ? wire47 : reg123)}))))
        begin
          for (forvar148 = (1'h0); (forvar148 < (1'h1)); forvar148 = (forvar148 + (1'h1)))
            begin
              reg149 = ((7'h45) ?
                  wire26[(2'h2):(1'h0)] : ((|$unsigned($signed(reg52))) << (8'hbb)));
              reg150 = ($signed(((^((7'h48) << reg138)) ^ $signed(((8'hba) ?
                      reg86 : reg136)))) ?
                  ((&($unsigned(reg60) ?
                      (!(7'h47)) : wire26)) > reg76[(4'hc):(4'ha)]) : ($signed(($signed(reg146) ?
                          ((8'hbc) ^ reg138) : (&reg144))) ?
                      $signed((|$signed(reg76))) : $signed({reg144, (8'ha7)})));
              reg151 = (+({reg32[(1'h1):(1'h1)]} ?
                  ($unsigned((|(8'hbc))) ?
                      $signed((reg81 <= (8'ha3))) : $unsigned(reg75[(2'h2):(1'h0)])) : $unsigned({(reg119 >>> reg120),
                      wire29})));
            end
          reg152 <= (reg139[(3'h4):(3'h4)] ?
              reg52 : ((~$signed(((8'ha4) ? reg131 : wire47))) ?
                  $unsigned(reg70) : $unsigned($unsigned({reg144}))));
        end
      else
        begin
          if ($unsigned(reg109[(3'h4):(2'h2)]))
            begin
              reg148 = (!$unsigned(wire47[(1'h1):(1'h0)]));
            end
          else
            begin
              reg152 <= ({$signed($signed((reg64 ~^ (8'ha7))))} >>> $signed($signed($unsigned({reg92}))));
              reg153 = ((~|{$unsigned($unsigned(wire49))}) ?
                  $unsigned((~&reg64)) : {($signed((8'hb1)) ?
                          ($signed(reg64) == (reg121 ?
                              reg104 : reg106)) : $unsigned((reg133 >> wire49)))});
              reg154 = $unsigned($signed((reg52[(1'h0):(1'h0)] || reg151[(3'h7):(3'h4)])));
            end
          for (forvar155 = (1'h0); (forvar155 < (1'h0)); forvar155 = (forvar155 + (1'h1)))
            begin
              reg156 = reg152;
              reg157 = reg154[(2'h3):(1'h0)];
              reg158 <= reg94[(1'h0):(1'h0)];
              reg159 = reg121[(4'ha):(3'h7)];
            end
          if ($signed((-$signed(reg55[(4'ha):(2'h2)]))))
            begin
              reg160 <= reg30;
              reg161 = $unsigned(reg97);
              reg162 = $unsigned($signed(reg60[(2'h3):(1'h1)]));
            end
          else
            begin
              reg161 = (-forvar148);
              reg163 <= $signed(((reg129[(5'h12):(3'h5)] <= ({(7'h46)} ?
                      reg153 : $signed(reg30))) ?
                  reg144[(2'h3):(2'h2)] : ($signed($unsigned(reg160)) ?
                      $unsigned((8'hab)) : $signed(reg94))));
            end
        end
      reg164 = (reg73[(3'h5):(1'h0)] ^~ ({(^(^(8'hbe)))} - reg82[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      for (forvar165 = (1'h0); (forvar165 < (2'h3)); forvar165 = (forvar165 + (1'h1)))
        begin
          if (reg56[(3'h7):(3'h7)])
            begin
              reg166 <= $unsigned((reg105 ?
                  $unsigned(($signed(reg82) ?
                      reg30 : {reg64})) : reg160[(1'h1):(1'h1)]));
              reg167 <= ({reg97} >= (reg166[(3'h6):(3'h5)] < reg166));
            end
          else
            begin
              reg166 <= $signed({($unsigned((reg56 ? reg105 : reg60)) == {reg76,
                      reg109[(3'h4):(2'h2)]}),
                  reg60[(1'h0):(1'h0)]});
              reg168 = ($signed(reg112[(4'ha):(3'h7)]) & reg40[(4'h8):(4'h8)]);
            end
        end
      for (forvar169 = (1'h0); (forvar169 < (1'h1)); forvar169 = (forvar169 + (1'h1)))
        begin
          reg170 = $unsigned((reg81[(1'h1):(1'h1)] ?
              $signed(reg105[(4'h9):(3'h4)]) : $unsigned($unsigned($signed(reg123)))));
        end
      reg171 <= (($unsigned(reg147[(2'h2):(1'h1)]) >>> $unsigned($signed((reg82 - reg51)))) ?
          reg123[(2'h3):(2'h2)] : reg44);
      reg172 <= {((~(reg90[(2'h2):(1'h0)] ?
              $signed(reg94) : (8'hb9))) >> $signed(((reg131 || (8'hab)) ?
              {reg84} : $signed(reg86)))),
          {$signed(($signed(reg136) <<< $unsigned(reg102)))}};
    end
  assign wire173 = wire29;
  always
    @(posedge clk) begin
      reg174 <= $signed((~|($signed(wire143) <= reg73[(1'h1):(1'h1)])));
    end
  always
    @(posedge clk) begin
      reg175 <= ({$unsigned((8'ha5))} ~^ $signed($unsigned(reg101)));
      reg176 = reg112[(2'h3):(1'h0)];
      if ($unsigned((+$signed(reg139[(1'h1):(1'h1)]))))
        begin
          for (forvar177 = (1'h0); (forvar177 < (2'h2)); forvar177 = (forvar177 + (1'h1)))
            begin
              reg178 = reg32;
              reg179 <= $unsigned({$signed($unsigned(reg90)),
                  reg75[(2'h2):(1'h0)]});
              reg180 = {(reg125[(3'h7):(3'h5)] ?
                      $signed($signed($signed(reg152))) : {((+wire49) ?
                              $unsigned(reg70) : $signed(reg172))})};
              reg181 <= reg178;
            end
          reg182 = reg53;
          for (forvar183 = (1'h0); (forvar183 < (1'h1)); forvar183 = (forvar183 + (1'h1)))
            begin
              reg184 <= $signed((~^{((~|reg73) < (wire95 ^ reg160))}));
              reg185 <= (~|$signed((wire28[(3'h6):(3'h5)] ?
                  reg101 : reg139[(3'h5):(1'h1)])));
              reg186 <= $unsigned($unsigned((((~wire142) >> $signed(reg40)) > ({reg120} <= reg129[(3'h5):(1'h0)]))));
              reg187 <= reg106;
              reg188 = ((7'h44) ? reg178 : $unsigned(reg53[(2'h3):(1'h0)]));
            end
          for (forvar189 = (1'h0); (forvar189 < (3'h4)); forvar189 = (forvar189 + (1'h1)))
            begin
              reg190 <= $signed($signed({(7'h48),
                  $signed((reg56 <<< (7'h47)))}));
              reg191 <= $unsigned(reg101);
              reg192 <= reg31[(2'h2):(1'h0)];
              reg193 = (|(^~(^reg60)));
            end
          if (reg187[(5'h12):(4'h9)])
            begin
              reg194 <= reg60;
              reg195 <= {reg101[(2'h2):(2'h2)]};
              reg196 = $signed({wire47});
              reg197 <= $signed({$signed(reg136[(5'h11):(5'h10)]),
                  $signed({$signed(reg158), reg79})});
            end
          else
            begin
              reg196 = {(reg61 ?
                      (($unsigned(forvar189) << $signed(reg92)) ?
                          reg121[(4'hc):(2'h2)] : $signed((+reg105))) : (~|wire26))};
              reg197 <= (reg158[(5'h10):(4'hf)] ?
                  reg92[(5'h13):(5'h12)] : reg131[(5'h11):(4'hf)]);
              reg198 <= $signed(reg188[(4'h9):(3'h7)]);
              reg199 <= wire95[(1'h1):(1'h1)];
              reg200 <= $signed((((!(^reg53)) ?
                      (wire142[(3'h5):(3'h4)] ~^ reg79[(2'h3):(1'h0)]) : reg192[(5'h12):(2'h2)]) ?
                  (((reg194 <= reg193) < $unsigned(reg56)) ^ {reg182[(3'h7):(2'h2)],
                      $signed((8'ha6))}) : $signed($unsigned(((8'had) <= wire27)))));
            end
        end
      else
        begin
          reg177 <= $unsigned($signed($unsigned((reg51[(4'h9):(1'h1)] ?
              (&reg82) : reg193[(3'h6):(3'h4)]))));
          for (forvar178 = (1'h0); (forvar178 < (1'h0)); forvar178 = (forvar178 + (1'h1)))
            begin
              reg180 = reg113[(2'h3):(1'h0)];
              reg182 = (^reg133[(3'h4):(3'h4)]);
              reg183 <= (8'hb6);
              reg188 = $signed({reg194, reg102[(3'h5):(2'h3)]});
              reg189 = reg60[(2'h2):(2'h2)];
            end
          reg193 = (wire47[(4'ha):(3'h4)] ?
              $unsigned(reg31[(4'ha):(1'h0)]) : (~({$signed(reg60)} * (~^$signed(reg197)))));
        end
      reg201 = $signed(wire45[(3'h7):(3'h4)]);
    end
  always
    @(posedge clk) begin
      reg202 = $signed(((reg130 <= ($unsigned((8'h9d)) << (reg200 ~^ reg125))) ?
          $unsigned(($signed(reg199) <= {reg171,
              reg44})) : ($unsigned($signed(reg147)) ^ {$signed(reg90),
              (reg79 ? (8'hbb) : reg76)})));
      reg203 <= $signed(((reg43[(3'h6):(3'h4)] || reg187) <<< reg56[(2'h2):(1'h0)]));
    end
  always
    @(posedge clk) begin
      for (forvar204 = (1'h0); (forvar204 < (1'h1)); forvar204 = (forvar204 + (1'h1)))
        begin
          reg205 = (|((reg123 > reg136[(5'h13):(3'h5)]) || reg123[(4'h8):(4'h8)]));
        end
      if ((((reg109[(3'h6):(3'h6)] ? reg119[(2'h2):(2'h2)] : {$signed(reg97)}) ?
              reg97 : $unsigned($unsigned($unsigned((8'ha2))))) ?
          ((wire48 - $unsigned((!(7'h43)))) ?
              (~(!reg190[(4'h8):(3'h7)])) : reg76) : reg139))
        begin
          reg206 = reg187;
          reg207 <= ((reg109 - ($unsigned(reg139[(3'h4):(1'h0)]) <<< $unsigned((~reg175)))) < $unsigned({reg163,
              $unsigned($unsigned((8'hbb)))}));
          for (forvar208 = (1'h0); (forvar208 < (1'h1)); forvar208 = (forvar208 + (1'h1)))
            begin
              reg209 <= ({(8'hae)} + (&((~&$signed((7'h48))) ~^ (^~$unsigned(reg191)))));
              reg210 <= (8'hbf);
              reg211 = reg186[(4'hb):(4'h8)];
            end
          if ((reg187[(2'h2):(1'h1)] ?
              ((|{reg166,
                  (reg185 <<< (8'h9c))}) < (+($signed(wire95) == (reg200 < reg177)))) : reg84))
            begin
              reg212 <= (($signed((~^$signed(reg86))) || (8'hb8)) ?
                  {reg94} : $unsigned(((8'ha4) ?
                      reg79[(5'h14):(4'h8)] : (-(^wire45)))));
              reg213 <= reg211;
              reg214 = reg119;
              reg215 <= $unsigned(reg174);
              reg216 = {reg113, reg43[(1'h0):(1'h0)]};
            end
          else
            begin
              reg212 <= reg90;
              reg214 = $unsigned(((wire26 - {$signed(wire142)}) ?
                  reg79 : ({$signed(reg192)} ?
                      ({reg133,
                          reg138} < $signed(reg205)) : (((8'haa) && reg174) ?
                          $signed(reg174) : (-reg213)))));
              reg216 = reg102;
              reg217 = reg190[(3'h4):(2'h3)];
            end
          reg218 = ($unsigned(((reg105 ?
              (reg123 >>> reg138) : $unsigned((8'ha4))) <= reg53[(3'h5):(2'h2)])) >> reg52);
        end
      else
        begin
          for (forvar206 = (1'h0); (forvar206 < (1'h0)); forvar206 = (forvar206 + (1'h1)))
            begin
              reg208 = reg131;
            end
          if ($signed((reg139[(1'h0):(1'h0)] | (forvar208[(3'h4):(1'h1)] ?
              $unsigned({reg210}) : $signed({reg113})))))
            begin
              reg209 <= $signed((&reg207));
              reg210 <= {reg185[(2'h2):(1'h1)], reg185[(1'h0):(1'h0)]};
              reg211 = ((~^$unsigned(((~&forvar208) >= wire26))) ?
                  (-reg51) : {$unsigned($unsigned((reg112 <= (8'ha8))))});
              reg212 <= (reg41[(2'h3):(2'h2)] ?
                  ($signed(reg82[(5'h10):(4'h9)]) <= (-{(reg123 ?
                          reg68 : reg109)})) : $signed($unsigned(($unsigned(reg172) ?
                      reg184[(4'ha):(1'h0)] : {reg113}))));
              reg213 <= reg64[(4'h8):(3'h5)];
            end
          else
            begin
              reg211 = ($signed({((reg73 ?
                      forvar204 : reg133) || $signed(reg192)),
                  reg121[(5'h10):(4'h9)]}) + {(reg119 ? reg84 : reg102)});
              reg214 = wire26;
            end
        end
      if (($signed({((reg152 ? reg183 : reg102) ?
                  $signed(reg208) : reg112[(4'h9):(3'h7)])}) ?
          reg119 : ((($unsigned(wire29) >>> {reg191, reg94}) ? reg55 : reg192) ?
              (reg104 - $signed((8'hbe))) : (+(((8'ha5) ~^ reg32) ^ $signed(reg31))))))
        begin
          if ((^~reg86))
            begin
              reg219 <= wire142;
              reg220 <= reg61[(5'h10):(5'h10)];
            end
          else
            begin
              reg221 = (|reg79);
              reg222 <= ((8'hb7) >>> reg214);
              reg223 <= ((&$unsigned((reg191 ?
                  (reg54 & reg139) : reg163[(1'h1):(1'h0)]))) << ((7'h45) ?
                  (reg174 >= {(-reg214)}) : reg172));
              reg224 <= $signed($unsigned({reg212, reg73[(1'h0):(1'h0)]}));
            end
          if ((8'hb4))
            begin
              reg225 <= (wire48[(2'h2):(2'h2)] << $signed(reg221));
              reg226 = reg86[(4'hb):(4'h9)];
            end
          else
            begin
              reg226 = $unsigned(reg105);
              reg227 = reg133;
            end
          for (forvar228 = (1'h0); (forvar228 < (1'h0)); forvar228 = (forvar228 + (1'h1)))
            begin
              reg229 = reg41[(4'h8):(2'h3)];
            end
        end
      else
        begin
          if ($unsigned(((~|$signed({wire173, reg220})) | {(+((8'ha6) ?
                  reg208 : (8'hbb)))})))
            begin
              reg219 <= reg147[(4'hc):(1'h0)];
            end
          else
            begin
              reg219 <= $signed((~^reg171[(2'h3):(1'h1)]));
              reg221 = reg223[(3'h7):(3'h4)];
              reg222 <= $signed((~|$signed((^~$signed(reg102)))));
              reg226 = $unsigned({reg121[(3'h4):(3'h4)],
                  (reg177[(2'h2):(1'h1)] << $signed((reg208 & reg222)))});
            end
        end
      reg230 = (^~reg70[(3'h5):(1'h1)]);
      for (forvar231 = (1'h0); (forvar231 < (2'h3)); forvar231 = (forvar231 + (1'h1)))
        begin
          reg232 = (reg229 + $unsigned(((~|reg121[(1'h0):(1'h0)]) ?
              wire142[(2'h3):(1'h1)] : ($signed(reg75) | reg211))));
        end
    end
  always
    @(posedge clk) begin
      reg233 <= (^~{reg181});
      reg234 = reg70;
      reg235 = (+$signed((~&reg220)));
    end
  assign wire236 = (((&reg97[(1'h0):(1'h0)]) > (~|{(wire95 == reg219)})) >= reg43[(4'hc):(3'h6)]);
  module237 #() modinst333 (.wire240(reg167), .wire241(reg60), .wire242(reg112), .wire238(reg186), .clk(clk), .wire239(reg86), .y(wire332));
  assign wire334 = {reg75[(2'h2):(1'h1)]};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module237
#(parameter param330 = ((|((~((8'hb2) ? (7'h44) : (8'hbc))) ? {(|(8'hab)), {(7'h48)}} : {(+(8'h9e)), ((7'h4a) ? (8'had) : (7'h42))})) ? (~|({(^~(8'h9d))} << (^~((7'h43) ? (8'hb0) : (8'hb3))))) : ((-(((8'hbe) || (8'hb7)) ? ((8'hb8) ^~ (8'hab)) : ((7'h49) ? (8'ha4) : (8'hbe)))) ? (({(8'haa)} ? ((8'hab) == (8'hb9)) : {(8'haf), (7'h45)}) && (~^((7'h45) ^ (7'h46)))) : ((^(~(8'ha0))) ? (7'h44) : (((8'ha2) ? (8'hb4) : (8'hb5)) ? ((7'h49) ? (8'hab) : (8'hb2)) : (~|(8'ha4)))))), 
parameter param331 = param330)
(y, clk, wire242, wire241, wire240, wire239, wire238);
  output wire [(32'h49a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire242;
  input wire [(5'h15):(1'h0)] wire241;
  input wire [(5'h17):(1'h0)] wire240;
  input wire signed [(3'h7):(1'h0)] wire239;
  input wire [(4'hd):(1'h0)] wire238;
  wire [(4'hc):(1'h0)] wire321;
  wire signed [(5'h13):(1'h0)] wire320;
  wire [(3'h4):(1'h0)] wire288;
  wire signed [(2'h2):(1'h0)] wire284;
  wire signed [(5'h18):(1'h0)] wire283;
  wire [(5'h17):(1'h0)] wire273;
  wire signed [(4'hf):(1'h0)] wire244;
  wire signed [(4'hb):(1'h0)] wire243;
  reg signed [(2'h2):(1'h0)] reg329 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg327 = (1'h0);
  reg [(5'h13):(1'h0)] reg326 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg325 = (1'h0);
  reg [(4'hb):(1'h0)] reg322 = (1'h0);
  reg [(2'h2):(1'h0)] reg319 = (1'h0);
  reg [(5'h18):(1'h0)] reg312 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg310 = (1'h0);
  reg [(5'h10):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg306 = (1'h0);
  reg [(3'h6):(1'h0)] reg305 = (1'h0);
  reg [(3'h4):(1'h0)] reg304 = (1'h0);
  reg [(5'h11):(1'h0)] reg303 = (1'h0);
  reg [(4'he):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg298 = (1'h0);
  reg [(5'h10):(1'h0)] reg297 = (1'h0);
  reg [(5'h12):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg292 = (1'h0);
  reg [(4'ha):(1'h0)] reg291 = (1'h0);
  reg [(4'hf):(1'h0)] reg286 = (1'h0);
  reg [(5'h18):(1'h0)] reg282 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg281 = (1'h0);
  reg [(5'h14):(1'h0)] reg280 = (1'h0);
  reg [(5'h12):(1'h0)] reg279 = (1'h0);
  reg [(4'he):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg271 = (1'h0);
  reg [(4'he):(1'h0)] reg267 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg265 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg263 = (1'h0);
  reg [(5'h16):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg261 = (1'h0);
  reg [(4'hb):(1'h0)] reg259 = (1'h0);
  reg [(5'h18):(1'h0)] reg258 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg256 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg255 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg249 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg248 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg246 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg328 = (1'h0);
  reg [(5'h15):(1'h0)] reg324 = (1'h0);
  reg [(3'h6):(1'h0)] forvar323 = (1'h0);
  reg [(4'h8):(1'h0)] reg318 = (1'h0);
  reg [(5'h13):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg316 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg315 = (1'h0);
  reg [(5'h11):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg313 = (1'h0);
  reg [(5'h12):(1'h0)] reg309 = (1'h0);
  reg [(5'h13):(1'h0)] forvar308 = (1'h0);
  reg [(5'h17):(1'h0)] reg301 = (1'h0);
  reg [(4'hb):(1'h0)] reg300 = (1'h0);
  reg [(4'hc):(1'h0)] reg299 = (1'h0);
  reg [(4'hc):(1'h0)] reg296 = (1'h0);
  reg [(3'h7):(1'h0)] reg295 = (1'h0);
  reg [(5'h13):(1'h0)] reg293 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg290 = (1'h0);
  reg [(3'h5):(1'h0)] forvar289 = (1'h0);
  reg [(4'h9):(1'h0)] reg287 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg285 = (1'h0);
  reg [(4'hf):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar276 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg275 = (1'h0);
  reg [(5'h14):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg270 = (1'h0);
  reg [(4'h9):(1'h0)] reg269 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar268 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar260 = (1'h0);
  reg [(4'ha):(1'h0)] reg257 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg254 = (1'h0);
  reg [(4'h9):(1'h0)] reg253 = (1'h0);
  reg [(5'h17):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg247 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar245 = (1'h0);
  assign y = {wire321,
                 wire320,
                 wire288,
                 wire284,
                 wire283,
                 wire273,
                 wire244,
                 wire243,
                 reg329,
                 reg327,
                 reg326,
                 reg325,
                 reg322,
                 reg319,
                 reg312,
                 reg311,
                 reg310,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg298,
                 reg297,
                 reg294,
                 reg292,
                 reg291,
                 reg286,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg274,
                 reg271,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg259,
                 reg258,
                 reg256,
                 reg255,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg246,
                 reg328,
                 reg324,
                 forvar323,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg309,
                 forvar308,
                 reg301,
                 reg300,
                 reg299,
                 reg296,
                 reg295,
                 reg293,
                 reg290,
                 forvar289,
                 reg287,
                 reg285,
                 reg278,
                 reg277,
                 forvar276,
                 reg275,
                 reg272,
                 reg270,
                 reg269,
                 forvar268,
                 reg260,
                 forvar260,
                 reg257,
                 reg254,
                 reg253,
                 reg252,
                 reg247,
                 forvar245,
                 (1'h0)};
  assign wire243 = ($signed($unsigned((wire239 ?
                           (wire240 + wire241) : (wire240 >= wire239)))) ?
                       ((!{(|wire242), (wire240 ? (8'hb0) : wire242)}) ?
                           wire240 : wire239) : wire242);
  assign wire244 = $signed((~|wire239));
  always
    @(posedge clk) begin
      for (forvar245 = (1'h0); (forvar245 < (1'h1)); forvar245 = (forvar245 + (1'h1)))
        begin
          reg246 <= {$signed(wire244),
              ({($signed(wire240) ? wire239 : (wire241 ? wire239 : wire240)),
                  wire241[(5'h15):(3'h5)]} ^~ (wire238 ?
                  wire242[(4'hf):(4'he)] : (wire242 ?
                      wire243[(3'h7):(3'h6)] : (wire240 << (8'hbb)))))};
          if (wire242[(4'he):(4'hc)])
            begin
              reg247 = ($unsigned(wire238[(4'h8):(3'h4)]) && $unsigned(wire242[(3'h5):(2'h2)]));
            end
          else
            begin
              reg248 <= forvar245;
              reg249 <= $unsigned(((wire239[(1'h0):(1'h0)] * ((wire238 ^ (8'hb5)) ?
                      $unsigned(reg246) : $signed(wire238))) ?
                  (7'h45) : ({(wire239 & wire241)} > wire243)));
            end
        end
      reg250 <= ((^~(^$signed({(8'hb0)}))) + $signed((wire239 == (-reg246[(1'h1):(1'h0)]))));
      if (wire238[(1'h0):(1'h0)])
        begin
          if (wire242)
            begin
              reg251 <= $signed(reg247);
              reg252 = ($unsigned(((~&wire240) <= wire244)) ?
                  (((wire238 ? reg249 : (wire240 * (8'ha4))) ^~ (8'hb6)) ?
                      (forvar245[(1'h1):(1'h0)] < ({wire243,
                          (7'h45)} >>> wire239)) : wire242) : {($unsigned(reg246[(2'h2):(2'h2)]) ?
                          $signed(((8'hb8) ^~ reg249)) : (wire242 ?
                              $unsigned(wire243) : reg250[(3'h7):(3'h6)]))});
              reg253 = $unsigned($unsigned(reg249[(5'h10):(3'h6)]));
            end
          else
            begin
              reg252 = wire244;
            end
          reg254 = reg249;
          if ($signed(wire239))
            begin
              reg255 <= (^wire239[(3'h4):(1'h1)]);
              reg256 <= $signed(wire242[(4'hc):(2'h3)]);
              reg257 = ($unsigned($signed(reg256[(1'h1):(1'h0)])) ?
                  (^~$unsigned($signed($unsigned(wire238)))) : (|(~&((^~wire239) >>> $unsigned(wire238)))));
              reg258 <= $unsigned($unsigned($unsigned(reg256)));
            end
          else
            begin
              reg255 <= $signed((&(~|reg251)));
              reg256 <= wire239[(1'h1):(1'h1)];
              reg258 <= ((~$unsigned({reg251})) ?
                  (!wire239) : reg250[(2'h3):(2'h3)]);
            end
          reg259 <= reg255[(2'h2):(1'h0)];
          for (forvar260 = (1'h0); (forvar260 < (2'h3)); forvar260 = (forvar260 + (1'h1)))
            begin
              reg261 <= {((8'ha9) ? {$unsigned(wire238)} : (8'ha9))};
              reg262 <= $signed($signed((reg251[(3'h5):(2'h2)] ?
                  (|$unsigned(reg253)) : $unsigned($signed(reg258)))));
              reg263 <= reg257[(4'ha):(3'h7)];
            end
        end
      else
        begin
          reg252 = (^~(8'hb4));
          reg253 = ($unsigned(((^~(wire243 ?
              (8'haf) : reg259)) < wire238)) - ((($signed((8'ha7)) >> $signed(reg253)) - (8'hb5)) ?
              reg255[(1'h0):(1'h0)] : $signed((reg250[(4'hb):(3'h6)] <= (|forvar260)))));
          reg255 <= $unsigned($unsigned($signed((|reg261))));
          if (($unsigned((((-reg263) ?
                  $unsigned(reg263) : (wire242 ^ (8'ha0))) ~^ reg262[(5'h11):(4'hc)])) ?
              (^~reg261) : $signed(reg255[(2'h2):(2'h2)])))
            begin
              reg257 = {(7'h47)};
              reg258 <= (reg261 || $unsigned(reg257));
              reg259 <= (reg256[(3'h5):(3'h5)] <= $signed((wire240 ?
                  forvar245[(3'h5):(1'h0)] : $signed((-reg258)))));
              reg260 = $signed($unsigned((7'h43)));
              reg261 <= $signed($signed(((reg260 ~^ reg247) > $signed((reg258 ?
                  reg246 : reg249)))));
            end
          else
            begin
              reg257 = (reg247[(4'h8):(3'h4)] - $unsigned($signed({reg247,
                  $unsigned((8'hae))})));
              reg260 = (8'hae);
              reg261 <= reg263[(3'h7):(2'h3)];
            end
        end
      reg264 <= ($signed((wire242[(2'h2):(1'h1)] ? wire242 : (8'h9d))) ?
          (8'ha3) : $signed((~^(reg251[(3'h7):(1'h1)] ?
              (!reg251) : (wire240 || wire243)))));
      if ($unsigned(reg262[(3'h5):(1'h1)]))
        begin
          reg265 <= ($signed(((+(wire242 ? (7'h45) : reg246)) >= ({reg248,
                  wire242} ?
              $signed(reg251) : ((8'ha7) ?
                  reg257 : (8'hac))))) == reg247[(1'h0):(1'h0)]);
          reg266 <= {wire240[(2'h3):(1'h1)],
              ($signed(((8'hbe) | reg254[(1'h1):(1'h1)])) - wire242)};
          reg267 <= ((($unsigned({reg249, reg264}) ?
              (^~((7'h43) ?
                  reg253 : reg259)) : reg249[(4'hc):(4'hc)]) >> {reg260}) <<< (((+(reg251 ?
                      reg250 : reg258)) ?
                  ((wire243 ? reg264 : (8'had)) ?
                      (reg246 >= wire243) : $signed((7'h43))) : $unsigned($unsigned((8'ha0)))) ?
              (((reg266 >>> reg262) ?
                      (wire240 ? wire238 : reg265) : (reg259 ?
                          wire238 : wire238)) ?
                  (~&(^~wire240)) : reg263[(1'h0):(1'h0)]) : $unsigned(reg257[(1'h1):(1'h1)])));
          for (forvar268 = (1'h0); (forvar268 < (3'h4)); forvar268 = (forvar268 + (1'h1)))
            begin
              reg269 = reg252;
              reg270 = $signed(reg247[(4'h9):(1'h0)]);
              reg271 <= $unsigned(($signed(wire242) >>> reg246));
              reg272 = (+{$signed((7'h43))});
            end
        end
      else
        begin
          reg265 <= {$signed($unsigned($unsigned($signed(reg271)))),
              $unsigned(wire238[(4'hd):(4'h8)])};
        end
    end
  assign wire273 = ((^~{($unsigned(wire238) ?
                               $signed(reg271) : (reg259 ? reg246 : reg265))}) ?
                       (7'h47) : reg267[(4'hb):(4'ha)]);
  always
    @(posedge clk) begin
      reg274 <= reg259;
      reg275 = $signed((reg263 >= (^$unsigned({reg259, (7'h42)}))));
      for (forvar276 = (1'h0); (forvar276 < (1'h0)); forvar276 = (forvar276 + (1'h1)))
        begin
          if (forvar276)
            begin
              reg277 = ((((reg275 ? (^~wire244) : {(7'h44), reg275}) ?
                  wire273 : reg263) | reg271) - ((((^wire239) <<< (~|wire244)) ?
                  ((~|reg264) ?
                      reg261 : (+reg261)) : (8'hb1)) << $unsigned(({wire244,
                      wire240} ?
                  $unsigned(reg250) : reg258))));
              reg278 = (reg275 != $signed($unsigned({(reg258 ?
                      (8'hb4) : reg275),
                  (|reg265)})));
            end
          else
            begin
              reg279 <= wire242[(3'h7):(1'h0)];
              reg280 <= ((8'hbc) >> $signed((~|(-$unsigned(wire273)))));
            end
        end
      reg281 <= (^($unsigned($unsigned((~reg279))) ?
          ($signed($signed(reg263)) ?
              wire241[(4'ha):(2'h3)] : $unsigned(wire239[(3'h6):(3'h6)])) : ($signed(reg267) ?
              {(reg251 - reg264)} : ({reg264} ?
                  (wire273 >= reg271) : $unsigned(reg266)))));
      reg282 <= $signed(reg248[(5'h11):(4'ha)]);
    end
  assign wire283 = $unsigned(wire239[(3'h7):(3'h7)]);
  assign wire284 = $unsigned(wire244);
  always
    @(posedge clk) begin
      if (wire244)
        begin
          if ((~reg250))
            begin
              reg285 = ((wire239 ^ (7'h4a)) ?
                  reg251[(3'h7):(3'h6)] : $signed((~&wire283)));
            end
          else
            begin
              reg285 = {$signed((((wire239 > reg281) <= reg280[(1'h0):(1'h0)]) ?
                      (~&wire244) : reg246)),
                  reg282[(5'h18):(5'h11)]};
            end
          reg286 <= $unsigned(wire284);
          reg287 = $unsigned(wire273);
        end
      else
        begin
          reg285 = (8'hb2);
        end
    end
  assign wire288 = $signed($signed(($unsigned((|reg274)) + ({wire239} + (~^reg279)))));
  always
    @(posedge clk) begin
      for (forvar289 = (1'h0); (forvar289 < (2'h2)); forvar289 = (forvar289 + (1'h1)))
        begin
          reg290 = $unsigned(reg259[(3'h6):(3'h5)]);
          if ((+$signed(wire243)))
            begin
              reg291 <= $signed((+{reg264}));
              reg292 <= ((~|(((7'h48) > ((7'h45) ? wire238 : wire288)) ?
                      reg265[(2'h3):(2'h3)] : (wire273[(5'h12):(4'hb)] != (reg261 ?
                          reg267 : reg282)))) ?
                  wire238[(3'h7):(3'h5)] : (reg246 + $signed(($unsigned(reg264) >> $unsigned(wire238)))));
              reg293 = $unsigned($unsigned((+$signed(reg286[(4'hc):(3'h7)]))));
              reg294 <= wire243[(1'h1):(1'h1)];
              reg295 = $unsigned((wire242 ?
                  {wire241,
                      {reg248[(4'ha):(2'h3)],
                          wire283}} : ($unsigned($signed(reg280)) <<< (8'hbd))));
            end
          else
            begin
              reg293 = $unsigned($signed($unsigned(reg264)));
              reg295 = (8'h9e);
              reg296 = reg267[(4'hb):(4'h8)];
              reg297 <= (&$unsigned(($signed((reg274 ? reg286 : reg295)) ?
                  $unsigned($unsigned(reg255)) : (reg262 ?
                      ((8'hb6) ? reg248 : reg292) : (!reg274)))));
              reg298 <= $unsigned(((~^($signed(reg294) ~^ reg264)) & reg282));
            end
          if ($signed(reg274[(4'h9):(3'h4)]))
            begin
              reg299 = $unsigned((7'h48));
              reg300 = reg271[(1'h0):(1'h0)];
              reg301 = (reg291[(2'h2):(1'h0)] * wire243[(4'h9):(4'h9)]);
            end
          else
            begin
              reg302 <= ((wire240 ?
                  (reg258 ?
                      (((8'hbc) ?
                          reg256 : reg295) <<< {reg279}) : reg296) : ((8'hba) ?
                      wire273[(4'he):(2'h2)] : $unsigned($unsigned(wire283)))) + (7'h49));
              reg303 <= {$unsigned(wire243)};
              reg304 <= (reg302[(4'hc):(3'h4)] ?
                  ($unsigned((reg281 ? reg280 : reg290)) <<< {(8'hbe),
                      (reg280[(5'h13):(2'h3)] ?
                          reg295 : $unsigned(reg301))}) : ($unsigned($signed((reg281 * wire288))) ?
                      wire283[(3'h7):(3'h7)] : (((reg280 ? reg259 : reg261) ?
                          $unsigned(reg251) : (-reg297)) | wire283[(5'h17):(5'h11)])));
              reg305 <= wire240;
              reg306 <= (8'h9f);
            end
          reg307 <= reg282;
        end
      for (forvar308 = (1'h0); (forvar308 < (2'h3)); forvar308 = (forvar308 + (1'h1)))
        begin
          reg309 = ({$unsigned(($signed(reg282) ?
                  (|reg305) : (+(8'hb3))))} >> (reg299 ?
              (^$signed(reg293)) : (~^$signed({reg265}))));
          reg310 <= $unsigned($unsigned((($signed(wire284) >= reg299[(4'hc):(1'h1)]) >> reg305)));
          reg311 <= reg290;
          if ($unsigned((~|reg263[(4'ha):(4'h8)])))
            begin
              reg312 <= (~^reg302[(3'h5):(2'h2)]);
              reg313 = $unsigned(wire288);
            end
          else
            begin
              reg313 = {($signed(reg255) && reg301[(4'hb):(3'h6)]),
                  reg310[(1'h1):(1'h0)]};
            end
          if ($signed((!$signed({(reg264 ? reg250 : reg246)}))))
            begin
              reg314 = (~reg303);
              reg315 = ($unsigned(reg250) - $unsigned((~^((^~reg264) != (wire241 ?
                  reg266 : wire239)))));
              reg316 = (&reg258[(4'hb):(4'hb)]);
              reg317 = $signed($signed({($signed(reg304) * $unsigned((8'hb4))),
                  ((-(7'h40)) - reg282)}));
              reg318 = (reg298 * (wire240[(1'h1):(1'h1)] ~^ (wire238 ?
                  (~|((8'hae) ?
                      reg290 : reg265)) : $signed($unsigned(reg267)))));
            end
          else
            begin
              reg319 <= (reg250 ?
                  {((8'hb0) ? (~|{reg318}) : (reg280 + reg251[(1'h1):(1'h1)])),
                      reg251[(3'h7):(3'h7)]} : $signed((((reg309 || wire273) ?
                          {reg246} : (^reg315)) ?
                      wire273[(1'h1):(1'h1)] : {$signed(reg292),
                          $signed(reg304)})));
            end
        end
    end
  assign wire320 = ($unsigned($unsigned(({reg291, reg306} ?
                       $signed(reg258) : reg248[(1'h0):(1'h0)]))) <<< {(reg294 | (!$signed(reg266))),
                       $unsigned((~^$unsigned(reg302)))});
  assign wire321 = {reg266};
  always
    @(posedge clk) begin
      reg322 <= (!reg267);
      for (forvar323 = (1'h0); (forvar323 < (1'h1)); forvar323 = (forvar323 + (1'h1)))
        begin
          if ($signed($signed((^($unsigned(wire243) ?
              (reg264 ? reg305 : wire243) : forvar323)))))
            begin
              reg324 = $unsigned($unsigned(reg249[(4'h8):(3'h5)]));
            end
          else
            begin
              reg325 <= wire242;
              reg326 <= $unsigned($signed((~|$unsigned((reg255 ?
                  (8'h9d) : reg292)))));
              reg327 <= ((reg298 >>> reg307) ?
                  reg302[(4'he):(4'hd)] : (!reg248[(4'ha):(3'h7)]));
              reg328 = $signed(($unsigned($unsigned((|reg249))) + reg310));
            end
        end
      reg329 <= $unsigned((^$signed(wire273[(3'h6):(3'h4)])));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module852  (y, clk, wire853, wire854, wire855, wire856);
  output wire [(32'hbb9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire853;
  input wire signed [(5'h11):(1'h0)] wire854;
  input wire [(5'h17):(1'h0)] wire855;
  input wire [(5'h14):(1'h0)] wire856;
  wire [(5'h13):(1'h0)] wire1593;
  wire signed [(5'h17):(1'h0)] wire1556;
  wire signed [(2'h2):(1'h0)] wire1553;
  wire signed [(4'h9):(1'h0)] wire1550;
  wire [(5'h12):(1'h0)] wire1303;
  wire [(5'h18):(1'h0)] wire1057;
  wire signed [(4'h8):(1'h0)] wire1090;
  wire signed [(5'h16):(1'h0)] wire1091;
  wire [(4'ha):(1'h0)] wire1092;
  wire [(3'h5):(1'h0)] wire1093;
  wire signed [(5'h15):(1'h0)] wire1094;
  wire signed [(4'he):(1'h0)] wire1095;
  wire [(5'h16):(1'h0)] wire1290;
  reg signed [(3'h5):(1'h0)] reg1576 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1592 = (1'h0);
  reg [(2'h3):(1'h0)] reg1590 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1589 = (1'h0);
  reg [(3'h7):(1'h0)] reg1586 = (1'h0);
  reg [(5'h11):(1'h0)] reg1584 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1578 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1577 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1573 = (1'h0);
  reg [(5'h13):(1'h0)] reg1572 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1570 = (1'h0);
  reg [(4'hb):(1'h0)] reg1567 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1566 = (1'h0);
  reg [(5'h12):(1'h0)] reg1564 = (1'h0);
  reg [(3'h5):(1'h0)] reg1562 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1561 = (1'h0);
  reg [(4'h9):(1'h0)] reg1559 = (1'h0);
  reg [(2'h3):(1'h0)] reg1557 = (1'h0);
  reg [(5'h14):(1'h0)] reg1314 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1313 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1311 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1309 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1306 = (1'h0);
  reg [(5'h17):(1'h0)] reg1301 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1299 = (1'h0);
  reg [(4'hf):(1'h0)] reg1298 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1295 = (1'h0);
  reg [(4'hf):(1'h0)] reg1293 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1217 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1213 = (1'h0);
  reg [(4'he):(1'h0)] reg1209 = (1'h0);
  reg [(3'h6):(1'h0)] reg1203 = (1'h0);
  reg [(3'h6):(1'h0)] reg1201 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1199 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1195 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1193 = (1'h0);
  reg [(4'ha):(1'h0)] reg1187 = (1'h0);
  reg [(3'h7):(1'h0)] reg1186 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1183 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1179 = (1'h0);
  reg [(4'hf):(1'h0)] reg1178 = (1'h0);
  reg [(4'ha):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1173 = (1'h0);
  reg [(5'h11):(1'h0)] reg1172 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1168 = (1'h0);
  reg [(4'ha):(1'h0)] reg1166 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1163 = (1'h0);
  reg [(5'h11):(1'h0)] reg1157 = (1'h0);
  reg [(4'ha):(1'h0)] reg1156 = (1'h0);
  reg [(4'h9):(1'h0)] reg1153 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1150 = (1'h0);
  reg [(5'h13):(1'h0)] reg1148 = (1'h0);
  reg [(4'he):(1'h0)] reg1146 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1142 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1141 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1125 = (1'h0);
  reg [(3'h7):(1'h0)] reg1135 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1133 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1132 = (1'h0);
  reg [(2'h2):(1'h0)] reg1129 = (1'h0);
  reg [(3'h7):(1'h0)] reg1128 = (1'h0);
  reg [(4'hb):(1'h0)] reg1126 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1118 = (1'h0);
  reg [(3'h5):(1'h0)] reg1116 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1114 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1113 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1112 = (1'h0);
  reg [(5'h14):(1'h0)] reg1110 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1109 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1108 = (1'h0);
  reg [(3'h4):(1'h0)] reg1107 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1104 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1100 = (1'h0);
  reg [(3'h5):(1'h0)] reg1099 = (1'h0);
  reg [(4'hb):(1'h0)] reg1089 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1085 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1082 = (1'h0);
  reg [(4'hd):(1'h0)] reg1081 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1078 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1076 = (1'h0);
  reg [(5'h17):(1'h0)] reg1075 = (1'h0);
  reg [(5'h18):(1'h0)] reg1071 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1068 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1067 = (1'h0);
  reg [(5'h14):(1'h0)] reg1065 = (1'h0);
  reg [(5'h17):(1'h0)] reg1064 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1062 = (1'h0);
  reg [(3'h7):(1'h0)] reg1061 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1585 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1591 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1588 = (1'h0);
  reg [(5'h13):(1'h0)] reg1587 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1585 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1583 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1582 = (1'h0);
  reg [(5'h11):(1'h0)] reg1581 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1580 = (1'h0);
  reg [(3'h5):(1'h0)] reg1579 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1576 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1575 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1574 = (1'h0);
  reg [(4'ha):(1'h0)] reg1571 = (1'h0);
  reg [(4'h9):(1'h0)] reg1569 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1568 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1565 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1563 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1560 = (1'h0);
  reg [(4'he):(1'h0)] reg1558 = (1'h0);
  reg [(5'h14):(1'h0)] reg1555 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1554 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1552 = (1'h0);
  reg [(3'h6):(1'h0)] reg1316 = (1'h0);
  reg [(4'hb):(1'h0)] reg1315 = (1'h0);
  reg [(5'h12):(1'h0)] reg1312 = (1'h0);
  reg [(5'h15):(1'h0)] reg1310 = (1'h0);
  reg [(4'hc):(1'h0)] reg1308 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1307 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1305 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1304 = (1'h0);
  reg [(4'hf):(1'h0)] reg1302 = (1'h0);
  reg [(5'h15):(1'h0)] reg1300 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1297 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1292 = (1'h0);
  reg [(5'h16):(1'h0)] reg1296 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1294 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1292 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1216 = (1'h0);
  reg [(2'h2):(1'h0)] reg1215 = (1'h0);
  reg [(4'h8):(1'h0)] reg1214 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1212 = (1'h0);
  reg [(3'h4):(1'h0)] reg1211 = (1'h0);
  reg [(4'hd):(1'h0)] reg1210 = (1'h0);
  reg [(3'h7):(1'h0)] reg1208 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1207 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1206 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1205 = (1'h0);
  reg [(5'h10):(1'h0)] reg1204 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1202 = (1'h0);
  reg [(2'h3):(1'h0)] reg1200 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1198 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1197 = (1'h0);
  reg [(4'h9):(1'h0)] reg1196 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1194 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1192 = (1'h0);
  reg [(3'h5):(1'h0)] reg1191 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1190 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1189 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1188 = (1'h0);
  reg [(4'he):(1'h0)] reg1185 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1184 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1182 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1181 = (1'h0);
  reg [(5'h11):(1'h0)] reg1180 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1177 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1175 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1174 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1166 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1171 = (1'h0);
  reg [(3'h5):(1'h0)] reg1170 = (1'h0);
  reg [(4'h8):(1'h0)] reg1169 = (1'h0);
  reg [(4'he):(1'h0)] reg1167 = (1'h0);
  reg [(4'hd):(1'h0)] reg1144 = (1'h0);
  reg [(4'hb):(1'h0)] reg1165 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1164 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1162 = (1'h0);
  reg [(4'hf):(1'h0)] reg1161 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1160 = (1'h0);
  reg [(4'ha):(1'h0)] reg1159 = (1'h0);
  reg [(5'h13):(1'h0)] reg1158 = (1'h0);
  reg [(3'h4):(1'h0)] reg1155 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1154 = (1'h0);
  reg [(5'h11):(1'h0)] reg1152 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1151 = (1'h0);
  reg [(4'h8):(1'h0)] reg1149 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1147 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1145 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1144 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1143 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1140 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1139 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1138 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1126 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1137 = (1'h0);
  reg [(4'hd):(1'h0)] reg1136 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1134 = (1'h0);
  reg [(4'hd):(1'h0)] reg1131 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1130 = (1'h0);
  reg [(4'ha):(1'h0)] reg1127 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1125 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1124 = (1'h0);
  reg [(5'h13):(1'h0)] reg1123 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1122 = (1'h0);
  reg [(4'hc):(1'h0)] reg1121 = (1'h0);
  reg [(5'h12):(1'h0)] reg1120 = (1'h0);
  reg [(4'hc):(1'h0)] reg1119 = (1'h0);
  reg [(5'h17):(1'h0)] reg1117 = (1'h0);
  reg [(3'h7):(1'h0)] reg1115 = (1'h0);
  reg [(4'h9):(1'h0)] reg1111 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1106 = (1'h0);
  reg [(4'hd):(1'h0)] reg1105 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1103 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1102 = (1'h0);
  reg [(4'h9):(1'h0)] reg1101 = (1'h0);
  reg [(4'hc):(1'h0)] reg1098 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1097 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1096 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1088 = (1'h0);
  reg [(4'he):(1'h0)] reg1087 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1086 = (1'h0);
  reg [(4'hf):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1083 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1080 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1079 = (1'h0);
  reg [(2'h2):(1'h0)] reg1077 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1074 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1073 = (1'h0);
  reg [(2'h3):(1'h0)] reg1072 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1070 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1069 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1066 = (1'h0);
  reg [(3'h7):(1'h0)] reg1063 = (1'h0);
  reg [(5'h17):(1'h0)] reg1060 = (1'h0);
  reg [(5'h14):(1'h0)] reg1059 = (1'h0);
  assign y = {wire1593,
                 wire1556,
                 wire1553,
                 wire1550,
                 wire1303,
                 wire1057,
                 wire1090,
                 wire1091,
                 wire1092,
                 wire1093,
                 wire1094,
                 wire1095,
                 wire1290,
                 reg1576,
                 reg1592,
                 reg1590,
                 reg1589,
                 reg1586,
                 reg1584,
                 reg1578,
                 reg1577,
                 reg1573,
                 reg1572,
                 reg1570,
                 reg1567,
                 reg1566,
                 reg1564,
                 reg1562,
                 reg1561,
                 reg1559,
                 reg1557,
                 reg1314,
                 reg1313,
                 reg1311,
                 reg1309,
                 reg1306,
                 reg1301,
                 reg1299,
                 reg1298,
                 reg1295,
                 reg1293,
                 reg1217,
                 reg1213,
                 reg1209,
                 reg1203,
                 reg1201,
                 reg1199,
                 reg1195,
                 reg1193,
                 reg1187,
                 reg1186,
                 reg1183,
                 reg1179,
                 reg1178,
                 reg1176,
                 reg1173,
                 reg1172,
                 reg1168,
                 reg1166,
                 reg1163,
                 reg1157,
                 reg1156,
                 reg1153,
                 reg1150,
                 reg1148,
                 reg1146,
                 reg1142,
                 reg1141,
                 reg1125,
                 reg1135,
                 reg1133,
                 reg1132,
                 reg1129,
                 reg1128,
                 reg1126,
                 reg1118,
                 reg1116,
                 reg1114,
                 reg1113,
                 reg1112,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1107,
                 reg1104,
                 reg1100,
                 reg1099,
                 reg1089,
                 reg1085,
                 reg1082,
                 reg1081,
                 reg1078,
                 reg1076,
                 reg1075,
                 reg1071,
                 reg1068,
                 reg1067,
                 reg1065,
                 reg1064,
                 reg1062,
                 reg1061,
                 forvar1585,
                 reg1591,
                 reg1588,
                 reg1587,
                 reg1585,
                 reg1583,
                 reg1582,
                 reg1581,
                 reg1580,
                 reg1579,
                 forvar1576,
                 reg1575,
                 reg1574,
                 reg1571,
                 reg1569,
                 reg1568,
                 reg1565,
                 reg1563,
                 reg1560,
                 reg1558,
                 reg1555,
                 reg1554,
                 reg1552,
                 reg1316,
                 reg1315,
                 reg1312,
                 reg1310,
                 reg1308,
                 reg1307,
                 forvar1305,
                 forvar1304,
                 reg1302,
                 reg1300,
                 forvar1297,
                 forvar1292,
                 reg1296,
                 reg1294,
                 reg1292,
                 reg1216,
                 reg1215,
                 reg1214,
                 forvar1212,
                 reg1211,
                 reg1210,
                 reg1208,
                 forvar1207,
                 reg1206,
                 reg1205,
                 reg1204,
                 reg1202,
                 reg1200,
                 forvar1198,
                 reg1197,
                 reg1196,
                 reg1194,
                 reg1192,
                 reg1191,
                 reg1190,
                 reg1189,
                 reg1188,
                 reg1185,
                 forvar1184,
                 forvar1182,
                 forvar1181,
                 reg1180,
                 reg1177,
                 reg1175,
                 forvar1174,
                 forvar1166,
                 reg1171,
                 reg1170,
                 reg1169,
                 reg1167,
                 reg1144,
                 reg1165,
                 reg1164,
                 reg1162,
                 reg1161,
                 forvar1160,
                 reg1159,
                 reg1158,
                 reg1155,
                 reg1154,
                 reg1152,
                 reg1151,
                 reg1149,
                 reg1147,
                 reg1145,
                 forvar1144,
                 reg1143,
                 reg1140,
                 reg1139,
                 forvar1138,
                 forvar1126,
                 reg1137,
                 reg1136,
                 reg1134,
                 reg1131,
                 reg1130,
                 reg1127,
                 forvar1125,
                 reg1124,
                 reg1123,
                 forvar1122,
                 reg1121,
                 reg1120,
                 reg1119,
                 reg1117,
                 reg1115,
                 reg1111,
                 reg1106,
                 reg1105,
                 reg1103,
                 reg1102,
                 reg1101,
                 reg1098,
                 forvar1097,
                 reg1096,
                 reg1088,
                 reg1087,
                 reg1086,
                 reg1084,
                 reg1083,
                 forvar1080,
                 forvar1079,
                 reg1077,
                 forvar1074,
                 reg1073,
                 reg1072,
                 reg1070,
                 forvar1069,
                 forvar1066,
                 reg1063,
                 reg1060,
                 reg1059,
                 (1'h0)};
  module857 #() modinst1058 (.wire858(wire855), .y(wire1057), .wire860(wire856), .wire861(wire853), .wire859(wire854), .clk(clk));
  always
    @(posedge clk) begin
      reg1059 = ($unsigned(({((8'hb9) * wire853)} ?
          wire853 : (7'h40))) <<< $unsigned((wire854 <<< wire855)));
      if ((^(~^$signed($signed({wire855, (8'ha3)})))))
        begin
          reg1060 = {wire854[(4'hc):(4'h8)]};
          reg1061 <= ((($signed((wire855 < wire854)) ?
              $unsigned($signed(reg1059)) : (8'hb0)) > wire853[(2'h2):(1'h1)]) != wire854);
          reg1062 <= (~&wire854[(3'h5):(2'h3)]);
        end
      else
        begin
          if (wire1057[(5'h15):(5'h12)])
            begin
              reg1060 = $signed(((wire854 ?
                      (~^$unsigned(reg1059)) : (reg1060[(5'h12):(1'h1)] >> $unsigned(wire854))) ?
                  $unsigned(((reg1060 ? wire1057 : (8'h9f)) ?
                      reg1062 : $signed(wire1057))) : ($unsigned($signed(reg1061)) >> (((8'hbc) <= reg1062) == $unsigned(wire854)))));
              reg1063 = reg1060[(4'h8):(3'h6)];
              reg1064 <= wire855[(4'h8):(1'h0)];
            end
          else
            begin
              reg1061 <= $unsigned(wire1057);
              reg1062 <= $unsigned($signed((~|{(wire855 ^ wire855),
                  wire855[(5'h14):(3'h6)]})));
              reg1064 <= ((wire854 ?
                  $signed((^reg1062[(3'h6):(3'h6)])) : ($unsigned((reg1062 >>> (7'h4a))) ?
                      wire854 : {(wire854 ?
                              wire1057 : reg1063)})) > ($signed((-wire1057)) <<< reg1059[(3'h4):(1'h0)]));
              reg1065 <= $unsigned(reg1061[(3'h4):(2'h2)]);
            end
          for (forvar1066 = (1'h0); (forvar1066 < (2'h2)); forvar1066 = (forvar1066 + (1'h1)))
            begin
              reg1067 <= reg1064[(5'h10):(1'h1)];
              reg1068 <= wire855;
            end
          for (forvar1069 = (1'h0); (forvar1069 < (2'h3)); forvar1069 = (forvar1069 + (1'h1)))
            begin
              reg1070 = $unsigned((reg1063[(2'h2):(1'h0)] ?
                  {(&wire1057[(3'h6):(3'h5)]),
                      (wire853[(3'h6):(3'h4)] ^~ (wire854 >= reg1060))} : reg1065));
              reg1071 <= reg1067[(4'h8):(3'h7)];
              reg1072 = wire1057;
            end
          reg1073 = ((&(&($signed(wire1057) ?
              ((8'hb7) ?
                  wire856 : wire854) : wire853))) >= $signed(reg1059[(4'hf):(3'h6)]));
          for (forvar1074 = (1'h0); (forvar1074 < (1'h0)); forvar1074 = (forvar1074 + (1'h1)))
            begin
              reg1075 <= $signed($unsigned(reg1061));
              reg1076 <= {($signed(reg1067) ^~ (((forvar1066 || wire856) >= (forvar1074 <<< reg1067)) >= ((reg1059 + reg1073) ?
                      reg1063[(3'h6):(1'h0)] : (~|wire856))))};
            end
        end
      reg1077 = (reg1059 ?
          $unsigned($unsigned($signed({reg1073}))) : (forvar1069 * $unsigned(((wire853 ?
              reg1067 : reg1071) == reg1068[(3'h4):(1'h0)]))));
    end
  always
    @(posedge clk) begin
      reg1078 <= $unsigned(reg1065);
      for (forvar1079 = (1'h0); (forvar1079 < (1'h0)); forvar1079 = (forvar1079 + (1'h1)))
        begin
          for (forvar1080 = (1'h0); (forvar1080 < (1'h1)); forvar1080 = (forvar1080 + (1'h1)))
            begin
              reg1081 <= (~|{{(reg1078 | reg1065)},
                  (($signed(reg1067) ~^ (wire1057 ^~ reg1068)) || (^wire1057))});
              reg1082 <= (~&(((-forvar1079[(4'hc):(3'h7)]) + wire1057) ~^ ((reg1076 + $unsigned(reg1071)) >> $unsigned((^forvar1080)))));
              reg1083 = (8'hae);
              reg1084 = {forvar1079,
                  $unsigned({$signed($unsigned(reg1065)), wire853})};
            end
          if ($signed(((-$unsigned(reg1078)) ?
              (wire855[(5'h15):(4'h9)] >= reg1064) : $unsigned($unsigned(reg1075[(5'h14):(3'h6)])))))
            begin
              reg1085 <= (reg1081[(3'h7):(1'h0)] ?
                  $unsigned($signed($signed((forvar1079 ?
                      (8'ha6) : wire853)))) : $unsigned($signed($unsigned($signed(wire854)))));
            end
          else
            begin
              reg1086 = reg1082[(1'h1):(1'h0)];
              reg1087 = (&$signed(reg1061[(2'h3):(2'h3)]));
              reg1088 = (-$unsigned((~^((reg1086 ?
                  (8'hab) : reg1082) | (~reg1067)))));
            end
        end
      reg1089 <= ({reg1076[(5'h12):(5'h12)]} >>> $signed((!$unsigned((~|wire854)))));
    end
  assign wire1090 = ((reg1075[(4'hd):(4'ha)] == (~((~|reg1076) + reg1075[(4'hc):(2'h2)]))) || {((wire1057 ?
                                (reg1081 ?
                                    reg1067 : reg1081) : reg1078[(3'h5):(1'h1)]) ?
                            (~reg1061) : (^reg1076))});
  assign wire1091 = reg1064;
  assign wire1092 = $signed({$unsigned(reg1065[(4'ha):(3'h4)])});
  assign wire1093 = $signed($unsigned($unsigned(({wire855, (7'h48)} ?
                        (+(8'hb7)) : (reg1065 ? reg1062 : wire1092)))));
  assign wire1094 = $signed(((^~reg1065) < ((wire856 ?
                        wire1092 : $unsigned(reg1082)) * (8'h9e))));
  assign wire1095 = (8'hbf);
  always
    @(posedge clk) begin
      reg1096 = (reg1064[(5'h17):(2'h2)] | ({wire855[(4'ha):(1'h0)]} >= $signed((wire1092[(4'h9):(3'h7)] ?
          $unsigned(reg1078) : $signed(reg1089)))));
      for (forvar1097 = (1'h0); (forvar1097 < (3'h4)); forvar1097 = (forvar1097 + (1'h1)))
        begin
          reg1098 = reg1067;
          reg1099 <= $signed(wire1091);
          reg1100 <= $signed($unsigned({reg1062}));
          reg1101 = (~wire1057[(3'h4):(1'h1)]);
          if ($signed($unsigned((~^({reg1085, reg1085} ?
              (|reg1082) : (^~wire1091))))))
            begin
              reg1102 = $signed($unsigned($unsigned(reg1075)));
              reg1103 = (7'h46);
              reg1104 <= (!$signed(($signed(reg1103[(1'h0):(1'h0)]) != $unsigned($signed(wire856)))));
              reg1105 = reg1098[(4'ha):(3'h6)];
            end
          else
            begin
              reg1104 <= reg1081[(4'hb):(4'ha)];
              reg1105 = reg1104[(4'he):(4'hb)];
              reg1106 = $signed(reg1089[(4'h8):(3'h5)]);
            end
        end
      if ($signed(reg1078[(5'h17):(4'hd)]))
        begin
          reg1107 <= ($unsigned($signed(($unsigned(wire1094) << (reg1096 ?
                  reg1076 : wire1057)))) ?
              reg1065 : wire853[(4'hb):(3'h6)]);
          reg1108 <= ({$signed(reg1081[(4'ha):(3'h7)]),
                  $signed({(reg1075 >= reg1075)})} ?
              $unsigned(reg1098) : wire1090);
          reg1109 <= (!forvar1097[(2'h3):(1'h1)]);
          reg1110 <= ($signed(($signed((^reg1098)) ?
                  wire853 : (wire1092 ? {reg1108} : $signed(wire1093)))) ?
              $unsigned(reg1096) : {$unsigned($unsigned((reg1081 ^~ reg1106))),
                  wire1094});
        end
      else
        begin
          if ((~$signed(((&{reg1109}) ?
              $signed(reg1067[(4'h8):(2'h2)]) : reg1105[(1'h1):(1'h1)]))))
            begin
              reg1111 = (reg1102 && reg1099);
              reg1112 <= (&{$unsigned(({(8'h9e), wire1092} - reg1064))});
              reg1113 <= $signed(wire856);
              reg1114 <= {(^(wire855[(4'he):(3'h5)] ?
                      $unsigned($unsigned((8'ha8))) : $signed(reg1062[(3'h7):(3'h5)]))),
                  ($signed({(~&reg1068)}) <= wire853)};
              reg1115 = $unsigned(reg1068[(1'h0):(1'h0)]);
            end
          else
            begin
              reg1107 <= (!((($unsigned(wire1092) + (reg1099 <<< wire1091)) ?
                      reg1100 : (^((8'h9d) * reg1111))) ?
                  reg1104 : reg1113[(4'he):(4'hc)]));
            end
          reg1116 <= (reg1104[(4'hb):(4'h8)] & ($unsigned(reg1103[(3'h4):(2'h3)]) ?
              ((8'h9d) >>> $unsigned((!(8'hb0)))) : $unsigned(({wire1092} ?
                  {reg1113, (7'h41)} : $signed(wire856)))));
          reg1117 = $signed($signed(($unsigned(reg1068) - wire1090)));
          reg1118 <= $unsigned($signed(($unsigned($signed(reg1112)) * ($unsigned(wire1093) ?
              reg1115 : (-(7'h43))))));
          reg1119 = $unsigned(wire1090);
        end
    end
  always
    @(posedge clk) begin
      reg1120 = ((reg1112[(1'h0):(1'h0)] + $unsigned({reg1118,
              $signed(wire853)})) ?
          $signed((~^({reg1116,
              reg1100} <= $unsigned(wire1057)))) : ($unsigned(reg1076[(4'ha):(2'h3)]) * reg1075));
      reg1121 = $signed($signed(($signed(reg1061) ?
          ($unsigned(reg1067) ?
              reg1061 : $unsigned(reg1109)) : (^~(^~wire856)))));
      if (((~^$unsigned(({reg1067, reg1081} >> wire856))) ?
          (~&$unsigned((+(reg1078 ? reg1109 : reg1067)))) : reg1113))
        begin
          for (forvar1122 = (1'h0); (forvar1122 < (2'h2)); forvar1122 = (forvar1122 + (1'h1)))
            begin
              reg1123 = wire1095[(4'he):(3'h4)];
            end
          reg1124 = (reg1118 ?
              ($unsigned((((8'h9c) ? reg1108 : reg1120) ?
                      $unsigned(reg1099) : $unsigned(reg1116))) ?
                  reg1108 : $unsigned((~forvar1122))) : ($signed(($unsigned((7'h47)) >= $signed(reg1085))) && (8'hba)));
          for (forvar1125 = (1'h0); (forvar1125 < (1'h1)); forvar1125 = (forvar1125 + (1'h1)))
            begin
              reg1126 <= (!{reg1081,
                  (((wire1094 && (8'hb8)) > (reg1082 ? (8'hb8) : reg1120)) ?
                      $unsigned((wire1094 + reg1108)) : $signed((wire1095 ^ wire854)))});
              reg1127 = (|(($unsigned(reg1071[(5'h10):(4'h9)]) <<< (+$unsigned(wire853))) ?
                  (reg1078 << reg1076) : wire853[(1'h1):(1'h0)]));
            end
          if (($signed(wire1090[(3'h7):(1'h1)]) || $unsigned((-(~^reg1120)))))
            begin
              reg1128 <= (reg1109 > (~&$signed(reg1061)));
              reg1129 <= (^~{($signed((reg1108 ? reg1128 : reg1064)) ?
                      ($unsigned(forvar1122) ?
                          (reg1085 ?
                              reg1100 : wire853) : $signed(reg1062)) : wire1090)});
              reg1130 = (wire853 ?
                  reg1113[(4'h9):(4'h8)] : $unsigned(($signed(forvar1125) < (~|(reg1124 >> wire1092)))));
              reg1131 = $unsigned((7'h45));
              reg1132 <= (reg1085[(3'h5):(1'h0)] + (-($unsigned(wire1095[(3'h6):(1'h1)]) ~^ (~&$unsigned(wire1092)))));
            end
          else
            begin
              reg1128 <= $signed($signed($unsigned((8'hba))));
              reg1129 <= $unsigned($signed((reg1099 > (&$signed(reg1131)))));
            end
          if ((-(~^reg1107[(1'h0):(1'h0)])))
            begin
              reg1133 <= reg1124;
              reg1134 = $signed((^{(8'hac)}));
              reg1135 <= reg1065;
              reg1136 = ($signed(reg1118[(4'h8):(1'h1)]) == $unsigned($unsigned($signed(reg1135[(2'h2):(1'h1)]))));
              reg1137 = reg1124;
            end
          else
            begin
              reg1133 <= forvar1122[(3'h4):(2'h2)];
            end
        end
      else
        begin
          for (forvar1122 = (1'h0); (forvar1122 < (2'h3)); forvar1122 = (forvar1122 + (1'h1)))
            begin
              reg1125 <= reg1108[(4'h9):(1'h0)];
            end
          for (forvar1126 = (1'h0); (forvar1126 < (1'h0)); forvar1126 = (forvar1126 + (1'h1)))
            begin
              reg1128 <= {((-(!$unsigned(reg1107))) ?
                      {{forvar1126[(4'ha):(4'h8)],
                              (reg1076 ? wire1094 : reg1124)},
                          $signed($unsigned(reg1113))} : reg1130[(1'h0):(1'h0)])};
            end
          reg1130 = $unsigned(wire1093);
        end
    end
  always
    @(posedge clk) begin
      for (forvar1138 = (1'h0); (forvar1138 < (2'h3)); forvar1138 = (forvar1138 + (1'h1)))
        begin
          if ($unsigned((~^(wire1057 ?
              reg1125[(2'h3):(2'h2)] : ((-wire1094) ?
                  $unsigned(wire855) : $unsigned((8'ha8)))))))
            begin
              reg1139 = (reg1062 <= $unsigned((((7'h47) <= $signed(reg1068)) ?
                  reg1099 : {(reg1113 < reg1085)})));
              reg1140 = $signed((!$signed($signed($unsigned(reg1076)))));
              reg1141 <= wire853;
            end
          else
            begin
              reg1141 <= (~&((|(+(wire1095 >>> forvar1138))) ?
                  $signed(reg1068[(2'h3):(2'h2)]) : (($unsigned(wire1094) ~^ (~reg1081)) || $unsigned($signed((8'hbe))))));
              reg1142 <= (+(~|reg1071[(3'h7):(3'h6)]));
              reg1143 = {(&{(8'ha7)})};
            end
        end
      if (($unsigned({reg1065}) ?
          reg1071 : $unsigned($signed((|$signed(reg1082))))))
        begin
          for (forvar1144 = (1'h0); (forvar1144 < (3'h4)); forvar1144 = (forvar1144 + (1'h1)))
            begin
              reg1145 = reg1139;
              reg1146 <= $unsigned({((((8'hb4) << reg1126) ?
                      $unsigned((8'h9f)) : $signed(reg1085)) <= $signed(reg1064[(4'hb):(3'h6)]))});
              reg1147 = $signed($signed({$signed(reg1078[(5'h11):(4'hf)])}));
            end
          if ($signed(reg1099))
            begin
              reg1148 <= $unsigned(reg1062);
              reg1149 = $unsigned($unsigned(reg1132[(1'h1):(1'h1)]));
            end
          else
            begin
              reg1148 <= $unsigned(reg1100[(4'ha):(3'h7)]);
              reg1149 = $signed(wire1094);
              reg1150 <= (reg1100[(4'hf):(4'h9)] ?
                  {reg1081[(3'h7):(1'h0)]} : $unsigned($unsigned($unsigned($signed(reg1112)))));
            end
          if (reg1135)
            begin
              reg1151 = $unsigned($unsigned((({wire854} ?
                      reg1150[(1'h1):(1'h0)] : (reg1071 ? (7'h4a) : reg1116)) ?
                  {reg1133, (reg1067 && wire1090)} : ((reg1064 ?
                      reg1146 : reg1139) != (wire1095 ? reg1068 : (7'h40))))));
              reg1152 = {$signed(reg1061[(1'h1):(1'h0)]),
                  $unsigned((((reg1128 ? reg1081 : reg1128) ?
                          (reg1100 >= reg1128) : $signed(reg1062)) ?
                      (reg1150[(4'h8):(2'h2)] ?
                          reg1145 : $signed((8'hba))) : ($signed(reg1133) ~^ reg1128)))};
              reg1153 <= ({($signed((~|(8'hb8))) ?
                      {$unsigned(reg1065),
                          $signed(reg1149)} : reg1145)} <<< ($unsigned({wire1091,
                      $signed(reg1146)}) ?
                  ((~(reg1132 ? reg1078 : reg1081)) ?
                      reg1075[(5'h17):(4'he)] : (+reg1150[(4'h8):(4'h8)])) : (8'hbc)));
              reg1154 = (((8'ha8) * $unsigned((reg1104[(5'h10):(4'h8)] ?
                      (reg1142 ? wire854 : wire1057) : (|(8'hb4))))) ?
                  (8'h9e) : (^~{$unsigned(((8'hbb) | reg1126)), (~^reg1068)}));
              reg1155 = {(!$signed($unsigned($signed(reg1085)))),
                  forvar1138[(4'hc):(4'h9)]};
            end
          else
            begin
              reg1151 = $signed(reg1118);
              reg1153 <= $unsigned(reg1150[(4'ha):(1'h1)]);
              reg1156 <= {reg1078[(3'h4):(1'h1)]};
              reg1157 <= ((((wire1095[(3'h7):(3'h6)] == reg1142) != $signed(reg1142[(1'h0):(1'h0)])) ^~ $unsigned($signed(reg1116))) ?
                  $signed(reg1143) : reg1128[(3'h7):(1'h0)]);
              reg1158 = (((reg1078 ?
                      {wire1091[(3'h6):(3'h4)],
                          ((8'hba) >> reg1099)} : $signed((8'haa))) & $unsigned($unsigned(reg1078[(5'h14):(2'h2)]))) ?
                  ((8'hbf) ?
                      ({forvar1144,
                          $unsigned(reg1109)} >>> (~(&wire1093))) : {(+$unsigned(wire1094)),
                          ((reg1065 >> reg1114) ?
                              (|reg1139) : $signed(wire1093))}) : (reg1129 & reg1100[(4'h9):(4'h9)]));
            end
          reg1159 = ((((reg1140 ?
                      (~&reg1154) : (reg1158 ^ reg1125)) * $unsigned($unsigned(wire1057))) ?
                  ((wire1095[(1'h0):(1'h0)] < reg1145[(1'h1):(1'h1)]) ?
                      $unsigned($signed((8'hb4))) : ((~^reg1132) ?
                          $signed(reg1109) : $unsigned(reg1071))) : $signed(((&reg1116) << (~^reg1107)))) ?
              wire1091 : $unsigned($unsigned($signed($unsigned((8'ha9))))));
          for (forvar1160 = (1'h0); (forvar1160 < (3'h4)); forvar1160 = (forvar1160 + (1'h1)))
            begin
              reg1161 = {reg1153};
              reg1162 = $signed($unsigned($unsigned((^reg1150))));
              reg1163 <= wire856[(2'h2):(2'h2)];
              reg1164 = $signed({(~|({reg1068, reg1162} && (reg1161 ?
                      reg1075 : wire855)))});
              reg1165 = ((~&((~^$signed(reg1154)) * (!wire1095))) << reg1110[(5'h13):(1'h0)]);
            end
        end
      else
        begin
          if ((|reg1152))
            begin
              reg1144 = (8'ha5);
            end
          else
            begin
              reg1146 <= (reg1085 ?
                  (+({{reg1067}, $unsigned(reg1109)} ?
                      (!(reg1107 != reg1108)) : ((+reg1140) ?
                          reg1151[(4'h8):(1'h1)] : reg1144[(3'h7):(3'h5)]))) : (reg1146[(1'h0):(1'h0)] >>> (($unsigned(reg1157) - (reg1148 ?
                      wire1092 : reg1154)) > $unsigned(wire853[(4'h9):(2'h3)]))));
              reg1147 = ($unsigned(reg1145) != reg1062[(3'h5):(2'h2)]);
              reg1149 = reg1118[(4'ha):(1'h1)];
              reg1150 <= wire854[(3'h6):(1'h0)];
              reg1153 <= forvar1138;
            end
          reg1154 = (reg1081 <<< $signed((($unsigned(reg1132) != (reg1099 - reg1110)) ?
              reg1114 : $signed({reg1140, reg1162}))));
        end
      if ($unsigned($unsigned(reg1148[(2'h3):(1'h0)])))
        begin
          if ($unsigned(forvar1138))
            begin
              reg1166 <= reg1156[(3'h6):(1'h0)];
              reg1167 = $unsigned({$signed(reg1129[(1'h1):(1'h1)]),
                  (((reg1068 ? reg1085 : reg1108) + reg1078) >= (-(wire1057 ?
                      reg1146 : reg1157)))});
              reg1168 <= reg1128;
              reg1169 = reg1164[(1'h0):(1'h0)];
            end
          else
            begin
              reg1166 <= (8'hac);
              reg1167 = (!{reg1071, $signed((~$signed(reg1141)))});
              reg1169 = reg1139[(2'h3):(1'h0)];
              reg1170 = reg1064;
              reg1171 = {$unsigned($unsigned(($signed(reg1152) ?
                      (reg1078 ? reg1061 : reg1169) : (|reg1133)))),
                  (reg1065 ?
                      (-$signed($unsigned((8'hac)))) : ($unsigned((^reg1116)) ?
                          wire854[(1'h1):(1'h0)] : $unsigned(reg1128[(3'h7):(3'h7)])))};
            end
          reg1172 <= forvar1144[(2'h3):(1'h0)];
        end
      else
        begin
          for (forvar1166 = (1'h0); (forvar1166 < (1'h1)); forvar1166 = (forvar1166 + (1'h1)))
            begin
              reg1168 <= (^~reg1129);
              reg1172 <= {$signed(reg1085)};
              reg1173 <= (~^(reg1161 <= (!(wire1094 ?
                  (reg1143 || wire853) : reg1147[(3'h4):(3'h4)]))));
            end
          for (forvar1174 = (1'h0); (forvar1174 < (2'h3)); forvar1174 = (forvar1174 + (1'h1)))
            begin
              reg1175 = $unsigned((^$signed(((~&reg1168) ^~ $signed(forvar1160)))));
              reg1176 <= wire1092;
              reg1177 = {reg1076[(3'h4):(1'h0)], (|(8'hbf))};
              reg1178 <= reg1114;
              reg1179 <= $signed((((^~(^reg1176)) ?
                  $unsigned((reg1158 ?
                      reg1169 : reg1100)) : reg1163) ~^ $signed((-$signed(reg1153)))));
            end
          reg1180 = (^~(~^$signed((reg1065 ? $unsigned(reg1132) : reg1126))));
        end
      for (forvar1181 = (1'h0); (forvar1181 < (1'h1)); forvar1181 = (forvar1181 + (1'h1)))
        begin
          for (forvar1182 = (1'h0); (forvar1182 < (2'h3)); forvar1182 = (forvar1182 + (1'h1)))
            begin
              reg1183 <= reg1154;
            end
        end
      for (forvar1184 = (1'h0); (forvar1184 < (3'h4)); forvar1184 = (forvar1184 + (1'h1)))
        begin
          reg1185 = $signed((({$unsigned(reg1152)} ?
                  $signed(reg1128[(1'h0):(1'h0)]) : {(!reg1108), wire853}) ?
              $signed(reg1089[(2'h3):(2'h3)]) : reg1099));
          reg1186 <= (({($unsigned(reg1161) ? forvar1181 : $signed(reg1173))} ?
              (+(&reg1132)) : $unsigned(reg1104[(4'h8):(3'h6)])) ~^ reg1169);
          reg1187 <= (|forvar1181[(4'hb):(3'h7)]);
        end
    end
  always
    @(posedge clk) begin
      reg1188 = reg1104;
      if ($unsigned($signed(wire1093)))
        begin
          reg1189 = {(|(((~reg1068) ^~ $signed(reg1067)) ?
                  ((8'hbd) + (~|reg1100)) : {reg1157}))};
          reg1190 = (reg1189 - ($signed((|(reg1178 ? reg1183 : reg1110))) ?
              (reg1129 ? reg1188 : reg1075) : reg1173[(1'h0):(1'h0)]));
          reg1191 = reg1157[(4'h9):(2'h2)];
          if ((reg1081 ?
              ($unsigned($unsigned((reg1176 ? reg1071 : reg1191))) ?
                  $signed((~^$signed(reg1062))) : ($unsigned({(8'hb0)}) <= {reg1187[(3'h6):(2'h2)]})) : wire1092[(3'h7):(2'h2)]))
            begin
              reg1192 = reg1168;
            end
          else
            begin
              reg1193 <= $unsigned((!(^~((wire854 & reg1166) ^~ reg1188[(3'h4):(2'h2)]))));
              reg1194 = $signed($unsigned(($unsigned((7'h49)) < $unsigned(reg1067[(4'hd):(4'hc)]))));
              reg1195 <= $unsigned($signed((({reg1065} ?
                  (-reg1178) : (~&reg1193)) < {$unsigned(reg1179),
                  (reg1067 <<< reg1099)})));
              reg1196 = ({reg1141[(4'hd):(4'h9)],
                  reg1089} || reg1062[(2'h3):(1'h0)]);
              reg1197 = {(($signed(reg1150) ?
                          $signed((&(8'hb7))) : {(reg1188 ?
                                  wire856 : reg1191)}) ?
                      ((~reg1146) ?
                          $unsigned($unsigned((8'hb5))) : $signed(reg1082)) : $signed($signed($unsigned(reg1194))))};
            end
        end
      else
        begin
          reg1193 <= $unsigned($signed($signed($signed(reg1081))));
        end
      for (forvar1198 = (1'h0); (forvar1198 < (2'h3)); forvar1198 = (forvar1198 + (1'h1)))
        begin
          reg1199 <= $unsigned({reg1085[(1'h1):(1'h0)],
              $signed($signed($signed(reg1071)))});
        end
      if ((((reg1118 ?
              $unsigned((^wire1095)) : $signed($unsigned(reg1186))) <<< ((reg1109[(5'h12):(4'h8)] != wire853[(2'h3):(2'h2)]) <= reg1141)) ?
          $unsigned($signed(reg1196)) : (reg1100[(1'h0):(1'h0)] > reg1183)))
        begin
          reg1200 = ((|(reg1197[(2'h3):(2'h2)] ?
              $unsigned((reg1100 && reg1132)) : reg1126)) >>> reg1172);
          reg1201 <= ((reg1157[(5'h10):(3'h4)] >>> (~|wire1091[(4'h8):(4'h8)])) <= $signed((!$unsigned((reg1194 + (7'h49))))));
        end
      else
        begin
          if ((-$unsigned($signed(((reg1179 < reg1168) ?
              ((8'h9e) <= wire1090) : (reg1089 ? reg1082 : reg1199))))))
            begin
              reg1201 <= ((-reg1153[(3'h6):(3'h6)]) < ((reg1201[(1'h1):(1'h0)] >>> ((^reg1166) + (8'hb5))) <= ({reg1178,
                  (~reg1068)} < (reg1113 >= $signed(reg1065)))));
              reg1202 = $signed(wire854);
              reg1203 <= ((reg1135[(3'h4):(3'h4)] ?
                      ((|(-reg1179)) ?
                          ((reg1194 ?
                              reg1173 : (7'h49)) < $signed(wire1090)) : reg1082[(4'h8):(3'h7)]) : $unsigned($unsigned($unsigned(reg1195)))) ?
                  {($signed($signed(wire853)) ?
                          (reg1108 ?
                              (reg1196 | (8'ha5)) : ((7'h42) ^ (8'hb9))) : reg1104[(5'h15):(3'h5)]),
                      (($unsigned(wire1091) ~^ $signed(reg1196)) * $unsigned(wire1091[(1'h0):(1'h0)]))} : reg1081);
              reg1204 = (($unsigned({(reg1194 * reg1114),
                          reg1132[(2'h2):(1'h1)]}) ?
                      $signed(reg1082[(4'h8):(4'h8)]) : $unsigned((~(reg1192 ?
                          (8'hab) : reg1085)))) ?
                  $signed({$unsigned($signed(reg1166))}) : $unsigned($signed(reg1194[(3'h5):(3'h5)])));
              reg1205 = ($unsigned($signed((8'hb5))) < $signed($unsigned((!(reg1183 + reg1203)))));
            end
          else
            begin
              reg1200 = (|$signed((($unsigned(wire1090) & reg1183) ?
                  $signed($unsigned(reg1118)) : wire853[(3'h6):(3'h5)])));
            end
          reg1206 = $signed($unsigned(($signed((reg1064 ?
              reg1099 : reg1205)) <= $signed(reg1166))));
          for (forvar1207 = (1'h0); (forvar1207 < (3'h4)); forvar1207 = (forvar1207 + (1'h1)))
            begin
              reg1208 = reg1204[(3'h5):(2'h3)];
              reg1209 <= reg1075;
              reg1210 = reg1163;
              reg1211 = {$signed($signed((^reg1061)))};
            end
          for (forvar1212 = (1'h0); (forvar1212 < (2'h2)); forvar1212 = (forvar1212 + (1'h1)))
            begin
              reg1213 <= ((~|(8'hb7)) ?
                  ($unsigned(reg1187) ^~ reg1195[(3'h7):(3'h5)]) : (^$signed(($signed(forvar1198) + (reg1204 >= reg1089)))));
              reg1214 = (~&$unsigned((reg1178 ?
                  $signed((^~wire1057)) : ($unsigned(reg1195) ?
                      reg1156[(2'h3):(2'h2)] : reg1156))));
              reg1215 = reg1172;
              reg1216 = $signed($unsigned((~|$unsigned((~|reg1196)))));
              reg1217 <= ((~|reg1104[(1'h0):(1'h0)]) <<< ((reg1067 ?
                  (reg1200[(1'h1):(1'h0)] ?
                      reg1081 : (|reg1183)) : reg1197) <= ($signed(reg1100) * ($signed(reg1216) ?
                  reg1188[(5'h11):(4'ha)] : $signed(reg1067)))));
            end
        end
    end
  module1218 #() modinst1291 (wire1290, clk, reg1173, reg1142, wire1091, reg1178, reg1179);
  always
    @(posedge clk) begin
      if ((8'haf))
        begin
          reg1292 = reg1109[(4'h8):(2'h2)];
          if ((-$unsigned((7'h4a))))
            begin
              reg1293 <= reg1217[(1'h0):(1'h0)];
            end
          else
            begin
              reg1294 = (($unsigned($signed((|wire1092))) ?
                  wire854[(1'h0):(1'h0)] : reg1099) - (~^(((wire854 ?
                          reg1199 : reg1078) ?
                      ((8'hbb) ? (8'hae) : reg1132) : $signed(reg1118)) ?
                  ((+(7'h41)) && reg1146[(4'hd):(2'h3)]) : wire1095[(3'h7):(1'h1)])));
              reg1295 <= (+($signed((8'hab)) * $unsigned((7'h44))));
              reg1296 = (((reg1163[(2'h3):(1'h0)] ^~ reg1294[(2'h2):(1'h1)]) & ((((7'h47) <= reg1148) <= (reg1168 ?
                      (8'had) : reg1099)) << $signed($signed(reg1186)))) ?
                  ($unsigned(reg1108[(5'h12):(4'he)]) | (((reg1168 ^ wire1057) ?
                      (reg1125 >> reg1176) : reg1186[(3'h4):(2'h3)]) ~^ $unsigned({reg1186,
                      reg1183}))) : (-$unsigned($unsigned(((8'h9f) ^ reg1203)))));
            end
        end
      else
        begin
          for (forvar1292 = (1'h0); (forvar1292 < (1'h0)); forvar1292 = (forvar1292 + (1'h1)))
            begin
              reg1293 <= reg1142;
            end
          if ((!($signed(($signed((8'h9e)) ?
              $signed(reg1065) : {wire856,
                  reg1135})) >> ($unsigned((reg1176 <= reg1176)) ?
              wire856 : (~&((8'hbd) <<< reg1295))))))
            begin
              reg1294 = ($unsigned($signed(wire1091[(3'h5):(1'h1)])) ?
                  reg1176 : (^~(((-reg1293) <= reg1294) == ((reg1065 ?
                      reg1099 : reg1176) != $signed(reg1108)))));
            end
          else
            begin
              reg1295 <= {reg1178,
                  ({{{(8'h9d), reg1109}},
                          $signed(((8'ha8) ? reg1209 : reg1295))} ?
                      reg1085 : (~^{(~|forvar1292)}))};
            end
        end
      for (forvar1297 = (1'h0); (forvar1297 < (2'h2)); forvar1297 = (forvar1297 + (1'h1)))
        begin
          reg1298 <= {(reg1110 < reg1172)};
          reg1299 <= $unsigned($unsigned(({(wire1093 >>> reg1213),
                  $unsigned(reg1176)} ?
              $signed(reg1135[(3'h7):(2'h3)]) : (+(reg1132 ?
                  reg1085 : (8'haf))))));
          reg1300 = $signed(wire853);
          reg1301 <= $signed($signed($signed($signed((8'hbd)))));
          reg1302 = (-(reg1110 != $signed(reg1109)));
        end
    end
  assign wire1303 = (^reg1187[(2'h2):(1'h1)]);
  always
    @(posedge clk) begin
      for (forvar1304 = (1'h0); (forvar1304 < (1'h1)); forvar1304 = (forvar1304 + (1'h1)))
        begin
          for (forvar1305 = (1'h0); (forvar1305 < (1'h1)); forvar1305 = (forvar1305 + (1'h1)))
            begin
              reg1306 <= reg1295;
              reg1307 = {wire1091, $unsigned($unsigned((8'h9f)))};
              reg1308 = reg1156[(2'h2):(2'h2)];
              reg1309 <= $signed(wire1094);
            end
          if (($signed((^$signed($signed((8'h9f))))) ?
              (((~^$signed(reg1081)) ?
                      (|wire1091) : ((~^reg1099) ?
                          ((8'hb1) ?
                              reg1118 : (8'haa)) : (reg1126 << reg1183))) ?
                  wire854 : wire1090) : $signed({reg1076[(4'hc):(1'h0)],
                  (~|(reg1071 ? reg1082 : reg1298))})))
            begin
              reg1310 = $signed((reg1065 - ((reg1203 <= $signed(reg1150)) ?
                  {(reg1112 <<< reg1209),
                      $signed(wire1057)} : $signed((reg1081 ?
                      wire1057 : reg1306)))));
              reg1311 <= reg1104[(4'he):(2'h2)];
              reg1312 = forvar1304[(3'h5):(2'h3)];
              reg1313 <= (((8'hb1) || (!reg1142)) ?
                  (reg1183 || reg1168) : (&(reg1311 != $signed((8'h9d)))));
            end
          else
            begin
              reg1311 <= ({forvar1305} ?
                  (^~$unsigned(reg1156[(2'h3):(2'h3)])) : ($signed($signed($signed(reg1118))) ?
                      reg1173[(5'h17):(4'h9)] : $unsigned({(|(8'hbc))})));
              reg1313 <= (|{(8'h9e)});
              reg1314 <= reg1075[(5'h17):(5'h17)];
            end
          reg1315 = $signed(reg1153);
          reg1316 = (~^reg1082);
        end
    end
  module1317 #() modinst1551 (wire1550, clk, wire856, wire1094, reg1199, reg1125);
  always
    @(posedge clk) begin
      reg1552 = $signed((^~$signed((~^reg1125))));
    end
  assign wire1553 = {(reg1100 ?
                            wire1550 : (reg1076[(4'hf):(3'h6)] ?
                                $signed($unsigned(reg1081)) : ($signed(reg1173) ?
                                    $signed(reg1061) : (~(8'hb6))))),
                        ($unsigned(($signed((8'ha5)) == {reg1078})) & reg1173[(4'h9):(3'h4)])};
  always
    @(posedge clk) begin
      reg1554 = $signed(({((wire1095 ?
              reg1129 : reg1108) <= (reg1217 > reg1166)),
          reg1213} < $signed($signed((reg1071 ? reg1309 : reg1309)))));
      reg1555 = (~&(reg1203[(3'h5):(1'h0)] < $signed(reg1166[(3'h7):(2'h2)])));
    end
  assign wire1556 = reg1187[(4'h9):(1'h1)];
  always
    @(posedge clk) begin
      if ((8'hb9))
        begin
          reg1557 <= (|reg1109[(1'h0):(1'h0)]);
        end
      else
        begin
          if ((($unsigned(($signed(wire1290) > $signed(reg1112))) * $signed((-$unsigned(reg1168)))) + reg1141))
            begin
              reg1558 = (((~^(reg1293[(2'h3):(2'h2)] ?
                          (wire1091 <<< reg1187) : reg1148[(4'hd):(4'hc)])) ?
                      reg1071[(4'h8):(2'h3)] : $unsigned($unsigned($signed(reg1082)))) ?
                  $signed(((!(wire1093 ? reg1076 : reg1076)) ?
                      (^$unsigned(reg1157)) : (reg1099[(1'h1):(1'h1)] | reg1116[(2'h3):(2'h2)]))) : reg1067);
              reg1559 <= $unsigned(wire854[(4'ha):(4'h8)]);
              reg1560 = $unsigned(($unsigned(($unsigned(reg1213) ?
                  reg1089 : {reg1109, reg1082})) >> wire1290[(4'h8):(1'h0)]));
            end
          else
            begin
              reg1558 = reg1203;
            end
          if (((((-(reg1193 ? reg1311 : reg1195)) ?
                      {$signed(reg1195)} : reg1065[(4'he):(4'hd)]) ?
                  $signed({$signed((8'ha8)), (&reg1089)}) : (~|$signed({wire856,
                      reg1067}))) ?
              reg1195 : (+(^reg1213))))
            begin
              reg1561 <= {({(~&(7'h44))} ?
                      reg1209[(3'h7):(2'h3)] : reg1195[(3'h7):(1'h0)])};
              reg1562 <= $unsigned({$unsigned(reg1153),
                  reg1201[(2'h3):(1'h1)]});
              reg1563 = reg1128;
              reg1564 <= reg1558;
            end
          else
            begin
              reg1563 = ($unsigned((8'hb1)) * $signed($signed((^~((8'ha5) <= (7'h40))))));
              reg1564 <= ((({$signed(reg1141)} ?
                      reg1195[(3'h6):(3'h5)] : wire1090[(2'h3):(1'h1)]) ?
                  $signed(reg1100[(3'h4):(1'h1)]) : $signed({reg1561})) && (^~$unsigned($unsigned({reg1201}))));
              reg1565 = reg1559;
              reg1566 <= ((+(reg1561 + {((8'ha4) ?
                      wire1290 : wire1550)})) ^ $unsigned(reg1157));
            end
          reg1567 <= ($signed($signed(((~&wire1556) && reg1168[(3'h6):(3'h6)]))) <= {$signed($unsigned(((8'hbb) != (8'h9f))))});
          reg1568 = reg1150[(3'h4):(3'h4)];
          reg1569 = (((reg1110[(5'h10):(4'hf)] ?
                  reg1141[(1'h1):(1'h0)] : $signed(reg1116[(2'h2):(2'h2)])) ?
              ($signed($unsigned(reg1560)) <= (|(wire1553 ?
                  reg1110 : wire1094))) : ($unsigned(((8'hbb) ~^ reg1089)) ?
                  (8'ha0) : reg1195[(2'h2):(1'h0)])) == (~|($signed((8'hac)) || $signed(reg1201))));
        end
      reg1570 <= ({reg1199} > $unsigned((~|$signed((!(8'ha5))))));
      reg1571 = $signed($unsigned($unsigned(((|reg1107) ?
          reg1186 : $signed(reg1109)))));
      reg1572 <= (reg1209 || reg1082);
      reg1573 <= (8'h9c);
    end
  always
    @(posedge clk) begin
      reg1574 = (7'h45);
      reg1575 = reg1193[(1'h0):(1'h0)];
      if ($signed(reg1195))
        begin
          for (forvar1576 = (1'h0); (forvar1576 < (1'h0)); forvar1576 = (forvar1576 + (1'h1)))
            begin
              reg1577 <= ($signed((~(8'hab))) ?
                  {(reg1176[(3'h5):(2'h3)] >> $signed({reg1089}))} : reg1061);
            end
          reg1578 <= (~&(|$signed(($unsigned(reg1301) << (reg1179 ?
              reg1574 : reg1577)))));
          if (({$signed((reg1128[(2'h3):(1'h1)] << reg1577)),
              ($unsigned(((8'ha0) ?
                  reg1559 : reg1173)) > wire1091)} << $unsigned((-((wire1290 > reg1168) ?
              (-reg1313) : wire1095[(3'h7):(2'h3)])))))
            begin
              reg1579 = (8'had);
            end
          else
            begin
              reg1579 = reg1298;
              reg1580 = {$unsigned((((8'hbb) ?
                      (~^wire1093) : (8'h9d)) >> $unsigned($unsigned(wire1303)))),
                  $unsigned(reg1199[(2'h2):(1'h0)])};
              reg1581 = (~|reg1183[(3'h6):(2'h2)]);
              reg1582 = $signed(forvar1576[(3'h6):(2'h3)]);
            end
          if ($unsigned(($signed((~^wire854[(4'hc):(2'h2)])) < reg1172[(4'h8):(1'h0)])))
            begin
              reg1583 = (~^(~^$signed({(|reg1582)})));
              reg1584 <= reg1570[(1'h0):(1'h0)];
              reg1585 = ($signed($signed({{reg1146}})) ?
                  wire1550 : reg1583[(2'h2):(1'h0)]);
            end
          else
            begin
              reg1583 = reg1579[(2'h2):(2'h2)];
              reg1585 = wire854[(4'h8):(4'h8)];
              reg1586 <= (reg1108[(3'h7):(1'h0)] ?
                  (+((8'hb5) >= reg1173)) : (8'hbf));
              reg1587 = reg1559;
            end
          if ($unsigned((~|((~$unsigned(reg1108)) ?
              reg1109 : (~&(reg1583 < reg1582))))))
            begin
              reg1588 = $signed($signed($unsigned($unsigned($unsigned(reg1581)))));
              reg1589 <= (&$unsigned({((reg1298 ?
                      reg1065 : wire1303) ^ reg1575[(1'h1):(1'h1)])}));
              reg1590 <= reg1564;
            end
          else
            begin
              reg1588 = reg1112;
              reg1589 <= (wire1057[(4'ha):(4'ha)] - reg1199[(5'h11):(4'h9)]);
              reg1590 <= reg1566[(3'h6):(1'h1)];
              reg1591 = $unsigned(reg1187[(1'h0):(1'h0)]);
              reg1592 <= reg1148;
            end
        end
      else
        begin
          if (((reg1178[(3'h6):(3'h6)] ?
                  wire855[(3'h4):(2'h2)] : $unsigned($signed((reg1067 ?
                      reg1141 : (8'haa))))) ?
              ($signed(((7'h43) ? $signed((8'hbc)) : $unsigned(reg1082))) ?
                  $signed($signed((-reg1301))) : {$signed($unsigned(wire1090)),
                      reg1309[(1'h1):(1'h1)]}) : $unsigned(reg1591[(1'h1):(1'h1)])))
            begin
              reg1576 <= wire1094[(3'h6):(3'h5)];
              reg1579 = $signed(wire1290[(4'hb):(1'h1)]);
              reg1584 <= reg1065[(5'h10):(4'he)];
            end
          else
            begin
              reg1576 <= reg1108[(3'h6):(1'h0)];
              reg1577 <= ((+reg1585[(4'hc):(1'h0)]) << wire1090[(4'h8):(3'h4)]);
            end
          for (forvar1585 = (1'h0); (forvar1585 < (1'h0)); forvar1585 = (forvar1585 + (1'h1)))
            begin
              reg1586 <= (-(|$unsigned(((8'ha0) & $signed(wire1290)))));
              reg1589 <= (reg1142 ?
                  reg1071[(4'h9):(2'h3)] : $signed($signed(forvar1576)));
              reg1590 <= reg1578;
            end
        end
    end
  assign wire1593 = (((~&reg1199[(5'h12):(1'h1)]) * reg1068) ?
                        (reg1142 ?
                            (|(~reg1301[(5'h12):(2'h3)])) : reg1173) : $signed(wire1091[(4'he):(4'hd)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module376
#(parameter param717 = (((8'ha9) ? (&(((8'hb0) ? (7'h42) : (8'hbe)) ? {(8'hb1), (8'hbe)} : ((8'hac) ? (8'hbd) : (8'hac)))) : (({(7'h40), (8'ha1)} * (!(8'ha1))) <= (~^(8'hb2)))) + (((!((8'hb2) ? (8'hba) : (8'hba))) ? ((~(7'h46)) << (+(8'hbf))) : (8'hb3)) == (((|(8'hbb)) <= (7'h45)) ? {((8'hae) ? (8'hb1) : (7'h44)), {(8'hab)}} : ((+(8'haa)) >>> ((8'hb8) ? (8'h9e) : (8'ha9)))))), 
parameter param718 = (param717 ? ((^~param717) ^ ((((8'h9c) ~^ param717) >> param717) ? param717 : (~|(param717 - param717)))) : (!{param717, (~|param717)})))
(y, clk, wire377, wire378, wire379, wire380, wire381);
  output wire [(32'h93a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h18):(1'h0)] wire377;
  input wire [(5'h16):(1'h0)] wire378;
  input wire [(5'h11):(1'h0)] wire379;
  input wire [(5'h11):(1'h0)] wire380;
  input wire signed [(4'hc):(1'h0)] wire381;
  wire [(4'hd):(1'h0)] wire686;
  wire signed [(4'hf):(1'h0)] wire665;
  wire signed [(5'h18):(1'h0)] wire635;
  wire signed [(2'h3):(1'h0)] wire634;
  wire [(2'h2):(1'h0)] wire630;
  wire signed [(5'h11):(1'h0)] wire382;
  wire [(5'h13):(1'h0)] wire512;
  wire [(5'h11):(1'h0)] wire544;
  wire signed [(5'h14):(1'h0)] wire584;
  reg [(5'h14):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg710 = (1'h0);
  reg [(4'he):(1'h0)] reg709 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg708 = (1'h0);
  reg [(3'h4):(1'h0)] reg707 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg706 = (1'h0);
  reg [(4'ha):(1'h0)] reg702 = (1'h0);
  reg [(5'h16):(1'h0)] reg699 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg695 = (1'h0);
  reg [(4'he):(1'h0)] reg693 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg691 = (1'h0);
  reg [(5'h15):(1'h0)] reg687 = (1'h0);
  reg [(4'hb):(1'h0)] reg685 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg684 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg683 = (1'h0);
  reg [(5'h14):(1'h0)] reg676 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg666 = (1'h0);
  reg [(5'h17):(1'h0)] reg675 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg674 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg672 = (1'h0);
  reg [(5'h17):(1'h0)] reg668 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg667 = (1'h0);
  reg [(4'h8):(1'h0)] reg664 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg662 = (1'h0);
  reg [(4'he):(1'h0)] reg660 = (1'h0);
  reg [(5'h14):(1'h0)] reg658 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg655 = (1'h0);
  reg [(4'h9):(1'h0)] reg651 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg650 = (1'h0);
  reg [(5'h13):(1'h0)] reg647 = (1'h0);
  reg [(4'hb):(1'h0)] reg646 = (1'h0);
  reg [(5'h13):(1'h0)] reg644 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg643 = (1'h0);
  reg [(3'h6):(1'h0)] reg642 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg636 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg633 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg632 = (1'h0);
  reg [(4'hc):(1'h0)] reg631 = (1'h0);
  reg [(3'h6):(1'h0)] reg623 = (1'h0);
  reg [(3'h7):(1'h0)] reg622 = (1'h0);
  reg [(2'h3):(1'h0)] reg621 = (1'h0);
  reg [(3'h5):(1'h0)] reg620 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg616 = (1'h0);
  reg [(4'hd):(1'h0)] reg615 = (1'h0);
  reg [(2'h2):(1'h0)] reg613 = (1'h0);
  reg [(5'h16):(1'h0)] reg611 = (1'h0);
  reg [(4'h8):(1'h0)] reg610 = (1'h0);
  reg [(2'h3):(1'h0)] reg605 = (1'h0);
  reg [(5'h14):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg586 = (1'h0);
  reg [(4'h9):(1'h0)] reg599 = (1'h0);
  reg [(4'hd):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg595 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg594 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg591 = (1'h0);
  reg signed [(4'he):(1'h0)] reg590 = (1'h0);
  reg [(4'hb):(1'h0)] reg588 = (1'h0);
  reg [(5'h14):(1'h0)] reg542 = (1'h0);
  reg [(5'h11):(1'h0)] reg539 = (1'h0);
  reg [(3'h5):(1'h0)] reg535 = (1'h0);
  reg [(4'hc):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg526 = (1'h0);
  reg [(5'h12):(1'h0)] reg523 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg518 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg520 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg714 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg713 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg712 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg711 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg705 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg704 = (1'h0);
  reg [(4'hb):(1'h0)] forvar703 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg701 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg700 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar698 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg697 = (1'h0);
  reg signed [(4'he):(1'h0)] reg696 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg694 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar692 = (1'h0);
  reg [(3'h7):(1'h0)] reg690 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar689 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg689 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg688 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar687 = (1'h0);
  reg [(5'h16):(1'h0)] reg682 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar681 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg680 = (1'h0);
  reg [(5'h11):(1'h0)] forvar679 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg678 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar677 = (1'h0);
  reg [(4'hf):(1'h0)] reg673 = (1'h0);
  reg [(5'h11):(1'h0)] reg671 = (1'h0);
  reg [(4'ha):(1'h0)] forvar670 = (1'h0);
  reg [(3'h7):(1'h0)] reg669 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar666 = (1'h0);
  reg [(5'h16):(1'h0)] reg663 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar659 = (1'h0);
  reg [(4'h8):(1'h0)] reg657 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg656 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg654 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg653 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg652 = (1'h0);
  reg [(5'h11):(1'h0)] reg649 = (1'h0);
  reg [(3'h4):(1'h0)] reg648 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg645 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar645 = (1'h0);
  reg [(5'h14):(1'h0)] reg641 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg640 = (1'h0);
  reg [(4'h9):(1'h0)] reg639 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg638 = (1'h0);
  reg [(4'h9):(1'h0)] reg637 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg629 = (1'h0);
  reg [(5'h16):(1'h0)] reg628 = (1'h0);
  reg [(3'h5):(1'h0)] reg627 = (1'h0);
  reg [(4'h9):(1'h0)] forvar626 = (1'h0);
  reg [(5'h15):(1'h0)] reg625 = (1'h0);
  reg [(5'h13):(1'h0)] forvar624 = (1'h0);
  reg [(4'hd):(1'h0)] reg619 = (1'h0);
  reg [(4'hd):(1'h0)] reg618 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg617 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg614 = (1'h0);
  reg [(3'h6):(1'h0)] reg612 = (1'h0);
  reg signed [(4'he):(1'h0)] reg609 = (1'h0);
  reg [(4'he):(1'h0)] forvar608 = (1'h0);
  reg [(5'h11):(1'h0)] reg607 = (1'h0);
  reg [(4'hc):(1'h0)] reg606 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar603 = (1'h0);
  reg [(5'h16):(1'h0)] forvar587 = (1'h0);
  reg [(4'h9):(1'h0)] reg602 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg601 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar600 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg598 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar597 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg593 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg592 = (1'h0);
  reg [(5'h17):(1'h0)] reg589 = (1'h0);
  reg [(5'h11):(1'h0)] reg587 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar586 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg543 = (1'h0);
  reg [(4'he):(1'h0)] reg541 = (1'h0);
  reg [(4'he):(1'h0)] reg540 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg538 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg537 = (1'h0);
  reg [(3'h4):(1'h0)] reg536 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar535 = (1'h0);
  reg [(5'h14):(1'h0)] reg534 = (1'h0);
  reg [(4'h8):(1'h0)] reg533 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg532 = (1'h0);
  reg [(5'h16):(1'h0)] forvar531 = (1'h0);
  reg [(4'hc):(1'h0)] forvar530 = (1'h0);
  reg [(4'hb):(1'h0)] reg529 = (1'h0);
  reg [(2'h3):(1'h0)] forvar527 = (1'h0);
  reg [(4'hc):(1'h0)] reg525 = (1'h0);
  reg [(4'hb):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg522 = (1'h0);
  reg [(4'hb):(1'h0)] reg521 = (1'h0);
  reg [(4'hb):(1'h0)] reg519 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar518 = (1'h0);
  reg [(4'ha):(1'h0)] reg517 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg516 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar514 = (1'h0);
  assign y = {wire686,
                 wire665,
                 wire635,
                 wire634,
                 wire630,
                 wire382,
                 wire512,
                 wire544,
                 wire584,
                 reg716,
                 reg715,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 reg702,
                 reg699,
                 reg695,
                 reg693,
                 reg691,
                 reg687,
                 reg685,
                 reg684,
                 reg683,
                 reg676,
                 reg666,
                 reg675,
                 reg674,
                 reg672,
                 reg668,
                 reg667,
                 reg664,
                 reg662,
                 reg660,
                 reg658,
                 reg655,
                 reg651,
                 reg650,
                 reg647,
                 reg646,
                 reg644,
                 reg643,
                 reg642,
                 reg636,
                 reg633,
                 reg632,
                 reg631,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 reg616,
                 reg615,
                 reg613,
                 reg611,
                 reg610,
                 reg605,
                 reg604,
                 reg586,
                 reg599,
                 reg596,
                 reg595,
                 reg594,
                 reg591,
                 reg590,
                 reg588,
                 reg542,
                 reg539,
                 reg535,
                 reg528,
                 reg526,
                 reg523,
                 reg518,
                 reg520,
                 reg714,
                 reg713,
                 reg712,
                 reg711,
                 reg705,
                 reg704,
                 forvar703,
                 reg701,
                 reg700,
                 forvar698,
                 reg697,
                 reg696,
                 reg694,
                 forvar692,
                 reg690,
                 forvar689,
                 reg689,
                 reg688,
                 forvar687,
                 reg682,
                 forvar681,
                 reg680,
                 forvar679,
                 reg678,
                 forvar677,
                 reg673,
                 reg671,
                 forvar670,
                 reg669,
                 forvar666,
                 reg663,
                 reg661,
                 forvar659,
                 reg657,
                 reg656,
                 reg654,
                 reg653,
                 reg652,
                 reg649,
                 reg648,
                 reg645,
                 forvar645,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg629,
                 reg628,
                 reg627,
                 forvar626,
                 reg625,
                 forvar624,
                 reg619,
                 reg618,
                 reg617,
                 reg614,
                 reg612,
                 reg609,
                 forvar608,
                 reg607,
                 reg606,
                 forvar603,
                 forvar587,
                 reg602,
                 reg601,
                 forvar600,
                 reg598,
                 forvar597,
                 reg593,
                 reg592,
                 reg589,
                 reg587,
                 forvar586,
                 reg543,
                 reg541,
                 reg540,
                 reg538,
                 reg537,
                 reg536,
                 forvar535,
                 reg534,
                 reg533,
                 reg532,
                 forvar531,
                 forvar530,
                 reg529,
                 forvar527,
                 reg525,
                 reg524,
                 reg522,
                 reg521,
                 reg519,
                 forvar518,
                 reg517,
                 reg516,
                 reg515,
                 forvar514,
                 (1'h0)};
  assign wire382 = ((($unsigned((wire380 ? (8'ha1) : wire381)) ?
                               $signed(wire378[(5'h15):(2'h2)]) : $signed((wire380 > wire380))) ?
                           $unsigned($signed((~wire379))) : $signed($unsigned(wire381[(4'h9):(3'h7)]))) ?
                       wire377 : {$signed((~&$signed(wire377))),
                           ((&(~&wire380)) && $unsigned((wire377 ?
                               wire380 : wire379)))});
  module383 #() modinst513 (wire512, clk, wire382, wire380, wire379, wire378);
  always
    @(posedge clk) begin
      if (wire378)
        begin
          for (forvar514 = (1'h0); (forvar514 < (2'h3)); forvar514 = (forvar514 + (1'h1)))
            begin
              reg515 = (!wire512[(1'h1):(1'h0)]);
              reg516 = (&$unsigned($signed(wire380[(4'h8):(2'h2)])));
              reg517 = reg515;
            end
          for (forvar518 = (1'h0); (forvar518 < (3'h4)); forvar518 = (forvar518 + (1'h1)))
            begin
              reg519 = (&$unsigned(((&(~wire382)) > $unsigned((forvar518 != reg516)))));
            end
          if ((|($signed((wire382[(4'hd):(4'ha)] < (|reg516))) && forvar514[(5'h16):(2'h3)])))
            begin
              reg520 <= ($signed((~^reg517[(4'ha):(2'h2)])) ?
                  (&$signed(((~|reg516) ^~ forvar514[(4'h9):(1'h1)]))) : reg517[(3'h4):(1'h1)]);
              reg521 = wire512;
              reg522 = (-($signed(wire512) ?
                  $unsigned(reg520[(2'h2):(1'h1)]) : $signed((~|(forvar518 & wire380)))));
            end
          else
            begin
              reg521 = (~^(!reg520[(4'hd):(4'h9)]));
              reg522 = reg515[(4'h9):(1'h1)];
            end
        end
      else
        begin
          for (forvar514 = (1'h0); (forvar514 < (2'h2)); forvar514 = (forvar514 + (1'h1)))
            begin
              reg518 <= $unsigned($unsigned(wire382[(2'h3):(1'h1)]));
              reg519 = $signed(wire380);
            end
          reg520 <= $signed(($signed($unsigned((!wire382))) ?
              (((wire379 ? wire382 : forvar518) ?
                  (8'ha8) : wire382[(4'hb):(3'h5)]) + wire379[(5'h11):(5'h10)]) : $unsigned($signed(wire380[(5'h11):(4'hf)]))));
          if ((+reg517[(2'h3):(1'h0)]))
            begin
              reg521 = forvar514;
              reg523 <= ((-{wire512,
                      (forvar518 == (wire377 ? forvar518 : (8'hac)))}) ?
                  $signed(wire381) : $unsigned($unsigned(forvar518[(1'h0):(1'h0)])));
              reg524 = (~|({(8'h9f), (~^$signed(wire381))} << (reg523 ?
                  $unsigned((wire378 ?
                      forvar514 : reg521)) : reg519[(4'h9):(1'h0)])));
              reg525 = (($unsigned(wire379) == wire379[(4'ha):(3'h5)]) <= ($signed({(^~reg523)}) ?
                  (^~((reg524 | wire381) >> (!wire379))) : ({(+wire380)} ?
                      $unsigned((reg516 ?
                          reg520 : wire382)) : reg524[(3'h6):(2'h3)])));
              reg526 <= ({$unsigned(((8'hab) ?
                      (reg519 ~^ (8'hbd)) : (^reg524))),
                  (^~reg522)} == wire377[(4'hd):(2'h3)]);
            end
          else
            begin
              reg523 <= (((&($signed(wire381) ?
                      (~^reg516) : wire378[(4'he):(3'h6)])) ?
                  forvar514 : wire382[(4'hb):(1'h1)]) ^ wire378);
              reg524 = forvar518;
              reg525 = (^~(!$unsigned((^~{wire379}))));
            end
        end
      for (forvar527 = (1'h0); (forvar527 < (2'h2)); forvar527 = (forvar527 + (1'h1)))
        begin
          reg528 <= reg521;
        end
      reg529 = $signed((reg528[(3'h5):(2'h2)] & wire380[(2'h2):(1'h1)]));
    end
  always
    @(posedge clk) begin
      for (forvar530 = (1'h0); (forvar530 < (1'h0)); forvar530 = (forvar530 + (1'h1)))
        begin
          for (forvar531 = (1'h0); (forvar531 < (3'h4)); forvar531 = (forvar531 + (1'h1)))
            begin
              reg532 = $signed($unsigned(wire381[(4'hb):(1'h0)]));
              reg533 = wire380[(5'h10):(3'h5)];
              reg534 = (~^reg520);
            end
        end
    end
  always
    @(posedge clk) begin
      if (($unsigned((+((wire512 ? wire378 : (8'hae)) ?
              (reg523 ? wire382 : (7'h47)) : (wire378 < reg528)))) ?
          $unsigned({{{wire512}}, $unsigned(wire512)}) : $signed({wire381,
              (wire382 != (~|wire381))})))
        begin
          for (forvar535 = (1'h0); (forvar535 < (2'h3)); forvar535 = (forvar535 + (1'h1)))
            begin
              reg536 = $unsigned({reg526,
                  ({(wire379 ? wire379 : reg518)} | $unsigned(((8'ha6) ?
                      reg520 : (8'hb1))))});
              reg537 = (wire379[(1'h0):(1'h0)] == wire378[(2'h2):(1'h1)]);
              reg538 = (wire512[(3'h7):(1'h0)] ~^ reg520);
            end
        end
      else
        begin
          if ($unsigned({(+wire377),
              $unsigned((reg518[(1'h1):(1'h0)] << $signed(forvar535)))}))
            begin
              reg535 <= reg528;
              reg536 = reg535;
              reg537 = {reg535[(2'h3):(2'h3)],
                  $signed($unsigned((^~$signed(reg536))))};
            end
          else
            begin
              reg536 = reg518;
              reg539 <= wire380[(4'h9):(3'h6)];
              reg540 = reg538[(2'h3):(2'h3)];
            end
          reg541 = (~&((8'hab) ?
              (!$unsigned(forvar535)) : reg537[(1'h1):(1'h0)]));
        end
      reg542 <= $unsigned($unsigned(reg523));
      reg543 = (({(reg528 ? reg526[(1'h1):(1'h0)] : reg523[(4'hf):(4'hb)]),
          $signed(wire379[(2'h2):(1'h1)])} & (reg528 <= (8'h9d))) + (~|wire377));
    end
  assign wire544 = {(8'h9c)};
  module545 #() modinst585 (.wire549(reg539), .wire550(reg542), .y(wire584), .wire546(reg518), .wire548(wire512), .clk(clk), .wire547(reg528));
  always
    @(posedge clk) begin
      if (wire382)
        begin
          for (forvar586 = (1'h0); (forvar586 < (3'h4)); forvar586 = (forvar586 + (1'h1)))
            begin
              reg587 = ($signed($unsigned((~&reg523[(4'he):(4'he)]))) == $signed($signed({$unsigned(wire512)})));
              reg588 <= ((wire380 >> $signed(wire584[(5'h13):(5'h13)])) + $unsigned($unsigned(($signed(wire584) ?
                  wire512 : reg526))));
              reg589 = wire380[(3'h5):(1'h0)];
            end
          if (wire378)
            begin
              reg590 <= (8'ha3);
              reg591 <= reg518[(1'h1):(1'h1)];
            end
          else
            begin
              reg592 = ((((^wire380) ?
                      (reg542[(2'h3):(2'h2)] ?
                          (wire382 >= reg528) : (reg528 & wire382)) : wire379) <<< $signed(($signed(reg535) ?
                      (wire512 ? reg542 : reg588) : {(8'hbc), (7'h41)}))) ?
                  $unsigned(wire379) : reg518);
              reg593 = (-reg592);
              reg594 <= reg592[(3'h7):(1'h1)];
              reg595 <= $unsigned((7'h42));
              reg596 <= forvar586;
            end
          for (forvar597 = (1'h0); (forvar597 < (2'h2)); forvar597 = (forvar597 + (1'h1)))
            begin
              reg598 = (-({(((8'ha0) ? reg542 : reg590) ?
                          $unsigned(reg591) : wire379)} ?
                  (({reg526,
                      reg539} && $unsigned(wire379)) + forvar597) : (8'ha6)));
            end
          reg599 <= $unsigned(($signed((~&(wire382 - reg595))) + $unsigned($signed(forvar597))));
          for (forvar600 = (1'h0); (forvar600 < (1'h0)); forvar600 = (forvar600 + (1'h1)))
            begin
              reg601 = (~&({wire378, $signed((reg526 ? reg535 : wire381))} ?
                  (!$signed($signed(forvar586))) : (($signed((8'hba)) | wire381[(1'h1):(1'h0)]) < $signed($unsigned(wire544)))));
              reg602 = ((reg591 && ($signed(((8'ha8) ? wire512 : reg588)) ?
                      ((~reg587) || $signed((8'haf))) : reg593[(5'h14):(3'h4)])) ?
                  {(({reg518} | {reg518, wire379}) ?
                          reg590 : reg528)} : ((reg588 ?
                          $unsigned($signed((8'hb7))) : reg590[(2'h2):(1'h1)]) ?
                      (~({wire584, wire382} ?
                          (wire377 <= wire378) : (reg595 * reg518))) : reg598));
            end
        end
      else
        begin
          reg586 <= (+$signed($signed({$unsigned(reg528),
              $unsigned(wire381)})));
          for (forvar587 = (1'h0); (forvar587 < (2'h3)); forvar587 = (forvar587 + (1'h1)))
            begin
              reg588 <= $unsigned((~|$signed(wire379[(4'hc):(2'h2)])));
              reg590 <= $signed(($unsigned({((7'h42) <= wire378),
                  (reg591 - reg528)}) ~^ $signed($signed((~&(8'hbc))))));
              reg591 <= (wire377[(5'h11):(1'h0)] ?
                  $signed((((reg598 >= wire381) >>> {(8'ha9)}) << (~&wire381))) : ($unsigned($unsigned($signed(wire544))) && (!(+(reg598 == forvar586)))));
            end
          reg592 = $unsigned(((($signed(wire512) ?
                  forvar597 : $unsigned(reg593)) ?
              ((-forvar597) > (reg520 ?
                  reg526 : reg594)) : $unsigned($signed(reg589))) == {$unsigned((reg526 & reg598)),
              $signed({wire380})}));
          reg593 = {{$unsigned({(-wire584), reg594})}, (~|(8'hbf))};
          reg594 <= reg594[(1'h1):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar603 = (1'h0); (forvar603 < (1'h0)); forvar603 = (forvar603 + (1'h1)))
        begin
          if (({((~&$signed(reg599)) ? $signed((^wire512)) : (~^(8'ha7))),
              reg596} | reg590[(4'ha):(3'h6)]))
            begin
              reg604 <= ((-{wire377,
                  ($signed(reg590) <<< {(7'h4a), reg586})}) << (|reg594));
              reg605 <= (^~$signed((-$unsigned(wire584[(4'hc):(2'h3)]))));
              reg606 = ((|$signed(($unsigned(wire512) ?
                      $unsigned(reg604) : {reg520, wire379}))) ?
                  $signed($unsigned(reg588)) : reg520);
              reg607 = wire378[(5'h12):(4'hb)];
            end
          else
            begin
              reg604 <= wire381[(1'h1):(1'h1)];
            end
        end
      if ($unsigned((-reg518)))
        begin
          for (forvar608 = (1'h0); (forvar608 < (2'h3)); forvar608 = (forvar608 + (1'h1)))
            begin
              reg609 = reg520;
              reg610 <= reg595;
              reg611 <= $unsigned($unsigned((&reg590[(3'h5):(1'h0)])));
              reg612 = (+(|reg526));
              reg613 <= (wire381[(4'ha):(3'h6)] ?
                  {(~(~&(reg604 ? forvar608 : reg611))),
                      $signed({(wire512 ^ wire584)})} : ((~^(&(reg594 ?
                          (7'h45) : forvar608))) ?
                      (&$signed(reg595)) : wire379[(4'hd):(2'h3)]));
            end
        end
      else
        begin
          for (forvar608 = (1'h0); (forvar608 < (1'h0)); forvar608 = (forvar608 + (1'h1)))
            begin
              reg610 <= $signed(wire379);
              reg612 = (8'hbb);
              reg614 = forvar608[(1'h0):(1'h0)];
              reg615 <= (((~|$unsigned((wire381 ?
                      reg606 : wire381))) != ($unsigned((reg518 ?
                      wire378 : reg591)) < $signed((-reg539)))) ?
                  (^~(reg604[(2'h3):(2'h2)] ?
                      (~|(wire379 <<< wire544)) : ($unsigned(wire544) >> (reg609 ?
                          reg523 : wire382)))) : ((-({forvar603,
                          reg523} && (reg520 ? reg595 : wire381))) ?
                      $unsigned($signed(reg591)) : (reg588 == (reg606[(1'h0):(1'h0)] != wire544[(4'h8):(2'h2)]))));
              reg616 <= $unsigned(reg614[(3'h4):(1'h0)]);
            end
          reg617 = ({reg605[(2'h2):(1'h0)]} || $signed(($unsigned((~&(8'hb7))) ?
              {(reg605 ? reg594 : reg518),
                  (wire377 ? (7'h44) : reg526)} : $signed({reg604, reg594}))));
          if ({(~&$signed({reg604[(5'h13):(4'hb)]})),
              (+$unsigned((((8'haa) ^~ reg591) | {(7'h46)})))})
            begin
              reg618 = $signed($unsigned((~&((wire512 ?
                  (8'hbc) : forvar608) & (reg590 > reg615)))));
              reg619 = {forvar603, reg618};
              reg620 <= wire377[(4'hd):(4'ha)];
            end
          else
            begin
              reg618 = ({$signed($unsigned({reg518})),
                      ((~&(reg607 ? reg612 : reg606)) ?
                          $unsigned((&wire381)) : (reg620[(2'h3):(2'h3)] ?
                              ((8'hb0) <<< reg586) : ((7'h46) ?
                                  reg539 : wire512)))} ?
                  ({reg588[(3'h5):(1'h0)],
                      reg518} > {$unsigned($unsigned(reg542)),
                      ((|reg590) && $unsigned((7'h44)))}) : ($signed(wire512[(2'h2):(1'h0)]) ?
                      reg617[(3'h6):(2'h2)] : $signed($signed((reg610 == reg595)))));
              reg620 <= ($signed((~&{(~reg595)})) * {$signed($signed((reg523 ?
                      reg595 : reg599))),
                  {($unsigned((8'h9c)) ?
                          (wire544 >>> (8'ha7)) : (reg595 || reg611)),
                      ($unsigned(wire381) ?
                          (wire378 > reg595) : ((8'hb4) >>> forvar608))}});
              reg621 <= ($signed($unsigned($signed((8'hbe)))) ?
                  (($unsigned((|reg590)) != $unsigned((+reg606))) <= ((~&(reg614 ?
                      reg619 : reg588)) & (reg616[(1'h0):(1'h0)] ^~ (reg614 ?
                      wire584 : (8'hae))))) : ((&$unsigned((+(8'hbb)))) ?
                      reg539[(5'h11):(4'hc)] : reg528[(4'h9):(1'h0)]));
              reg622 <= {{$unsigned(reg518[(1'h1):(1'h0)]),
                      reg539[(1'h1):(1'h0)]}};
              reg623 <= (-$unsigned($unsigned($unsigned(wire512))));
            end
        end
      for (forvar624 = (1'h0); (forvar624 < (1'h0)); forvar624 = (forvar624 + (1'h1)))
        begin
          reg625 = ((reg599 != reg586[(5'h12):(3'h5)]) ? reg617 : reg612);
          for (forvar626 = (1'h0); (forvar626 < (1'h1)); forvar626 = (forvar626 + (1'h1)))
            begin
              reg627 = ($signed((reg610[(2'h3):(2'h3)] ^ ({reg618} || reg523[(1'h0):(1'h0)]))) ?
                  reg542 : $unsigned(reg542));
              reg628 = $unsigned((^reg523));
            end
        end
      reg629 = $signed((&$unsigned(reg606)));
    end
  assign wire630 = $unsigned(reg586[(4'hf):(3'h5)]);
  always
    @(posedge clk) begin
      reg631 <= {($signed($signed($signed(wire380))) ?
              {$unsigned((wire381 ?
                      (8'h9d) : reg610))} : $signed({$unsigned(wire584),
                  reg623[(2'h3):(2'h2)]})),
          reg605[(1'h0):(1'h0)]};
      reg632 <= (!(-$unsigned(reg604)));
      reg633 <= ((reg620[(3'h4):(2'h2)] ?
          {wire381[(3'h4):(1'h0)]} : (((8'h9d) ?
              reg611[(5'h15):(4'hc)] : (reg631 >= reg542)) * (~&(-reg632)))) > $signed(reg610));
    end
  assign wire634 = reg599;
  assign wire635 = reg632[(4'h8):(4'h8)];
  always
    @(posedge clk) begin
      reg636 <= (~((~{$signed(reg631),
          $unsigned(reg611)}) || reg633[(4'h9):(4'h8)]));
      if ($signed($unsigned($signed(reg632[(4'h9):(3'h6)]))))
        begin
          reg637 = (!(|(~|(reg590 ?
              $signed((8'hae)) : (reg636 ? reg596 : reg599)))));
          reg638 = (reg520 ? wire635 : {reg539[(4'ha):(4'h8)]});
          if (($unsigned((8'h9e)) ?
              (($signed($unsigned(wire584)) ?
                      (|(wire380 ?
                          reg610 : (8'hae))) : $unsigned($signed(wire381))) ?
                  wire380[(4'hd):(3'h4)] : $signed((&{wire544}))) : $unsigned($unsigned($unsigned((reg637 ?
                  reg615 : (8'hb4)))))))
            begin
              reg639 = (&{$unsigned(((&reg632) ?
                      ((8'h9e) && reg604) : (reg518 ? wire584 : (8'hae)))),
                  {{(reg518 ^ reg621), $unsigned(reg542)}}});
              reg640 = (~|$unsigned($signed(reg613)));
              reg641 = $unsigned(((8'hb9) >> reg613));
            end
          else
            begin
              reg639 = {reg611,
                  {(($unsigned(reg595) ?
                          reg637 : wire512[(5'h12):(4'hd)]) * (^(8'h9d))),
                      wire544}};
              reg640 = (({wire380} ?
                      $unsigned(reg596[(4'h9):(1'h1)]) : $signed((wire377[(5'h10):(4'ha)] ?
                          reg633 : $signed(reg594)))) ?
                  reg599[(2'h2):(1'h1)] : $unsigned($signed(reg588)));
              reg642 <= reg539;
              reg643 <= {$signed($signed($signed((~&reg616)))),
                  (~|((8'ha7) && (!reg636[(2'h3):(1'h1)])))};
              reg644 <= reg604[(2'h3):(2'h3)];
            end
          for (forvar645 = (1'h0); (forvar645 < (2'h3)); forvar645 = (forvar645 + (1'h1)))
            begin
              reg646 <= $signed(reg644);
              reg647 <= $unsigned($unsigned({reg637[(3'h5):(3'h4)],
                  (reg523 == $signed(reg595))}));
            end
        end
      else
        begin
          if (((wire544[(5'h11):(4'hf)] ?
              reg639 : $unsigned({(~wire630)})) == $unsigned(reg639[(3'h7):(2'h3)])))
            begin
              reg642 <= reg644;
              reg643 <= {((~&$unsigned(reg520)) < reg599[(2'h3):(2'h2)]),
                  ((((~&(8'hb5)) ^~ {reg646}) ?
                      ((reg632 <= reg542) != {reg604}) : ((~|reg637) ?
                          reg611[(2'h2):(1'h0)] : (^~reg623))) * $unsigned({(~|(8'hb0)),
                      reg623[(3'h5):(2'h2)]}))};
              reg644 <= $signed($signed(reg632[(3'h5):(2'h2)]));
              reg645 = wire379;
              reg646 <= (reg645[(3'h6):(1'h1)] ^~ $signed((^$unsigned($unsigned(reg615)))));
            end
          else
            begin
              reg642 <= $signed($signed(wire635));
              reg645 = $unsigned($signed(((~$unsigned((8'hab))) == ((reg595 ?
                  reg611 : reg535) >>> (|reg616)))));
              reg648 = reg588[(4'h9):(1'h1)];
              reg649 = ($signed(reg599[(3'h6):(3'h4)]) ^~ (reg645[(5'h12):(2'h3)] < $unsigned(reg518)));
              reg650 <= (~&reg594);
            end
          if ($signed((|$unsigned(reg526))))
            begin
              reg651 <= reg649;
              reg652 = (~^{(((wire380 <<< (7'h47)) ?
                      (reg615 ?
                          reg613 : reg613) : reg520[(4'hb):(2'h2)]) > reg644),
                  ($unsigned((reg535 < reg594)) | $unsigned($unsigned(reg643)))});
              reg653 = (((~&$unsigned(reg638[(3'h7):(1'h1)])) >= reg636) >= $unsigned(reg599));
              reg654 = $signed($unsigned(reg648[(1'h1):(1'h0)]));
              reg655 <= $unsigned((~wire584[(5'h10):(4'h9)]));
            end
          else
            begin
              reg651 <= reg637[(3'h4):(2'h2)];
              reg655 <= $unsigned($signed(reg642[(3'h6):(1'h0)]));
              reg656 = $signed($signed(reg638));
              reg657 = (^~$signed((+reg542[(4'hc):(2'h2)])));
              reg658 <= {$signed($signed((reg611 + (-reg539))))};
            end
          for (forvar659 = (1'h0); (forvar659 < (3'h4)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 <= reg644[(4'hc):(1'h0)];
              reg661 = (wire382[(3'h5):(1'h1)] - $signed(reg595[(4'hd):(4'h8)]));
              reg662 <= (($unsigned((^(reg654 <= reg616))) == (^~(!(wire378 ?
                      reg586 : reg648)))) ?
                  {(7'h4a)} : (reg650[(1'h0):(1'h0)] >= $unsigned($unsigned((reg648 + wire381)))));
              reg663 = reg632[(1'h0):(1'h0)];
            end
          reg664 <= ((+$signed(((reg615 ? (8'hb0) : wire380) ^ (wire634 ?
                  reg621 : reg591)))) ?
              (reg623[(3'h4):(2'h2)] ?
                  {(reg613[(1'h0):(1'h0)] != $unsigned((7'h48))),
                      reg661[(3'h7):(1'h1)]} : $signed(reg542[(4'he):(1'h1)])) : reg616[(3'h5):(1'h1)]);
        end
    end
  assign wire665 = {$signed(((reg623[(2'h2):(1'h0)] ?
                               $signed(reg526) : {wire630, reg662}) ?
                           $signed($signed(reg664)) : (&$signed(reg643)))),
                       (^~((|reg535) * ((reg643 << wire634) - $signed(reg616))))};
  always
    @(posedge clk) begin
      if ($signed(wire379[(4'h8):(3'h6)]))
        begin
          for (forvar666 = (1'h0); (forvar666 < (1'h1)); forvar666 = (forvar666 + (1'h1)))
            begin
              reg667 <= (~&$signed($signed(((~reg622) & (8'hbd)))));
              reg668 <= reg605[(2'h3):(1'h0)];
            end
          reg669 = reg596;
          for (forvar670 = (1'h0); (forvar670 < (3'h4)); forvar670 = (forvar670 + (1'h1)))
            begin
              reg671 = ((~({reg662[(2'h2):(1'h0)]} ?
                  (-(reg590 ? (8'h9d) : (8'hb0))) : ({wire377} ?
                      $signed(wire381) : (8'hb7)))) <= wire379[(4'ha):(4'h9)]);
              reg672 <= ($unsigned($unsigned((+(reg664 ?
                  reg633 : reg671)))) ~^ reg588);
              reg673 = $signed(reg586);
              reg674 <= forvar666[(3'h5):(2'h3)];
            end
          reg675 <= $signed($unsigned((~|reg633[(4'hc):(3'h6)])));
        end
      else
        begin
          reg666 <= (^~reg621);
          reg669 = ($signed(reg644[(2'h3):(1'h0)]) ?
              (reg631 >>> ($signed(reg616) - reg647[(5'h12):(1'h1)])) : {{$signed((reg594 > reg613)),
                      (~$unsigned(reg636))}});
          for (forvar670 = (1'h0); (forvar670 < (3'h4)); forvar670 = (forvar670 + (1'h1)))
            begin
              reg671 = reg646;
            end
          reg672 <= reg523[(5'h11):(4'he)];
          reg674 <= reg616;
        end
      reg676 <= (~&((((reg520 == reg643) >>> (~&reg667)) >= $unsigned($signed(reg613))) ?
          $unsigned((8'hac)) : $unsigned((8'hac))));
      for (forvar677 = (1'h0); (forvar677 < (2'h2)); forvar677 = (forvar677 + (1'h1)))
        begin
          reg678 = wire381;
          for (forvar679 = (1'h0); (forvar679 < (1'h0)); forvar679 = (forvar679 + (1'h1)))
            begin
              reg680 = (-$unsigned(reg668));
            end
          for (forvar681 = (1'h0); (forvar681 < (1'h0)); forvar681 = (forvar681 + (1'h1)))
            begin
              reg682 = (reg591[(2'h3):(1'h1)] ?
                  {$unsigned($signed((reg660 ?
                          (8'hb2) : (8'hb7))))} : (~$unsigned({$unsigned(reg596)})));
              reg683 <= wire634[(2'h3):(1'h0)];
              reg684 <= $signed({$signed(((|reg671) ?
                      wire382 : (reg674 ? wire635 : wire635)))});
            end
        end
    end
  always
    @(posedge clk) begin
      reg685 <= $signed($signed(reg651));
    end
  assign wire686 = $signed(reg658[(5'h10):(5'h10)]);
  always
    @(posedge clk) begin
      if (wire382[(1'h0):(1'h0)])
        begin
          for (forvar687 = (1'h0); (forvar687 < (1'h1)); forvar687 = (forvar687 + (1'h1)))
            begin
              reg688 = wire635;
            end
          reg689 = (|$unsigned((reg666 == (~&((8'haf) << reg528)))));
        end
      else
        begin
          reg687 <= (~&reg613);
          reg688 = reg523;
          for (forvar689 = (1'h0); (forvar689 < (2'h3)); forvar689 = (forvar689 + (1'h1)))
            begin
              reg690 = $unsigned(((~&$unsigned($unsigned(reg664))) ?
                  $signed((~&(reg590 >>> reg644))) : $signed(((^~reg683) < ((8'ha4) <<< reg676)))));
              reg691 <= $unsigned(reg542);
            end
          for (forvar692 = (1'h0); (forvar692 < (1'h1)); forvar692 = (forvar692 + (1'h1)))
            begin
              reg693 <= (((((reg691 <<< reg662) ~^ (|reg539)) ?
                          $signed((~&wire380)) : {$signed(wire635)}) ?
                      reg658 : $unsigned((|(-reg675)))) ?
                  (((wire634 | (^wire382)) ?
                          wire377 : (~|forvar687[(5'h11):(2'h2)])) ?
                      reg616[(2'h2):(2'h2)] : $signed($signed(reg616[(2'h3):(1'h1)]))) : $signed($signed($unsigned($signed(reg687)))));
              reg694 = ($signed(reg674) != (forvar692[(3'h7):(1'h0)] ?
                  wire686[(4'h9):(1'h0)] : $unsigned((((8'haf) & reg690) ?
                      (8'hb8) : (-wire382)))));
              reg695 <= $signed(reg643[(2'h3):(1'h0)]);
              reg696 = ((~&$unsigned($unsigned(reg662[(4'h8):(1'h1)]))) >>> $unsigned((reg586[(4'he):(2'h3)] >>> (^$signed(wire635)))));
              reg697 = $unsigned({reg695, ($unsigned((&forvar689)) && reg613)});
            end
          for (forvar698 = (1'h0); (forvar698 < (3'h4)); forvar698 = (forvar698 + (1'h1)))
            begin
              reg699 <= ($signed((($signed(reg684) + $signed(reg685)) ?
                  wire665 : reg526)) << $unsigned((8'ha6)));
              reg700 = (reg636 <<< reg599[(3'h6):(1'h0)]);
              reg701 = $signed($unsigned($unsigned(reg611)));
              reg702 <= $unsigned((reg662 - $unsigned(reg535)));
            end
        end
      for (forvar703 = (1'h0); (forvar703 < (3'h4)); forvar703 = (forvar703 + (1'h1)))
        begin
          reg704 = {$unsigned((wire630 ? reg621 : (-(~reg662))))};
          if (($unsigned(wire380[(4'hc):(1'h0)]) & ((&$unsigned(reg590)) ^ $signed(reg700))))
            begin
              reg705 = wire379;
            end
          else
            begin
              reg705 = (($signed(reg586) ^ ($signed((wire635 ?
                      forvar689 : reg688)) > reg610[(4'h8):(1'h0)])) ?
                  $unsigned(wire512[(5'h13):(2'h2)]) : forvar689[(2'h2):(2'h2)]);
              reg706 <= (((~^(~&$signed(reg694))) + reg611[(4'ha):(3'h5)]) <= (!(|reg620)));
              reg707 <= (~forvar698);
            end
          reg708 <= reg672;
          if (reg704)
            begin
              reg709 <= (reg662[(2'h3):(2'h3)] | $unsigned({$unsigned($unsigned(reg588)),
                  reg664}));
              reg710 <= $unsigned($unsigned({reg685[(3'h6):(1'h1)],
                  ((&(8'hac)) <= $unsigned(wire382))}));
              reg711 = reg616[(1'h1):(1'h1)];
            end
          else
            begin
              reg711 = reg666;
              reg712 = $signed($unsigned((reg700[(3'h5):(1'h1)] ?
                  {$unsigned(reg646),
                      ((8'hb2) ? (8'ha9) : reg660)} : $signed((!reg632)))));
              reg713 = $unsigned((((reg706[(2'h2):(2'h2)] << $unsigned(reg604)) == ($unsigned(reg704) ?
                      reg613 : (wire380 ? reg586 : reg631))) ?
                  $unsigned($signed(reg528[(3'h7):(3'h4)])) : (($signed((8'h9d)) ?
                      reg610 : ((8'hbd) ?
                          reg675 : reg599)) <<< reg528[(2'h2):(2'h2)])));
              reg714 = wire379;
              reg715 <= reg642;
            end
          reg716 <= reg518;
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module545
#(parameter param582 = (~^{(((8'hac) ? (7'h47) : ((7'h40) ? (8'hb9) : (8'ha1))) ^~ {((7'h45) || (8'hb7)), ((8'hbf) > (8'ha5))})}), 
parameter param583 = (-{(~^(param582 << (param582 & param582))), {(!(+param582))}}))
(y, clk, wire550, wire549, wire548, wire547, wire546);
  output wire [(32'h1af):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire550;
  input wire [(5'h11):(1'h0)] wire549;
  input wire signed [(5'h13):(1'h0)] wire548;
  input wire [(4'hb):(1'h0)] wire547;
  input wire [(3'h5):(1'h0)] wire546;
  wire signed [(4'hc):(1'h0)] wire581;
  reg [(4'hc):(1'h0)] reg580 = (1'h0);
  reg [(5'h14):(1'h0)] reg579 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg577 = (1'h0);
  reg [(5'h10):(1'h0)] reg575 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg573 = (1'h0);
  reg [(3'h7):(1'h0)] reg572 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg569 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg567 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg566 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg560 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg559 = (1'h0);
  reg [(3'h7):(1'h0)] reg557 = (1'h0);
  reg [(4'hb):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg551 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg578 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar576 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg574 = (1'h0);
  reg [(5'h12):(1'h0)] reg571 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar568 = (1'h0);
  reg [(2'h3):(1'h0)] forvar561 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar556 = (1'h0);
  reg signed [(4'he):(1'h0)] reg565 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg563 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar562 = (1'h0);
  reg [(4'ha):(1'h0)] reg561 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg555 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg553 = (1'h0);
  reg [(3'h6):(1'h0)] reg552 = (1'h0);
  assign y = {wire581,
                 reg580,
                 reg579,
                 reg577,
                 reg575,
                 reg573,
                 reg572,
                 reg570,
                 reg569,
                 reg567,
                 reg566,
                 reg562,
                 reg564,
                 reg560,
                 reg559,
                 reg557,
                 reg556,
                 reg551,
                 reg578,
                 forvar576,
                 reg574,
                 reg571,
                 forvar568,
                 forvar561,
                 forvar556,
                 reg565,
                 reg563,
                 forvar562,
                 reg561,
                 reg558,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg551 <= wire550[(3'h7):(2'h2)];
      reg552 = $signed((~wire547[(4'ha):(4'ha)]));
      reg553 = reg552;
    end
  always
    @(posedge clk) begin
      reg554 = $signed($unsigned(wire550));
      if ((~|(({(^wire548), $unsigned(wire550)} - wire550) ?
          $unsigned($unsigned(wire549)) : (wire550 ?
              wire550[(3'h5):(3'h5)] : {wire547, (&wire550)}))))
        begin
          if ($unsigned($signed((((wire546 ? wire550 : wire547) ?
                  (wire549 ? wire549 : wire550) : wire547[(4'ha):(4'h9)]) ?
              ({reg554, reg551} << (wire546 ?
                  wire546 : wire548)) : wire550[(1'h0):(1'h0)]))))
            begin
              reg555 = $unsigned((&wire546));
            end
          else
            begin
              reg556 <= reg551[(2'h2):(1'h1)];
              reg557 <= $signed(wire549);
              reg558 = (($unsigned((|(~|wire549))) & wire548[(4'h8):(1'h1)]) & (~(&$unsigned(reg557))));
              reg559 <= $unsigned(reg555[(5'h12):(4'he)]);
              reg560 <= (reg551[(4'h9):(1'h1)] ?
                  ((~(reg559 > reg555[(4'ha):(3'h5)])) ?
                      {(~|reg556)} : reg554[(4'h8):(2'h3)]) : $signed((($unsigned(reg555) ?
                          wire546[(1'h1):(1'h1)] : $unsigned((8'ha9))) ?
                      $signed($unsigned(wire550)) : $signed((wire547 > wire550)))));
            end
          reg561 = {reg560};
          for (forvar562 = (1'h0); (forvar562 < (3'h4)); forvar562 = (forvar562 + (1'h1)))
            begin
              reg563 = (reg551[(4'h8):(2'h2)] & $signed($unsigned({((7'h44) ?
                      reg551 : reg551),
                  reg554})));
            end
          reg564 <= forvar562;
          reg565 = $unsigned(reg560);
        end
      else
        begin
          reg555 = reg559;
          for (forvar556 = (1'h0); (forvar556 < (2'h2)); forvar556 = (forvar556 + (1'h1)))
            begin
              reg557 <= ((8'hb4) ~^ ((~&reg558[(4'h8):(1'h0)]) & (8'haf)));
              reg559 <= ($signed((8'hbe)) >>> {$unsigned(wire548), (-reg561)});
            end
          reg560 <= (|($unsigned(($unsigned(reg558) ?
                  (wire546 ? (7'h4a) : forvar556) : $signed(reg565))) ?
              ($signed(wire549[(3'h5):(1'h0)]) ?
                  ((reg554 ? reg559 : reg561) ?
                      $unsigned(wire547) : reg561[(3'h7):(3'h5)]) : ((!reg556) ?
                      wire546[(1'h1):(1'h0)] : wire550)) : $unsigned(((~|wire550) << (reg555 ?
                  reg554 : wire550)))));
          for (forvar561 = (1'h0); (forvar561 < (2'h3)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 <= $unsigned($signed((8'hb9)));
              reg563 = ((forvar556[(2'h2):(1'h1)] ?
                      $signed(wire550[(1'h1):(1'h1)]) : $signed(((wire549 ?
                              wire547 : reg556) ?
                          ((8'ha2) << reg560) : wire548))) ?
                  (($signed(((8'hbc) + wire547)) ?
                      $unsigned({reg560}) : $signed((reg563 ^~ (8'hb6)))) & ($unsigned($signed(reg559)) - ($unsigned(reg555) ?
                      reg554[(3'h4):(3'h4)] : (!(8'hb5))))) : $unsigned((~{((7'h4a) ^~ reg560),
                      $unsigned(wire547)})));
              reg565 = $unsigned((reg555 * $unsigned((8'ha6))));
              reg566 <= (+$unsigned((reg557 ~^ reg554[(2'h3):(1'h0)])));
              reg567 <= reg559[(4'hc):(4'ha)];
            end
          for (forvar568 = (1'h0); (forvar568 < (3'h4)); forvar568 = (forvar568 + (1'h1)))
            begin
              reg569 <= forvar562;
              reg570 <= reg567[(3'h5):(2'h3)];
              reg571 = (^(reg567[(2'h2):(2'h2)] ?
                  $unsigned((forvar561[(1'h1):(1'h1)] ?
                      reg565 : (reg558 + reg567))) : (((forvar568 >>> reg566) ?
                      (~&forvar556) : (|forvar568)) == reg567)));
              reg572 <= reg569;
              reg573 <= $unsigned((|$unsigned(reg561[(2'h3):(1'h1)])));
            end
        end
      reg574 = $unsigned($unsigned(wire546[(3'h4):(1'h1)]));
      reg575 <= {wire548[(1'h1):(1'h0)]};
    end
  always
    @(posedge clk) begin
      for (forvar576 = (1'h0); (forvar576 < (1'h0)); forvar576 = (forvar576 + (1'h1)))
        begin
          if ((((^~wire550) << ($unsigned(reg575[(4'hc):(4'hc)]) ?
              (|(7'h47)) : {reg575[(3'h5):(2'h3)]})) >>> $unsigned(reg570)))
            begin
              reg577 <= (~^$signed($unsigned((^((8'hb7) ^~ reg560)))));
              reg578 = {wire549[(4'hd):(2'h2)], wire549[(2'h2):(2'h2)]};
              reg579 <= reg569;
              reg580 <= (|$signed(reg579[(3'h5):(3'h5)]));
            end
          else
            begin
              reg577 <= $unsigned($signed($signed($signed((reg566 << wire550)))));
              reg578 = reg560;
              reg579 <= $unsigned((reg579[(4'hb):(2'h2)] ^ reg570[(1'h1):(1'h0)]));
              reg580 <= reg559[(4'h9):(1'h0)];
            end
        end
    end
  assign wire581 = reg559;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module383  (y, clk, wire387, wire386, wire385, wire384);
  output wire [(32'h640):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire387;
  input wire [(5'h11):(1'h0)] wire386;
  input wire signed [(5'h11):(1'h0)] wire385;
  input wire signed [(5'h10):(1'h0)] wire384;
  wire [(4'he):(1'h0)] wire475;
  wire signed [(5'h14):(1'h0)] wire457;
  wire [(3'h4):(1'h0)] wire456;
  wire [(4'hb):(1'h0)] wire455;
  wire signed [(5'h14):(1'h0)] wire454;
  reg signed [(4'hf):(1'h0)] reg510 = (1'h0);
  reg [(5'h12):(1'h0)] reg509 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg508 = (1'h0);
  reg [(5'h12):(1'h0)] reg507 = (1'h0);
  reg [(3'h7):(1'h0)] reg501 = (1'h0);
  reg [(3'h5):(1'h0)] reg500 = (1'h0);
  reg [(5'h16):(1'h0)] reg498 = (1'h0);
  reg [(4'hd):(1'h0)] reg497 = (1'h0);
  reg [(3'h5):(1'h0)] reg495 = (1'h0);
  reg [(4'hb):(1'h0)] reg494 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg493 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg491 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg490 = (1'h0);
  reg [(5'h15):(1'h0)] reg488 = (1'h0);
  reg [(3'h6):(1'h0)] reg486 = (1'h0);
  reg [(4'h8):(1'h0)] reg485 = (1'h0);
  reg [(4'ha):(1'h0)] reg484 = (1'h0);
  reg [(4'hf):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg481 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg479 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg478 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg469 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg468 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg465 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg464 = (1'h0);
  reg [(5'h12):(1'h0)] reg463 = (1'h0);
  reg [(4'h8):(1'h0)] reg460 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg458 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg453 = (1'h0);
  reg [(2'h2):(1'h0)] reg451 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg450 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg446 = (1'h0);
  reg [(4'hb):(1'h0)] reg445 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg441 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg437 = (1'h0);
  reg [(4'h9):(1'h0)] reg436 = (1'h0);
  reg [(3'h5):(1'h0)] reg435 = (1'h0);
  reg [(2'h3):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg431 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg430 = (1'h0);
  reg [(5'h15):(1'h0)] reg427 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg426 = (1'h0);
  reg [(4'hf):(1'h0)] reg424 = (1'h0);
  reg [(5'h17):(1'h0)] reg423 = (1'h0);
  reg [(4'h8):(1'h0)] reg422 = (1'h0);
  reg [(5'h17):(1'h0)] reg418 = (1'h0);
  reg [(2'h3):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg414 = (1'h0);
  reg [(4'hd):(1'h0)] reg413 = (1'h0);
  reg [(2'h2):(1'h0)] reg409 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg408 = (1'h0);
  reg [(5'h10):(1'h0)] reg405 = (1'h0);
  reg [(4'ha):(1'h0)] reg404 = (1'h0);
  reg [(5'h11):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg394 = (1'h0);
  reg [(2'h2):(1'h0)] reg392 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg511 = (1'h0);
  reg [(3'h5):(1'h0)] forvar510 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg506 = (1'h0);
  reg [(5'h12):(1'h0)] reg505 = (1'h0);
  reg [(5'h14):(1'h0)] forvar504 = (1'h0);
  reg [(5'h14):(1'h0)] reg503 = (1'h0);
  reg [(4'h9):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg502 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar499 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg496 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg492 = (1'h0);
  reg [(4'he):(1'h0)] forvar489 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg483 = (1'h0);
  reg [(3'h6):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar477 = (1'h0);
  reg [(5'h16):(1'h0)] forvar476 = (1'h0);
  reg [(3'h4):(1'h0)] reg474 = (1'h0);
  reg signed [(4'he):(1'h0)] reg473 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg471 = (1'h0);
  reg [(5'h15):(1'h0)] reg470 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg467 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg466 = (1'h0);
  reg [(3'h4):(1'h0)] forvar462 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg461 = (1'h0);
  reg [(3'h6):(1'h0)] reg447 = (1'h0);
  reg [(5'h10):(1'h0)] forvar452 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg448 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar447 = (1'h0);
  reg [(5'h14):(1'h0)] forvar444 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar443 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg442 = (1'h0);
  reg [(4'hd):(1'h0)] reg440 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg439 = (1'h0);
  reg [(2'h3):(1'h0)] reg438 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg434 = (1'h0);
  reg [(2'h3):(1'h0)] reg432 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg429 = (1'h0);
  reg [(3'h5):(1'h0)] forvar428 = (1'h0);
  reg [(4'hc):(1'h0)] reg425 = (1'h0);
  reg [(4'hc):(1'h0)] forvar421 = (1'h0);
  reg [(4'ha):(1'h0)] forvar409 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg420 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg419 = (1'h0);
  reg signed [(4'he):(1'h0)] reg417 = (1'h0);
  reg [(4'hd):(1'h0)] reg415 = (1'h0);
  reg [(5'h18):(1'h0)] reg412 = (1'h0);
  reg [(4'h8):(1'h0)] reg411 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg410 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg406 = (1'h0);
  reg [(4'h8):(1'h0)] reg402 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg401 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar397 = (1'h0);
  reg [(5'h18):(1'h0)] reg396 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar395 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg393 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg391 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg390 = (1'h0);
  reg [(5'h16):(1'h0)] forvar389 = (1'h0);
  reg [(3'h4):(1'h0)] forvar388 = (1'h0);
  assign y = {wire475,
                 wire457,
                 wire456,
                 wire455,
                 wire454,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg501,
                 reg500,
                 reg498,
                 reg497,
                 reg495,
                 reg494,
                 reg493,
                 reg491,
                 reg490,
                 reg488,
                 reg486,
                 reg485,
                 reg484,
                 reg482,
                 reg481,
                 reg479,
                 reg478,
                 reg472,
                 reg469,
                 reg468,
                 reg465,
                 reg464,
                 reg463,
                 reg460,
                 reg459,
                 reg458,
                 reg453,
                 reg451,
                 reg450,
                 reg449,
                 reg446,
                 reg445,
                 reg441,
                 reg437,
                 reg436,
                 reg435,
                 reg433,
                 reg431,
                 reg430,
                 reg427,
                 reg426,
                 reg424,
                 reg423,
                 reg422,
                 reg418,
                 reg416,
                 reg414,
                 reg413,
                 reg409,
                 reg408,
                 reg405,
                 reg404,
                 reg403,
                 reg400,
                 reg398,
                 reg394,
                 reg392,
                 reg511,
                 forvar510,
                 reg506,
                 reg505,
                 forvar504,
                 reg503,
                 reg499,
                 reg502,
                 forvar499,
                 reg496,
                 reg492,
                 forvar489,
                 reg487,
                 reg483,
                 reg480,
                 forvar477,
                 forvar476,
                 reg474,
                 reg473,
                 reg471,
                 reg470,
                 reg467,
                 reg466,
                 forvar462,
                 reg461,
                 reg447,
                 forvar452,
                 reg448,
                 forvar447,
                 forvar444,
                 forvar443,
                 reg442,
                 reg440,
                 reg439,
                 reg438,
                 reg434,
                 reg432,
                 reg429,
                 forvar428,
                 reg425,
                 forvar421,
                 forvar409,
                 reg420,
                 reg419,
                 reg417,
                 reg415,
                 reg412,
                 reg411,
                 reg410,
                 reg407,
                 reg406,
                 reg402,
                 reg401,
                 reg399,
                 forvar397,
                 reg396,
                 forvar395,
                 reg393,
                 reg391,
                 reg390,
                 forvar389,
                 forvar388,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar388 = (1'h0); (forvar388 < (2'h3)); forvar388 = (forvar388 + (1'h1)))
        begin
          for (forvar389 = (1'h0); (forvar389 < (1'h0)); forvar389 = (forvar389 + (1'h1)))
            begin
              reg390 = {($unsigned($signed(wire387[(4'he):(4'hc)])) ?
                      (wire387[(4'hd):(4'hc)] == ($signed(forvar388) ?
                          wire387 : $unsigned(forvar389))) : wire384)};
              reg391 = (&$unsigned(((((8'hb3) ? (8'had) : wire386) ?
                  $unsigned(forvar388) : (wire384 ?
                      forvar388 : (8'h9c))) == $unsigned((~&wire384)))));
              reg392 <= $signed(wire386);
            end
          reg393 = $unsigned(reg392[(2'h2):(1'h1)]);
          reg394 <= $unsigned((8'ha8));
        end
      for (forvar395 = (1'h0); (forvar395 < (1'h1)); forvar395 = (forvar395 + (1'h1)))
        begin
          reg396 = $signed(($signed((~(forvar389 * reg393))) << (reg391 ?
              ($unsigned(reg391) || (forvar388 << wire384)) : reg391[(3'h4):(2'h2)])));
          for (forvar397 = (1'h0); (forvar397 < (3'h4)); forvar397 = (forvar397 + (1'h1)))
            begin
              reg398 <= (~^wire387);
              reg399 = (|$signed((~|(^~(&forvar389)))));
              reg400 <= (7'h44);
              reg401 = (reg398 ? reg392 : {reg392[(1'h1):(1'h0)]});
              reg402 = $signed(($signed(((~forvar395) ?
                  reg401 : $signed(wire385))) >= (-($unsigned(reg401) < reg390))));
            end
          reg403 <= ((^~$signed(forvar395)) | (reg402 ?
              (($signed(reg390) ^~ wire386[(3'h5):(3'h4)]) + wire386) : $signed({$signed((8'ha3)),
                  $signed(reg390)})));
        end
      if (($unsigned($signed($unsigned($unsigned(reg402)))) - ((~|$signed(reg393[(4'h9):(1'h1)])) ~^ $signed({$unsigned(reg399)}))))
        begin
          if ($signed({($unsigned((~^wire387)) ?
                  $signed((+reg400)) : $unsigned((wire385 == forvar388))),
              {(^~(reg402 | reg393))}}))
            begin
              reg404 <= ($unsigned(wire387) | $signed(($unsigned((+reg393)) ?
                  {{reg396}} : reg400[(4'he):(4'hd)])));
              reg405 <= reg390[(3'h5):(2'h3)];
            end
          else
            begin
              reg404 <= $signed($unsigned(reg405));
              reg406 = (!$signed((^~forvar388)));
              reg407 = reg394[(4'hb):(3'h4)];
              reg408 <= ($unsigned($unsigned(((forvar389 <<< (8'hac)) - (reg401 + reg391)))) ?
                  reg406 : (((-{reg406, wire387}) ?
                          (reg391[(4'h9):(3'h5)] ?
                              reg390[(4'h8):(1'h0)] : {reg393,
                                  reg407}) : ((!wire384) & (forvar397 ?
                              forvar389 : reg398))) ?
                      reg392[(1'h1):(1'h1)] : (-reg391[(1'h0):(1'h0)])));
            end
          if (((7'h48) << $signed((~reg391[(1'h1):(1'h0)]))))
            begin
              reg409 <= {{(($unsigned(forvar388) ?
                              (reg404 ?
                                  reg404 : forvar395) : (reg404 ~^ reg404)) ?
                          $signed($signed((8'hb8))) : wire384),
                      (+$signed((7'h47)))},
                  (+{(~|(~^reg403)), $signed(forvar397)})};
            end
          else
            begin
              reg410 = $signed({$unsigned(reg391),
                  $signed($signed($unsigned(reg392)))});
            end
          reg411 = reg394;
          reg412 = reg394;
          if (((+reg401[(2'h2):(1'h1)]) <<< (8'hb5)))
            begin
              reg413 <= {$signed($unsigned(forvar389)),
                  {reg401,
                      ((^~$signed(reg402)) ?
                          ((reg392 ?
                              reg409 : reg394) | reg411[(3'h7):(2'h3)]) : $signed(wire387[(2'h2):(1'h1)]))}};
              reg414 <= $signed($unsigned($signed(((forvar395 ?
                      reg413 : reg413) ?
                  (reg413 ? reg405 : (8'hbc)) : (reg403 ^~ reg398)))));
              reg415 = ($signed((forvar395[(1'h1):(1'h0)] >>> forvar389)) == (reg407[(4'ha):(1'h0)] ?
                  forvar397[(2'h2):(1'h1)] : $signed(forvar397[(1'h0):(1'h0)])));
              reg416 <= wire385[(3'h7):(3'h4)];
            end
          else
            begin
              reg415 = (reg408 < reg413[(4'hd):(2'h3)]);
              reg417 = $signed((+$signed((reg390 ?
                  (~&reg407) : (reg413 ? reg390 : reg411)))));
              reg418 <= ($signed(((|reg392) >>> $unsigned($unsigned(reg402)))) & $signed((($unsigned(reg407) ?
                  reg415[(4'h9):(3'h5)] : (^~reg409)) == reg396[(4'ha):(4'h8)])));
              reg419 = (((reg415 ?
                      $signed($signed(reg405)) : (reg410[(4'h9):(1'h1)] ?
                          reg400[(3'h4):(2'h2)] : reg403[(5'h11):(4'hf)])) <<< $unsigned(forvar388)) ?
                  (~&forvar389[(1'h1):(1'h1)]) : (8'ha6));
              reg420 = $unsigned($unsigned($unsigned(((reg416 || wire387) ?
                  reg412 : $signed(reg407)))));
            end
        end
      else
        begin
          reg404 <= (($signed((&(reg390 & (7'h49)))) ?
                  reg407 : ($signed(reg392) ~^ reg409)) ?
              (reg401 ?
                  $unsigned($unsigned(reg410[(3'h6):(2'h2)])) : (^((~&wire387) ?
                      (reg418 && reg409) : reg405))) : (reg411[(4'h8):(3'h4)] ?
                  wire385 : ($signed((reg404 << reg402)) << (reg412[(3'h6):(3'h4)] ?
                      forvar395[(2'h2):(1'h0)] : (~|reg413)))));
          reg405 <= (($unsigned({reg401,
                  $unsigned(reg392)}) <= $unsigned(((&reg412) ?
                  (-reg391) : (8'hb5)))) ?
              (-$unsigned({reg408[(1'h0):(1'h0)],
                  (~|reg398)})) : $signed((+$unsigned((reg404 ?
                  wire387 : forvar389)))));
          reg408 <= (!((-$unsigned((~|reg390))) ?
              ($signed($unsigned(reg409)) == wire385[(4'h9):(4'h9)]) : (reg410 << $unsigned(wire386[(2'h3):(2'h3)]))));
          for (forvar409 = (1'h0); (forvar409 < (2'h2)); forvar409 = (forvar409 + (1'h1)))
            begin
              reg410 = reg399;
              reg413 <= $unsigned({(8'ha1),
                  $signed($signed(reg409[(2'h2):(1'h1)]))});
              reg414 <= (|(8'hb4));
            end
        end
      for (forvar421 = (1'h0); (forvar421 < (1'h0)); forvar421 = (forvar421 + (1'h1)))
        begin
          reg422 <= (($signed(({reg408} ?
                  (reg390 & reg409) : (reg414 ? reg393 : reg401))) ?
              reg394 : $unsigned((~reg391))) ^ ((wire385[(4'he):(2'h3)] ?
              $unsigned((reg413 ?
                  reg419 : forvar397)) : reg400[(4'ha):(3'h6)]) | forvar397));
          reg423 <= wire387[(2'h3):(1'h1)];
          reg424 <= (|(^(^~(&reg403))));
          reg425 = reg407[(2'h3):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      reg426 <= (reg403 < (&(^reg403[(5'h11):(3'h7)])));
      reg427 <= reg403;
    end
  always
    @(posedge clk) begin
      for (forvar428 = (1'h0); (forvar428 < (1'h1)); forvar428 = (forvar428 + (1'h1)))
        begin
          reg429 = (reg418 ?
              $unsigned($signed($signed((reg400 ?
                  reg392 : reg427)))) : (^~$unsigned($signed((|reg392)))));
          if (reg429[(1'h0):(1'h0)])
            begin
              reg430 <= reg422;
              reg431 <= reg414[(3'h5):(1'h1)];
              reg432 = (~^reg416);
              reg433 <= ((~|reg422) ?
                  {(reg400[(3'h5):(3'h4)] + ((~&wire386) ?
                          (reg422 | reg424) : (reg403 ?
                              (8'ha2) : (7'h41))))} : reg408);
              reg434 = ($unsigned((8'ha7)) ?
                  $signed($unsigned($unsigned({reg424}))) : ((wire385 || ($signed((8'ha8)) ?
                          $unsigned(reg414) : reg404)) ?
                      $unsigned($signed(forvar428[(2'h2):(2'h2)])) : ($unsigned((wire387 ?
                          reg403 : reg422)) && $unsigned((!wire387)))));
            end
          else
            begin
              reg430 <= $unsigned((+(reg422 ^ (^~reg416))));
              reg431 <= (8'hbc);
              reg433 <= ($signed($signed(reg400)) ?
                  reg427 : (reg432 ?
                      $signed($unsigned(reg400[(5'h13):(4'h8)])) : $signed((^~reg431[(3'h5):(2'h3)]))));
              reg435 <= ((wire384 ?
                  reg429[(1'h1):(1'h0)] : reg431) >>> ((+$unsigned(((8'ha0) + reg404))) ?
                  $unsigned((^reg403[(5'h11):(3'h4)])) : (wire387 <= (8'h9f))));
            end
          if ((((~&(wire384[(2'h2):(2'h2)] >> {reg424})) ?
              {(^~(reg409 ?
                      reg400 : wire386))} : reg429) << $signed($unsigned($unsigned(wire387[(1'h0):(1'h0)])))))
            begin
              reg436 <= $signed($unsigned(((reg418[(2'h3):(1'h0)] ?
                      reg403[(4'h9):(1'h0)] : $signed(reg430)) ?
                  (^reg400[(4'he):(1'h1)]) : reg416)));
              reg437 <= $signed(reg408);
            end
          else
            begin
              reg438 = reg413[(1'h1):(1'h1)];
              reg439 = reg424[(4'hd):(4'hb)];
              reg440 = ($unsigned((8'h9c)) >>> reg404[(4'h9):(4'h9)]);
            end
          reg441 <= (~|(|reg394));
          reg442 = $signed(reg439);
        end
      for (forvar443 = (1'h0); (forvar443 < (1'h0)); forvar443 = (forvar443 + (1'h1)))
        begin
          for (forvar444 = (1'h0); (forvar444 < (2'h2)); forvar444 = (forvar444 + (1'h1)))
            begin
              reg445 <= $signed($signed(({{reg430, reg416},
                      $signed(forvar428)} ?
                  reg429 : ((reg430 ? reg439 : reg432) ?
                      $unsigned(reg416) : $signed((7'h42))))));
            end
          reg446 <= $signed(forvar444);
        end
      if (($signed($unsigned($signed($unsigned(reg445)))) ?
          ($unsigned($signed((+reg435))) ^~ reg434) : $signed(reg422)))
        begin
          for (forvar447 = (1'h0); (forvar447 < (1'h0)); forvar447 = (forvar447 + (1'h1)))
            begin
              reg448 = reg430;
              reg449 <= reg445[(4'hb):(3'h6)];
            end
          reg450 <= ((forvar444 ?
              {{$unsigned(reg416)}} : (~^(forvar444[(5'h13):(1'h1)] * $signed(forvar443)))) >>> $signed($unsigned((^~(reg436 != (8'hab))))));
          reg451 <= ((|(($unsigned((8'hbd)) + $signed(reg439)) != $unsigned($signed(reg430)))) > forvar447[(3'h4):(3'h4)]);
          for (forvar452 = (1'h0); (forvar452 < (1'h1)); forvar452 = (forvar452 + (1'h1)))
            begin
              reg453 <= $unsigned((reg435[(2'h2):(2'h2)] ^~ (8'hb3)));
            end
        end
      else
        begin
          reg447 = ($unsigned((-$signed(reg450))) >= reg433[(2'h3):(2'h2)]);
          reg449 <= reg442;
        end
    end
  assign wire454 = (($signed({reg405}) ? reg422[(3'h7):(1'h0)] : (&(+reg418))) ?
                       $signed(reg422) : wire385[(1'h0):(1'h0)]);
  assign wire455 = (reg453[(3'h5):(1'h0)] ?
                       $signed((^~((reg409 ? reg450 : reg405) ?
                           $unsigned(wire387) : reg426[(4'ha):(4'h8)]))) : $unsigned((^((~^(8'hb9)) ?
                           (~^(8'hb8)) : wire454))));
  assign wire456 = $unsigned((!reg445));
  assign wire457 = {(($signed(reg422) | wire455) == wire385), reg408};
  always
    @(posedge clk) begin
      reg458 <= (|reg409);
      reg459 <= (!$unsigned((!(^~reg446))));
      if (reg398[(3'h7):(3'h6)])
        begin
          reg460 <= (((8'ha9) != reg414) >= (~&reg453));
          reg461 = $unsigned($unsigned((|$unsigned($signed((8'ha4))))));
        end
      else
        begin
          reg461 = {$signed($unsigned((~&reg416[(1'h0):(1'h0)]))),
              ({{reg431}, ((&reg459) ? (reg426 < reg398) : (8'hb8))} ?
                  wire455[(2'h2):(1'h1)] : ((reg405[(2'h3):(1'h0)] ?
                      (reg423 ?
                          reg414 : reg437) : $signed(wire386)) ^~ ($signed(reg446) ?
                      $unsigned(reg392) : ((8'hbe) ? reg403 : reg418))))};
        end
      for (forvar462 = (1'h0); (forvar462 < (1'h1)); forvar462 = (forvar462 + (1'h1)))
        begin
          if ((|(-($unsigned(reg409) ? {reg460[(2'h3):(1'h0)]} : (8'hbf)))))
            begin
              reg463 <= ($signed($signed(($unsigned(reg460) && reg446[(4'h8):(4'h8)]))) ^~ wire457[(4'he):(3'h5)]);
              reg464 <= wire385;
              reg465 <= (8'hb8);
              reg466 = {(reg450[(2'h3):(1'h1)] * $unsigned(((~reg414) <<< (reg463 <= reg446))))};
              reg467 = reg460[(2'h2):(1'h0)];
            end
          else
            begin
              reg466 = (~$signed((~^$signed((reg423 ? wire456 : reg446)))));
            end
          reg468 <= (wire454[(5'h14):(5'h12)] << $signed((((reg459 ?
                  reg413 : reg446) >= $unsigned(reg445)) ?
              $signed($unsigned(reg446)) : reg422[(3'h4):(3'h4)])));
          if ($unsigned(({reg459, reg465[(2'h3):(2'h2)]} ?
              (reg465 >> ((8'hae) ?
                  $signed(reg404) : reg416[(2'h2):(1'h0)])) : (~&$unsigned($signed(wire456))))))
            begin
              reg469 <= ({$signed(((reg427 < reg392) || (wire455 ?
                          wire384 : reg404))),
                      reg427} ?
                  (~^reg446) : reg405[(4'hc):(1'h1)]);
              reg470 = reg403;
              reg471 = (($unsigned(((|reg453) ?
                  (reg435 && wire386) : reg446)) != {$signed($unsigned(reg468)),
                  (+$signed(reg451))}) >= $signed({reg445,
                  $signed($signed(reg416))}));
            end
          else
            begin
              reg469 <= (8'h9e);
              reg472 <= reg408;
              reg473 = (-$signed(reg403[(2'h2):(1'h1)]));
            end
        end
      reg474 = (reg459 && ($signed(reg403) != $signed(({wire454, (8'hb1)} ?
          (!(7'h41)) : reg449))));
    end
  assign wire475 = (^~(|reg460[(2'h2):(1'h1)]));
  always
    @(posedge clk) begin
      for (forvar476 = (1'h0); (forvar476 < (2'h3)); forvar476 = (forvar476 + (1'h1)))
        begin
          for (forvar477 = (1'h0); (forvar477 < (2'h2)); forvar477 = (forvar477 + (1'h1)))
            begin
              reg478 <= (-reg398[(4'hd):(3'h5)]);
              reg479 <= ({reg418[(5'h12):(5'h10)],
                  (~reg427[(1'h1):(1'h0)])} | {(((|wire384) ?
                          reg459[(2'h2):(1'h1)] : (reg433 == (8'ha8))) ?
                      $signed($unsigned(reg403)) : reg405[(4'h9):(3'h4)])});
              reg480 = $signed((reg422 ?
                  reg472[(1'h0):(1'h0)] : (($signed(reg464) ?
                          $unsigned(reg436) : (reg460 ? reg404 : reg398)) ?
                      ($signed(reg414) * (~|forvar476)) : reg450)));
              reg481 <= reg424[(3'h6):(3'h4)];
            end
          if ($signed(reg430))
            begin
              reg482 <= (~forvar476[(5'h15):(1'h1)]);
              reg483 = $unsigned({reg405, reg458});
              reg484 <= $signed(reg453[(2'h2):(2'h2)]);
            end
          else
            begin
              reg483 = $signed(($unsigned(reg433) * reg404[(3'h6):(1'h1)]));
              reg484 <= reg469;
              reg485 <= reg468[(3'h4):(1'h0)];
              reg486 <= reg453;
              reg487 = $signed({(wire457 > reg422[(3'h7):(2'h3)])});
            end
          reg488 <= reg403;
          for (forvar489 = (1'h0); (forvar489 < (1'h1)); forvar489 = (forvar489 + (1'h1)))
            begin
              reg490 <= $signed($signed(reg398));
              reg491 <= ((~&(^reg484)) ? $signed(reg479) : wire386);
              reg492 = $signed($signed($signed(reg408)));
              reg493 <= reg400;
              reg494 <= reg483;
            end
          if ($signed(({(reg492[(5'h12):(4'ha)] ?
                      ((8'hb8) ~^ (8'ha4)) : reg465[(3'h6):(3'h6)])} ?
              (^$unsigned(((7'h41) | reg450))) : (((^~reg465) && $unsigned(reg431)) ?
                  (!$signed(reg398)) : reg430[(2'h3):(1'h1)]))))
            begin
              reg495 <= reg427;
            end
          else
            begin
              reg495 <= wire475;
              reg496 = ($unsigned((reg408 < reg481[(4'hb):(3'h5)])) <<< reg486[(1'h1):(1'h0)]);
              reg497 <= $signed($signed({(reg468 >>> {reg418})}));
              reg498 <= (({reg433[(2'h2):(1'h1)]} ?
                  {reg437[(3'h7):(3'h4)]} : ($signed($unsigned(reg433)) ?
                      (((8'hbb) ? reg409 : (8'hb1)) ?
                          $signed(reg416) : reg392[(2'h2):(1'h1)]) : ($unsigned(reg472) * $signed(reg424)))) - ($unsigned(reg449) << $signed($unsigned((wire457 ^ reg482)))));
            end
        end
    end
  always
    @(posedge clk) begin
      if (($signed($signed($unsigned(reg418))) ?
          (reg398[(4'h8):(2'h2)] || reg441[(1'h0):(1'h0)]) : $unsigned($signed((!reg481)))))
        begin
          for (forvar499 = (1'h0); (forvar499 < (1'h0)); forvar499 = (forvar499 + (1'h1)))
            begin
              reg500 <= (^~reg404[(4'h9):(3'h4)]);
              reg501 <= {reg453[(2'h2):(1'h1)], $unsigned(reg423)};
              reg502 = (^~((reg490 ?
                      $unsigned((reg423 ?
                          reg465 : wire385)) : (~&$signed(reg392))) ?
                  $signed(forvar499) : reg449[(3'h6):(3'h5)]));
            end
        end
      else
        begin
          reg499 = $signed(reg465);
        end
      reg503 = {{$signed(((&reg459) ? reg491 : (~(8'h9d))))}};
      for (forvar504 = (1'h0); (forvar504 < (3'h4)); forvar504 = (forvar504 + (1'h1)))
        begin
          reg505 = {($unsigned($unsigned($signed(reg427))) * $unsigned({(reg503 ?
                      (7'h46) : reg501)})),
              (+$unsigned(($unsigned(reg491) << (wire475 ? reg418 : reg398))))};
          if (reg405[(1'h0):(1'h0)])
            begin
              reg506 = ((($unsigned((~reg459)) ~^ reg458) ?
                      {(wire387[(3'h6):(1'h0)] ?
                              $unsigned(reg445) : $unsigned((7'h47))),
                          (^~(&reg490))} : reg413) ?
                  wire457 : $unsigned(reg394[(3'h6):(3'h5)]));
              reg507 <= ((&reg422) - (^$unsigned(reg490)));
              reg508 <= ($unsigned(wire384[(4'hf):(3'h7)]) ?
                  $signed(({reg502[(2'h3):(2'h3)]} ?
                      $unsigned((reg472 << (8'h9e))) : reg486)) : wire384);
            end
          else
            begin
              reg506 = (-{((reg449 ? reg436 : $unsigned(reg485)) ?
                      reg408 : reg488)});
            end
          reg509 <= (reg459 ?
              $unsigned($unsigned((8'hb8))) : $signed((reg468[(4'hd):(4'h9)] ?
                  {reg486[(3'h6):(3'h4)]} : (reg499 ^ {reg481, reg403}))));
        end
      if ((reg433 | reg506[(5'h15):(4'ha)]))
        begin
          for (forvar510 = (1'h0); (forvar510 < (2'h3)); forvar510 = (forvar510 + (1'h1)))
            begin
              reg511 = ($signed(reg426) ?
                  ((wire385 > wire454) | ({$signed(reg413)} ?
                      (!$unsigned(reg482)) : (~&reg450[(2'h3):(1'h0)]))) : $signed({reg509}));
            end
        end
      else
        begin
          reg510 <= $signed($signed(((^~reg422[(3'h7):(3'h7)]) ?
              ((+reg503) ?
                  (reg509 ? reg493 : (8'h9e)) : {reg485,
                      reg499}) : $unsigned({(8'ha1)}))));
          reg511 = wire455[(2'h3):(2'h3)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1317
#(parameter param1549 = {(({((8'h9c) ^ (8'hab))} >>> ({(8'hbf)} || {(8'ha2)})) | ((((8'hb8) & (8'ha1)) & ((8'ha8) || (7'h45))) ? {((8'h9e) <= (8'hae))} : ((-(8'ha4)) ? ((8'ha3) ? (8'hbb) : (7'h41)) : (^(8'ha0)))))})
(y, clk, wire1321, wire1320, wire1319, wire1318);
  output wire [(32'hb9a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire1321;
  input wire signed [(5'h15):(1'h0)] wire1320;
  input wire [(5'h14):(1'h0)] wire1319;
  input wire signed [(5'h11):(1'h0)] wire1318;
  wire signed [(3'h5):(1'h0)] wire1536;
  wire [(3'h6):(1'h0)] wire1535;
  wire signed [(3'h5):(1'h0)] wire1534;
  wire [(4'hf):(1'h0)] wire1390;
  wire signed [(4'ha):(1'h0)] wire1373;
  wire signed [(2'h3):(1'h0)] wire1353;
  wire [(4'h9):(1'h0)] wire1352;
  wire signed [(5'h15):(1'h0)] wire1334;
  wire [(5'h10):(1'h0)] wire1333;
  wire [(3'h6):(1'h0)] wire1331;
  wire [(4'ha):(1'h0)] wire1330;
  wire signed [(4'hc):(1'h0)] wire1325;
  reg [(4'hb):(1'h0)] reg1548 = (1'h0);
  reg [(4'hd):(1'h0)] reg1547 = (1'h0);
  reg [(5'h10):(1'h0)] reg1543 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1542 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1540 = (1'h0);
  reg [(2'h2):(1'h0)] reg1538 = (1'h0);
  reg [(5'h13):(1'h0)] reg1533 = (1'h0);
  reg [(5'h16):(1'h0)] reg1532 = (1'h0);
  reg [(5'h13):(1'h0)] reg1531 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1527 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1526 = (1'h0);
  reg [(4'hd):(1'h0)] reg1523 = (1'h0);
  reg [(5'h10):(1'h0)] reg1519 = (1'h0);
  reg [(4'hc):(1'h0)] reg1515 = (1'h0);
  reg [(4'ha):(1'h0)] reg1514 = (1'h0);
  reg [(3'h7):(1'h0)] reg1511 = (1'h0);
  reg [(5'h10):(1'h0)] reg1509 = (1'h0);
  reg [(5'h12):(1'h0)] reg1507 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1504 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1503 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1502 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1501 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1499 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1497 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1496 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1495 = (1'h0);
  reg [(5'h16):(1'h0)] reg1492 = (1'h0);
  reg [(4'hf):(1'h0)] reg1477 = (1'h0);
  reg [(4'h9):(1'h0)] reg1490 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1489 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1488 = (1'h0);
  reg [(4'hc):(1'h0)] reg1487 = (1'h0);
  reg [(4'hd):(1'h0)] reg1485 = (1'h0);
  reg [(5'h15):(1'h0)] reg1484 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1483 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1482 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1481 = (1'h0);
  reg [(4'hd):(1'h0)] reg1480 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1479 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1478 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1474 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1473 = (1'h0);
  reg [(4'hf):(1'h0)] reg1472 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1470 = (1'h0);
  reg [(5'h10):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1467 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1466 = (1'h0);
  reg [(3'h4):(1'h0)] reg1465 = (1'h0);
  reg [(5'h12):(1'h0)] reg1463 = (1'h0);
  reg [(4'ha):(1'h0)] reg1462 = (1'h0);
  reg [(3'h7):(1'h0)] reg1461 = (1'h0);
  reg [(3'h4):(1'h0)] reg1460 = (1'h0);
  reg [(4'h8):(1'h0)] reg1459 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1458 = (1'h0);
  reg [(5'h14):(1'h0)] reg1456 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1454 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1452 = (1'h0);
  reg [(4'he):(1'h0)] reg1444 = (1'h0);
  reg [(5'h15):(1'h0)] reg1450 = (1'h0);
  reg [(5'h18):(1'h0)] reg1448 = (1'h0);
  reg [(5'h12):(1'h0)] reg1445 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1443 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1442 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1441 = (1'h0);
  reg [(4'h9):(1'h0)] reg1439 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1436 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1435 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1433 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1432 = (1'h0);
  reg [(3'h5):(1'h0)] reg1429 = (1'h0);
  reg [(4'h9):(1'h0)] reg1428 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1424 = (1'h0);
  reg [(5'h13):(1'h0)] reg1423 = (1'h0);
  reg [(5'h12):(1'h0)] reg1422 = (1'h0);
  reg [(4'hb):(1'h0)] reg1420 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1419 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1417 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1416 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1415 = (1'h0);
  reg [(5'h14):(1'h0)] reg1414 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1412 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1403 = (1'h0);
  reg [(5'h14):(1'h0)] reg1401 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1399 = (1'h0);
  reg [(5'h16):(1'h0)] reg1396 = (1'h0);
  reg [(4'hd):(1'h0)] reg1395 = (1'h0);
  reg [(4'h8):(1'h0)] reg1389 = (1'h0);
  reg [(5'h14):(1'h0)] reg1388 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1387 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1386 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1385 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1382 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1375 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1372 = (1'h0);
  reg [(4'h9):(1'h0)] reg1371 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1369 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1366 = (1'h0);
  reg [(4'h9):(1'h0)] reg1365 = (1'h0);
  reg [(4'hf):(1'h0)] reg1362 = (1'h0);
  reg [(4'h9):(1'h0)] reg1360 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1359 = (1'h0);
  reg [(3'h7):(1'h0)] reg1357 = (1'h0);
  reg [(4'he):(1'h0)] reg1356 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1348 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1343 = (1'h0);
  reg [(2'h2):(1'h0)] reg1340 = (1'h0);
  reg [(4'hc):(1'h0)] reg1337 = (1'h0);
  reg [(4'h8):(1'h0)] reg1336 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1329 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1326 = (1'h0);
  reg [(2'h3):(1'h0)] reg1324 = (1'h0);
  reg [(4'hf):(1'h0)] reg1546 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1545 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1544 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1541 = (1'h0);
  reg [(3'h6):(1'h0)] reg1539 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1537 = (1'h0);
  reg [(3'h5):(1'h0)] reg1530 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1529 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1528 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1525 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1524 = (1'h0);
  reg [(2'h3):(1'h0)] reg1522 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1521 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1520 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1518 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1517 = (1'h0);
  reg [(4'hf):(1'h0)] reg1516 = (1'h0);
  reg [(5'h11):(1'h0)] reg1513 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1512 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1510 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1508 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1506 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1505 = (1'h0);
  reg [(4'h8):(1'h0)] reg1500 = (1'h0);
  reg [(5'h12):(1'h0)] reg1498 = (1'h0);
  reg [(4'h9):(1'h0)] reg1494 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1493 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1471 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1491 = (1'h0);
  reg [(5'h16):(1'h0)] reg1486 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1477 = (1'h0);
  reg [(2'h2):(1'h0)] reg1476 = (1'h0);
  reg [(5'h10):(1'h0)] reg1475 = (1'h0);
  reg [(5'h12):(1'h0)] reg1471 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1456 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1455 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1468 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1464 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1457 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1455 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1453 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1447 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1451 = (1'h0);
  reg [(4'ha):(1'h0)] reg1449 = (1'h0);
  reg [(3'h7):(1'h0)] reg1447 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1446 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1444 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1440 = (1'h0);
  reg [(3'h7):(1'h0)] reg1438 = (1'h0);
  reg [(5'h12):(1'h0)] reg1437 = (1'h0);
  reg [(3'h5):(1'h0)] reg1434 = (1'h0);
  reg [(5'h17):(1'h0)] reg1431 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1430 = (1'h0);
  reg [(3'h7):(1'h0)] reg1421 = (1'h0);
  reg [(2'h2):(1'h0)] reg1427 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1426 = (1'h0);
  reg [(2'h2):(1'h0)] reg1425 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1421 = (1'h0);
  reg [(3'h5):(1'h0)] reg1418 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1413 = (1'h0);
  reg [(5'h10):(1'h0)] reg1411 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1410 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1409 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1407 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1406 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1405 = (1'h0);
  reg [(2'h2):(1'h0)] reg1404 = (1'h0);
  reg [(5'h16):(1'h0)] reg1402 = (1'h0);
  reg [(5'h17):(1'h0)] reg1400 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1398 = (1'h0);
  reg [(5'h11):(1'h0)] reg1397 = (1'h0);
  reg [(4'hb):(1'h0)] reg1394 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1393 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1392 = (1'h0);
  reg [(4'he):(1'h0)] reg1391 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1383 = (1'h0);
  reg [(2'h3):(1'h0)] reg1381 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1380 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1379 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1378 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1377 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1376 = (1'h0);
  reg [(3'h5):(1'h0)] reg1374 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1370 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1368 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1367 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1361 = (1'h0);
  reg [(5'h10):(1'h0)] reg1364 = (1'h0);
  reg [(4'hf):(1'h0)] reg1363 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1361 = (1'h0);
  reg [(5'h10):(1'h0)] reg1358 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1355 = (1'h0);
  reg [(2'h2):(1'h0)] reg1354 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1351 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1350 = (1'h0);
  reg [(4'hd):(1'h0)] reg1349 = (1'h0);
  reg [(4'hd):(1'h0)] reg1347 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1346 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1345 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1338 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1344 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1342 = (1'h0);
  reg [(5'h18):(1'h0)] reg1341 = (1'h0);
  reg [(4'h8):(1'h0)] reg1339 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1338 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1335 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1332 = (1'h0);
  reg [(5'h18):(1'h0)] reg1328 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1327 = (1'h0);
  reg [(5'h12):(1'h0)] reg1323 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1322 = (1'h0);
  assign y = {wire1536,
                 wire1535,
                 wire1534,
                 wire1390,
                 wire1373,
                 wire1353,
                 wire1352,
                 wire1334,
                 wire1333,
                 wire1331,
                 wire1330,
                 wire1325,
                 reg1548,
                 reg1547,
                 reg1543,
                 reg1542,
                 reg1540,
                 reg1538,
                 reg1533,
                 reg1532,
                 reg1531,
                 reg1527,
                 reg1526,
                 reg1523,
                 reg1519,
                 reg1515,
                 reg1514,
                 reg1511,
                 reg1509,
                 reg1507,
                 reg1504,
                 reg1503,
                 reg1502,
                 reg1501,
                 reg1499,
                 reg1497,
                 reg1496,
                 reg1495,
                 reg1492,
                 reg1477,
                 reg1490,
                 reg1489,
                 reg1488,
                 reg1487,
                 reg1485,
                 reg1484,
                 reg1483,
                 reg1482,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1478,
                 reg1474,
                 reg1473,
                 reg1472,
                 reg1470,
                 reg1469,
                 reg1467,
                 reg1466,
                 reg1465,
                 reg1463,
                 reg1462,
                 reg1461,
                 reg1460,
                 reg1459,
                 reg1458,
                 reg1456,
                 reg1454,
                 reg1452,
                 reg1444,
                 reg1450,
                 reg1448,
                 reg1445,
                 reg1443,
                 reg1442,
                 reg1441,
                 reg1439,
                 reg1436,
                 reg1435,
                 reg1433,
                 reg1432,
                 reg1429,
                 reg1428,
                 reg1424,
                 reg1423,
                 reg1422,
                 reg1420,
                 reg1419,
                 reg1417,
                 reg1416,
                 reg1415,
                 reg1414,
                 reg1412,
                 reg1408,
                 reg1403,
                 reg1401,
                 reg1399,
                 reg1396,
                 reg1395,
                 reg1389,
                 reg1388,
                 reg1387,
                 reg1386,
                 reg1385,
                 reg1382,
                 reg1375,
                 reg1372,
                 reg1371,
                 reg1369,
                 reg1366,
                 reg1365,
                 reg1362,
                 reg1360,
                 reg1359,
                 reg1357,
                 reg1356,
                 reg1348,
                 reg1343,
                 reg1340,
                 reg1337,
                 reg1336,
                 reg1329,
                 reg1326,
                 reg1324,
                 reg1546,
                 reg1545,
                 reg1544,
                 forvar1541,
                 reg1539,
                 forvar1537,
                 reg1530,
                 forvar1529,
                 reg1528,
                 forvar1525,
                 reg1524,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1518,
                 reg1517,
                 reg1516,
                 reg1513,
                 reg1512,
                 forvar1510,
                 reg1508,
                 reg1506,
                 forvar1505,
                 reg1500,
                 reg1498,
                 reg1494,
                 forvar1493,
                 forvar1471,
                 reg1491,
                 reg1486,
                 forvar1477,
                 reg1476,
                 reg1475,
                 reg1471,
                 forvar1456,
                 reg1455,
                 forvar1468,
                 reg1464,
                 reg1457,
                 forvar1455,
                 reg1453,
                 forvar1447,
                 reg1451,
                 reg1449,
                 reg1447,
                 reg1446,
                 forvar1444,
                 reg1440,
                 reg1438,
                 reg1437,
                 reg1434,
                 reg1431,
                 reg1430,
                 reg1421,
                 reg1427,
                 reg1426,
                 reg1425,
                 forvar1421,
                 reg1418,
                 reg1413,
                 reg1411,
                 reg1410,
                 forvar1409,
                 forvar1407,
                 reg1406,
                 forvar1405,
                 reg1404,
                 reg1402,
                 reg1400,
                 reg1398,
                 reg1397,
                 reg1394,
                 forvar1393,
                 reg1392,
                 reg1391,
                 reg1384,
                 reg1383,
                 reg1381,
                 reg1380,
                 reg1379,
                 forvar1378,
                 forvar1377,
                 reg1376,
                 reg1374,
                 reg1370,
                 forvar1368,
                 reg1367,
                 reg1361,
                 reg1364,
                 reg1363,
                 forvar1361,
                 reg1358,
                 reg1355,
                 reg1354,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1347,
                 forvar1346,
                 forvar1345,
                 reg1338,
                 reg1344,
                 reg1342,
                 reg1341,
                 reg1339,
                 forvar1338,
                 reg1335,
                 reg1332,
                 reg1328,
                 reg1327,
                 reg1323,
                 reg1322,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1322 = ($unsigned((((+wire1320) < {wire1319}) >= {wire1318[(4'h8):(3'h7)],
              (~^(7'h40))})) ?
          $signed((8'ha7)) : {($signed($unsigned((8'ha0))) ?
                  ({wire1318} ?
                      $unsigned(wire1321) : wire1321[(3'h4):(3'h4)]) : $unsigned((8'had))),
              (((^~(8'hab)) >= (wire1320 ? (8'h9e) : wire1319)) ?
                  {$unsigned(wire1321)} : (((8'hbe) ^ wire1318) == wire1321[(5'h14):(4'hf)]))});
      reg1323 = (({wire1318} ?
              $signed(wire1320) : ((~|wire1319[(5'h10):(4'ha)]) * ({wire1319} ^~ (8'hb1)))) ?
          wire1319 : (+(~|({wire1319, wire1320} + $signed(reg1322)))));
      reg1324 <= ((&(wire1321 ?
          (8'haf) : ((wire1321 || wire1321) ?
              $signed(reg1323) : $unsigned(wire1320)))) & (|(~(^reg1322[(1'h1):(1'h0)]))));
    end
  assign wire1325 = wire1318;
  always
    @(posedge clk) begin
      reg1326 <= (-wire1325);
      reg1327 = (~(~($unsigned($unsigned(wire1318)) & $unsigned($unsigned(wire1321)))));
      reg1328 = $unsigned(($unsigned(((reg1327 == wire1321) | $signed((8'hb8)))) | ($signed((-wire1319)) >> reg1326[(2'h2):(1'h0)])));
      reg1329 <= $unsigned((~^$unsigned($signed((~|reg1326)))));
    end
  assign wire1330 = ($unsigned(((wire1318 & {wire1319}) ?
                            ((&(7'h44)) ?
                                $unsigned(reg1329) : $signed(reg1329)) : (&$unsigned(reg1326)))) ?
                        {reg1326, (8'ha4)} : {$signed(reg1326[(2'h3):(1'h0)]),
                            (~^{(~^(7'h47))})});
  assign wire1331 = (-(&$unsigned($signed($signed(wire1330)))));
  always
    @(posedge clk) begin
      reg1332 = (($signed((~|$signed(wire1321))) ?
              wire1331[(2'h2):(2'h2)] : wire1321[(4'h9):(1'h0)]) ?
          (~($unsigned((^reg1324)) ?
              $signed((wire1321 ?
                  wire1318 : wire1319)) : reg1326)) : $unsigned($unsigned($signed(wire1319[(4'ha):(3'h7)]))));
    end
  assign wire1333 = wire1321[(5'h12):(5'h12)];
  assign wire1334 = ((((~|$unsigned(wire1325)) ?
                                ($unsigned(reg1324) ^ $signed(wire1318)) : reg1324) ?
                            (($unsigned((8'hb0)) + {wire1331,
                                wire1321}) * ($signed(wire1333) | (wire1331 ?
                                wire1333 : wire1319))) : wire1333) ?
                        (wire1330 != ((reg1329[(4'ha):(4'h9)] != wire1319[(3'h6):(3'h5)]) ?
                            (-((8'ha0) >> reg1326)) : $signed((~^reg1324)))) : $unsigned((8'hae)));
  always
    @(posedge clk) begin
      if ($signed((~|$signed(reg1326[(2'h2):(1'h1)]))))
        begin
          reg1335 = $unsigned(wire1331[(1'h1):(1'h0)]);
          reg1336 <= ($signed(wire1330[(4'h9):(2'h2)]) ?
              $signed((~$unsigned(((7'h4a) << wire1331)))) : $signed((8'haa)));
          reg1337 <= wire1331;
          for (forvar1338 = (1'h0); (forvar1338 < (2'h2)); forvar1338 = (forvar1338 + (1'h1)))
            begin
              reg1339 = (wire1321[(4'hc):(4'h9)] ?
                  $signed(reg1335[(5'h11):(4'hf)]) : $unsigned(reg1324));
              reg1340 <= wire1321[(4'he):(3'h4)];
              reg1341 = reg1337[(4'hb):(3'h5)];
              reg1342 = reg1329[(4'ha):(3'h5)];
              reg1343 <= wire1331[(2'h3):(2'h2)];
            end
          reg1344 = ({(-reg1342)} ?
              {(wire1330[(2'h2):(1'h0)] ?
                      {$unsigned((8'ha4))} : (reg1335[(5'h13):(4'hf)] ?
                          (~|wire1320) : (!(8'hbf))))} : (+$unsigned((&(7'h48)))));
        end
      else
        begin
          if (((((~&(wire1331 ? reg1329 : wire1318)) ?
              (wire1325[(3'h6):(3'h4)] ?
                  $signed(reg1326) : {(8'hb7),
                      forvar1338}) : {(reg1326 >= wire1331),
                  $signed(reg1343)}) > (((reg1326 ? reg1344 : reg1326) ?
                  reg1344[(2'h2):(1'h1)] : {reg1326, reg1339}) ?
              (~|(reg1335 >> (8'hb2))) : (wire1321 >= (~&forvar1338)))) & (8'ha5)))
            begin
              reg1336 <= (({{reg1343[(2'h2):(1'h0)]},
                          {{wire1333, wire1321}, reg1326}} ?
                      wire1334[(3'h4):(2'h3)] : (~^{forvar1338, wire1321})) ?
                  ((!(8'ha8)) ?
                      (&reg1340) : $unsigned((+reg1336[(4'h8):(3'h5)]))) : $unsigned(reg1342[(1'h1):(1'h0)]));
            end
          else
            begin
              reg1336 <= (wire1319[(2'h3):(2'h3)] ?
                  ($signed($signed(reg1342)) && (wire1318 ?
                      $signed($unsigned((8'ha7))) : ($unsigned(reg1335) + reg1324[(1'h1):(1'h1)]))) : forvar1338[(2'h3):(1'h1)]);
              reg1337 <= (~&wire1321[(1'h1):(1'h0)]);
              reg1338 = $signed(reg1344[(2'h3):(2'h3)]);
              reg1339 = $unsigned($signed((~wire1333[(2'h2):(1'h1)])));
            end
        end
      for (forvar1345 = (1'h0); (forvar1345 < (1'h1)); forvar1345 = (forvar1345 + (1'h1)))
        begin
          for (forvar1346 = (1'h0); (forvar1346 < (3'h4)); forvar1346 = (forvar1346 + (1'h1)))
            begin
              reg1347 = $signed({wire1334[(4'h9):(2'h3)]});
              reg1348 <= (reg1337 <= $signed($unsigned(((~^reg1326) + (reg1347 + reg1337)))));
              reg1349 = (7'h47);
            end
          reg1350 = (7'h43);
          reg1351 = reg1336;
        end
    end
  assign wire1352 = reg1348[(2'h3):(2'h2)];
  assign wire1353 = ($unsigned(reg1348[(1'h1):(1'h1)]) ~^ (8'h9d));
  always
    @(posedge clk) begin
      if (($signed(reg1340[(1'h1):(1'h1)]) ?
          $unsigned(($signed($unsigned(reg1324)) ?
              wire1334 : $signed((wire1321 ?
                  wire1352 : reg1324)))) : $unsigned((-reg1337[(4'h9):(4'h8)]))))
        begin
          if ((8'hb1))
            begin
              reg1354 = (~&(!(|((wire1318 ? (8'h9f) : wire1321) ^ (wire1321 ?
                  (8'ha6) : reg1337)))));
              reg1355 = reg1343;
              reg1356 <= $unsigned({reg1355[(3'h5):(2'h2)]});
              reg1357 <= {reg1337[(3'h7):(1'h0)], reg1329};
              reg1358 = reg1354;
            end
          else
            begin
              reg1354 = wire1334;
              reg1355 = $signed(wire1352[(1'h1):(1'h1)]);
            end
          reg1359 <= reg1357[(1'h1):(1'h1)];
          if ($unsigned(wire1320))
            begin
              reg1360 <= $signed(((|((&reg1324) ?
                      (reg1355 == (7'h45)) : (wire1353 ? reg1343 : wire1321))) ?
                  $signed($signed($unsigned(wire1331))) : $signed($signed((wire1319 ?
                      reg1359 : reg1356)))));
            end
          else
            begin
              reg1360 <= $unsigned({$unsigned(((wire1334 ? wire1320 : reg1357) ?
                      (wire1330 ? reg1354 : wire1321) : $signed(wire1353)))});
            end
          for (forvar1361 = (1'h0); (forvar1361 < (2'h2)); forvar1361 = (forvar1361 + (1'h1)))
            begin
              reg1362 <= ($signed(($unsigned(reg1358) >>> (+(8'ha0)))) ?
                  reg1354[(1'h0):(1'h0)] : $signed((~$unsigned(wire1321[(4'ha):(3'h6)]))));
              reg1363 = ($unsigned(reg1326) ?
                  (reg1337[(4'hc):(4'hc)] ?
                      $unsigned(({reg1358,
                          reg1362} ^~ (reg1340 & wire1321))) : $unsigned(((^reg1348) ^~ (reg1329 ?
                          reg1326 : wire1319)))) : $signed(reg1356[(4'he):(4'ha)]));
              reg1364 = $unsigned(wire1319);
              reg1365 <= $unsigned((~{(reg1326 ?
                      (wire1334 ? reg1340 : reg1359) : (reg1324 < wire1334)),
                  (reg1348 ? {reg1364, (7'h45)} : wire1318[(4'ha):(2'h3)])}));
            end
          if ($signed(reg1365[(2'h2):(1'h0)]))
            begin
              reg1366 <= ({(forvar1361[(4'hb):(4'ha)] ?
                      ($signed(reg1329) >>> reg1355) : (reg1363 ?
                          $unsigned(forvar1361) : reg1343[(2'h2):(1'h0)]))} >>> ((&(8'hbb)) & ((^~$signed(reg1326)) ?
                  $unsigned({wire1334}) : ($signed(wire1320) ?
                      wire1320 : (reg1364 ? wire1330 : reg1358)))));
            end
          else
            begin
              reg1366 <= (($signed(reg1355[(3'h5):(1'h0)]) ?
                  reg1355 : ((((8'hbc) & reg1359) ?
                      (+(8'ha4)) : wire1352[(4'h9):(1'h0)]) - {wire1353[(1'h1):(1'h0)],
                      $signed(wire1319)})) != $signed($signed(reg1366[(3'h4):(2'h3)])));
            end
        end
      else
        begin
          if ((|wire1352))
            begin
              reg1354 = $unsigned({wire1333[(1'h0):(1'h0)]});
              reg1355 = $signed($unsigned(wire1325[(3'h7):(3'h7)]));
              reg1356 <= ({$unsigned(wire1352[(3'h5):(3'h4)])} ?
                  (-((wire1330 ?
                      $signed((8'haf)) : {reg1356}) + $signed({wire1334,
                      (8'hae)}))) : ($signed((~&{reg1337})) ?
                      reg1356[(3'h5):(2'h3)] : reg1360[(1'h0):(1'h0)]));
              reg1357 <= $signed($signed($unsigned($signed($unsigned(reg1343)))));
              reg1358 = {({wire1330,
                          ((reg1357 ?
                              reg1364 : forvar1361) || (reg1355 <<< reg1337))} ?
                      wire1330 : $unsigned(reg1360))};
            end
          else
            begin
              reg1356 <= (^~((8'hb3) ?
                  (|((reg1365 >> wire1321) * (reg1343 ^~ wire1319))) : reg1364[(1'h1):(1'h0)]));
            end
          if (wire1319[(1'h1):(1'h1)])
            begin
              reg1361 = reg1354[(1'h1):(1'h1)];
              reg1363 = (&(^~{$unsigned({reg1355, wire1330}),
                  {(reg1343 ? wire1352 : reg1358), (^~reg1348)}}));
              reg1364 = $unsigned($unsigned(({wire1334[(1'h1):(1'h0)]} ?
                  (8'hab) : reg1360[(2'h3):(1'h0)])));
              reg1365 <= (^$signed((reg1363[(3'h6):(2'h2)] ?
                  reg1343 : $signed((~|wire1320)))));
              reg1367 = {(-$signed($unsigned($signed((8'h9e)))))};
            end
          else
            begin
              reg1361 = wire1320[(5'h13):(5'h13)];
              reg1363 = $signed((reg1355[(3'h5):(1'h0)] ?
                  (|wire1319) : $unsigned(wire1353)));
              reg1365 <= $signed((~$unsigned((8'hbd))));
              reg1367 = $signed({($unsigned((~^wire1319)) ?
                      (~$unsigned(wire1353)) : $unsigned(reg1329[(3'h5):(2'h2)])),
                  (-reg1359[(1'h0):(1'h0)])});
            end
          for (forvar1368 = (1'h0); (forvar1368 < (1'h1)); forvar1368 = (forvar1368 + (1'h1)))
            begin
              reg1369 <= {$signed((($unsigned(reg1358) >= (reg1329 ^~ reg1356)) ~^ wire1320)),
                  reg1363[(4'hb):(3'h5)]};
              reg1370 = $signed((((^(wire1353 - wire1318)) + (|$signed(reg1340))) ^ ($signed(wire1330[(2'h2):(2'h2)]) + $signed(reg1358))));
              reg1371 <= $unsigned(reg1359);
            end
          reg1372 <= {wire1353};
        end
    end
  assign wire1373 = ($unsigned({{(~&reg1362),
                            $unsigned(wire1330)}}) << wire1353[(1'h1):(1'h0)]);
  always
    @(posedge clk) begin
      reg1374 = $signed($signed(reg1359[(2'h2):(1'h1)]));
      reg1375 <= $signed((((^$unsigned(wire1334)) ?
              $signed((reg1371 != wire1353)) : $signed(wire1373)) ?
          (~&((wire1373 ^~ reg1360) ?
              $signed(reg1365) : reg1371[(1'h1):(1'h1)])) : (8'ha4)));
      reg1376 = $unsigned(((8'h9e) ?
          (7'h46) : $unsigned({(wire1333 ? (8'h9e) : (7'h42))})));
      for (forvar1377 = (1'h0); (forvar1377 < (2'h2)); forvar1377 = (forvar1377 + (1'h1)))
        begin
          for (forvar1378 = (1'h0); (forvar1378 < (1'h1)); forvar1378 = (forvar1378 + (1'h1)))
            begin
              reg1379 = wire1319[(5'h11):(4'hc)];
              reg1380 = (~&{$unsigned(((reg1366 ? (8'had) : (8'hbd)) ?
                      {reg1326} : $unsigned(reg1357)))});
              reg1381 = reg1324;
            end
          reg1382 <= (({$unsigned(reg1371)} ?
                  (&($signed(forvar1378) ?
                      {reg1362} : $unsigned(reg1371))) : ((|(^~reg1375)) <<< (-reg1376))) ?
              wire1321[(5'h12):(2'h2)] : $signed($signed({(~^reg1329),
                  (&reg1359)})));
          reg1383 = $signed((reg1375 < reg1357[(3'h6):(3'h6)]));
          if (($signed(reg1356[(3'h7):(3'h5)]) ?
              reg1376 : (~{(wire1352 ?
                      $signed(reg1340) : (wire1321 ? (8'hac) : reg1365)),
                  $signed((+reg1337))})))
            begin
              reg1384 = wire1331;
            end
          else
            begin
              reg1385 <= (+$signed({((reg1384 ? reg1382 : wire1330) ?
                      $unsigned((8'haa)) : reg1384)}));
              reg1386 <= ($unsigned(reg1360[(3'h4):(1'h0)]) & (8'ha6));
              reg1387 <= ((reg1356 >> ((7'h43) ?
                  ((+reg1356) << $unsigned(forvar1377)) : wire1318)) + ((8'hae) >> $unsigned((!(~(8'ha9))))));
              reg1388 <= $signed(({wire1319[(4'hf):(4'hf)],
                      ((reg1383 > reg1371) ?
                          (reg1380 - forvar1377) : (reg1329 * reg1362))} ?
                  reg1383 : $signed((+(+wire1334)))));
            end
          reg1389 <= $unsigned($signed((reg1371[(4'h8):(3'h5)] ?
              ($signed(reg1326) ?
                  $unsigned(forvar1377) : forvar1377) : $unsigned({reg1380,
                  reg1387}))));
        end
    end
  assign wire1390 = {(-{($unsigned(reg1329) | (|wire1352)),
                            (((8'ha6) ? wire1318 : reg1362) >= (reg1359 ?
                                wire1321 : wire1320))})};
  always
    @(posedge clk) begin
      reg1391 = (({$signed(((8'hbb) - reg1371))} ?
          $unsigned(reg1386[(2'h2):(2'h2)]) : $unsigned(((wire1321 ~^ wire1373) ?
              ((7'h42) ?
                  wire1321 : reg1375) : wire1353[(2'h2):(1'h1)]))) || $signed(wire1321[(4'he):(3'h7)]));
      reg1392 = $unsigned({reg1385,
          (^($unsigned(reg1324) ? $signed(reg1360) : reg1366[(2'h2):(1'h0)]))});
      for (forvar1393 = (1'h0); (forvar1393 < (2'h2)); forvar1393 = (forvar1393 + (1'h1)))
        begin
          reg1394 = reg1388[(4'he):(1'h1)];
          if (($signed($unsigned(($signed(reg1388) && (reg1329 ?
                  reg1348 : reg1343)))) ?
              reg1387 : $unsigned((reg1337 ?
                  $signed($signed(reg1362)) : reg1359))))
            begin
              reg1395 <= $unsigned($signed((wire1325[(4'h9):(4'h8)] ?
                  {(reg1343 > (8'ha7))} : $unsigned(reg1385))));
              reg1396 <= $unsigned($signed((~^(wire1352 ?
                  (8'ha8) : $unsigned(wire1320)))));
              reg1397 = reg1386;
              reg1398 = (7'h40);
            end
          else
            begin
              reg1397 = (^$signed({reg1395, {$signed(reg1394), reg1357}}));
            end
          if ((((8'hb9) <<< (|reg1372[(1'h0):(1'h0)])) <<< reg1365[(2'h3):(1'h1)]))
            begin
              reg1399 <= wire1373;
            end
          else
            begin
              reg1399 <= ($signed($unsigned($signed($signed(reg1343)))) ?
                  $signed(($signed($unsigned(wire1330)) ?
                      $unsigned((7'h46)) : wire1330)) : wire1319[(1'h1):(1'h1)]);
              reg1400 = reg1336[(3'h5):(2'h3)];
              reg1401 <= wire1390[(4'hd):(3'h5)];
            end
          if ($signed((($unsigned((^wire1330)) >>> $signed(reg1362[(1'h0):(1'h0)])) == $unsigned(reg1371[(1'h0):(1'h0)]))))
            begin
              reg1402 = {$signed($unsigned(wire1325[(4'hc):(4'hb)]))};
              reg1403 <= ((~|(8'hb2)) ?
                  wire1331[(3'h4):(2'h3)] : (((7'h40) ?
                          $unsigned(reg1366[(1'h0):(1'h0)]) : wire1320) ?
                      wire1321 : $unsigned(((reg1360 ? reg1357 : reg1375) ?
                          ((8'ha1) + reg1329) : (reg1391 ?
                              reg1400 : reg1343)))));
            end
          else
            begin
              reg1402 = wire1331;
            end
        end
      reg1404 = {(7'h46)};
      for (forvar1405 = (1'h0); (forvar1405 < (1'h0)); forvar1405 = (forvar1405 + (1'h1)))
        begin
          reg1406 = (^(!$signed(reg1343)));
          for (forvar1407 = (1'h0); (forvar1407 < (1'h1)); forvar1407 = (forvar1407 + (1'h1)))
            begin
              reg1408 <= $signed($unsigned((reg1391 ?
                  reg1406[(3'h6):(3'h6)] : ($signed(reg1360) ?
                      (+reg1356) : (wire1321 >> reg1382)))));
            end
          for (forvar1409 = (1'h0); (forvar1409 < (1'h1)); forvar1409 = (forvar1409 + (1'h1)))
            begin
              reg1410 = reg1402;
              reg1411 = $unsigned($unsigned(((!reg1356) >> $unsigned(((8'ha5) <<< (8'ha4))))));
              reg1412 <= ($signed(wire1325[(3'h7):(3'h6)]) ?
                  ((+($signed(wire1334) ?
                          wire1320[(2'h2):(1'h0)] : (reg1408 ?
                              reg1411 : reg1396))) ?
                      (~^$unsigned(reg1388[(4'ha):(4'h8)])) : ({forvar1405[(1'h0):(1'h0)],
                              $signed(reg1371)} ?
                          (((8'ha5) && reg1403) ?
                              $unsigned(wire1319) : $signed(reg1392)) : (!(reg1403 ?
                              reg1387 : reg1411)))) : reg1343[(1'h0):(1'h0)]);
              reg1413 = $unsigned(wire1331[(3'h4):(1'h1)]);
            end
          if (reg1385[(3'h6):(2'h3)])
            begin
              reg1414 <= {reg1395[(3'h5):(3'h5)], wire1334[(5'h15):(4'he)]};
              reg1415 <= forvar1407;
              reg1416 <= reg1406;
              reg1417 <= $unsigned((reg1400[(4'h8):(3'h6)] ?
                  ((|(+reg1406)) > (8'hab)) : ((&reg1416) ?
                      wire1352[(1'h0):(1'h0)] : $unsigned((reg1404 != wire1318)))));
            end
          else
            begin
              reg1414 <= (+$unsigned($signed(($signed((8'ha0)) ?
                  reg1375[(2'h2):(2'h2)] : $signed(forvar1409)))));
              reg1415 <= ((-(reg1326[(2'h3):(1'h1)] - (^~(~^(7'h49))))) ~^ $unsigned(((~$unsigned(reg1336)) << {reg1329[(2'h3):(1'h0)]})));
              reg1418 = reg1414[(3'h7):(1'h1)];
              reg1419 <= $unsigned(((reg1369 ?
                      (wire1333[(4'hf):(3'h4)] ^ (reg1403 ?
                          reg1394 : forvar1407)) : ($unsigned(reg1410) << (forvar1405 < (8'haa)))) ?
                  reg1412[(1'h0):(1'h0)] : $unsigned(reg1357[(3'h5):(1'h1)])));
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned(($signed($unsigned({wire1330, reg1366})) ?
          (reg1326 ?
              ({reg1359,
                  reg1348} >= $unsigned(reg1359)) : wire1325[(4'hc):(3'h5)]) : wire1373[(3'h6):(1'h1)])))
        begin
          reg1420 <= reg1395;
          for (forvar1421 = (1'h0); (forvar1421 < (2'h2)); forvar1421 = (forvar1421 + (1'h1)))
            begin
              reg1422 <= $unsigned(reg1385);
              reg1423 <= wire1390;
              reg1424 <= ($unsigned(($signed({wire1331, wire1321}) ?
                  $unsigned({(8'h9d),
                      reg1412}) : reg1375)) == $unsigned(((wire1334 >= $signed(reg1362)) ?
                  (-reg1419) : (^(~reg1356)))));
              reg1425 = $unsigned(($signed(wire1330) ?
                  $unsigned($signed(wire1331[(3'h6):(1'h1)])) : (~|$unsigned($unsigned((8'hae))))));
              reg1426 = ($signed((reg1324 > (~&wire1325[(3'h7):(3'h6)]))) ?
                  {reg1422, (-(8'hb5))} : reg1408);
            end
          reg1427 = (!wire1353);
        end
      else
        begin
          reg1421 = $signed($signed((^~(reg1396[(4'ha):(4'h9)] ?
              reg1427[(1'h1):(1'h1)] : $unsigned(wire1333)))));
          reg1425 = wire1320[(5'h12):(5'h12)];
          if (($unsigned(reg1360) ?
              (((|(reg1385 - reg1348)) ?
                      $signed(reg1420[(2'h2):(2'h2)]) : (forvar1421 == reg1422)) ?
                  $unsigned((~&reg1389)) : (!{(8'hb1)})) : {($unsigned(reg1360[(3'h5):(1'h0)]) ^ ($unsigned(wire1373) & {reg1343}))}))
            begin
              reg1428 <= reg1375;
              reg1429 <= $unsigned({($unsigned($unsigned(reg1428)) >= ($signed((8'ha5)) > $signed(wire1373))),
                  ($unsigned((reg1403 ? reg1359 : reg1360)) ?
                      $signed(wire1331) : (^~$unsigned(reg1366)))});
            end
          else
            begin
              reg1426 = reg1372;
              reg1428 <= (reg1362 >= (|(+$unsigned(reg1424))));
              reg1429 <= reg1415;
            end
          if ($unsigned(wire1352[(4'h8):(1'h0)]))
            begin
              reg1430 = $unsigned({$unsigned((-reg1360))});
              reg1431 = $unsigned(wire1352[(3'h7):(2'h2)]);
              reg1432 <= (^~$signed($signed((~|reg1431[(2'h3):(2'h3)]))));
              reg1433 <= (&reg1396);
            end
          else
            begin
              reg1432 <= $signed((&(8'hab)));
              reg1433 <= wire1325;
            end
        end
      reg1434 = $unsigned(($signed(((&reg1415) == $signed(wire1325))) ?
          ($signed($unsigned((8'hbb))) ?
              (!reg1419) : (reg1389[(3'h4):(2'h3)] ?
                  $signed(reg1429) : {reg1343})) : $unsigned(wire1353)));
      if ((($unsigned(reg1426) && $unsigned(((^~reg1372) ?
              {reg1387, (8'ha7)} : reg1414[(5'h12):(2'h2)]))) ?
          reg1408 : wire1373))
        begin
          reg1435 <= (7'h47);
          reg1436 <= (($unsigned(($signed(wire1390) ?
                      {reg1387, reg1396} : {(8'ha3)})) ?
                  $signed({$unsigned(reg1432)}) : (({(8'hb9)} ?
                          ((8'hb6) ? wire1390 : (7'h45)) : $signed((8'hb0))) ?
                      ({(7'h41), (7'h4a)} ~^ {reg1420}) : reg1432)) ?
              (($unsigned($unsigned(reg1348)) < $signed($unsigned(reg1399))) >= ($signed(reg1382[(4'h9):(4'h8)]) ?
                  $unsigned((~reg1419)) : (8'ha9))) : $signed(($unsigned($unsigned(reg1336)) <<< $unsigned(reg1348))));
          reg1437 = $unsigned((wire1320[(4'hc):(3'h6)] ?
              $signed((reg1429[(1'h0):(1'h0)] ?
                  reg1387[(1'h1):(1'h1)] : (reg1336 <= wire1321))) : reg1422));
          if ($unsigned(reg1425))
            begin
              reg1438 = reg1366[(4'h8):(3'h6)];
              reg1439 <= $signed(($unsigned((8'h9f)) <<< reg1324[(2'h3):(2'h3)]));
            end
          else
            begin
              reg1438 = $signed(reg1408[(3'h7):(1'h0)]);
              reg1440 = (({{(reg1425 ? reg1359 : reg1401),
                          (wire1352 ? (8'hb0) : reg1359)},
                      wire1353} ?
                  (~|({reg1329} ?
                      (reg1359 ?
                          reg1420 : reg1423) : $signed(reg1357))) : ($signed((reg1387 >> wire1325)) ?
                      reg1422 : (reg1382[(1'h0):(1'h0)] ^ (reg1360 ?
                          reg1389 : (8'ha3))))) >= wire1330);
              reg1441 <= wire1373[(1'h0):(1'h0)];
              reg1442 <= (~|{$unsigned($unsigned(reg1326[(2'h2):(2'h2)]))});
            end
        end
      else
        begin
          if (reg1386[(4'h9):(1'h0)])
            begin
              reg1437 = (((reg1386[(2'h3):(1'h0)] ?
                      ($unsigned((8'hb3)) + (reg1435 ?
                          reg1440 : wire1330)) : reg1365) ?
                  $unsigned(((wire1334 ?
                      reg1395 : (8'hb7)) ~^ $signed(wire1325))) : ((~&(^forvar1421)) ?
                      (~|$signed(reg1417)) : {reg1436[(3'h7):(2'h3)]})) < reg1421);
            end
          else
            begin
              reg1437 = (reg1421 > $unsigned((+reg1428)));
              reg1439 <= ($signed(reg1356) ?
                  ({wire1330[(3'h6):(3'h5)]} != ({((8'haf) ? reg1420 : reg1389),
                      $signed(wire1325)} < $signed($unsigned(wire1330)))) : (7'h46));
              reg1441 <= {($unsigned((8'ha6)) ?
                      $unsigned($signed({reg1366, reg1433})) : reg1434)};
              reg1442 <= reg1371[(2'h3):(1'h1)];
              reg1443 <= $unsigned(wire1330);
            end
        end
      if (wire1331[(2'h3):(1'h0)])
        begin
          for (forvar1444 = (1'h0); (forvar1444 < (2'h3)); forvar1444 = (forvar1444 + (1'h1)))
            begin
              reg1445 <= wire1352;
              reg1446 = forvar1421;
              reg1447 = {reg1441[(2'h2):(1'h1)]};
              reg1448 <= wire1334;
            end
          reg1449 = $unsigned($unsigned((~(~^(reg1439 ? (7'h48) : reg1396)))));
          reg1450 <= reg1417;
          reg1451 = (^($unsigned($signed((^(8'hbc)))) ~^ $unsigned((-(reg1401 & wire1390)))));
        end
      else
        begin
          reg1444 <= reg1337[(4'hc):(2'h3)];
          reg1445 <= $signed(reg1439);
          reg1446 = reg1356[(1'h0):(1'h0)];
          for (forvar1447 = (1'h0); (forvar1447 < (2'h2)); forvar1447 = (forvar1447 + (1'h1)))
            begin
              reg1448 <= ((^(reg1399 ?
                  forvar1444 : $unsigned({(7'h47)}))) <<< (reg1442 ~^ $unsigned(((reg1382 << reg1372) ^ (+reg1360)))));
              reg1450 <= $signed($unsigned((8'haa)));
              reg1451 = (^~reg1416[(2'h3):(2'h2)]);
              reg1452 <= wire1318;
              reg1453 = (-(8'hb3));
            end
          reg1454 <= reg1415[(3'h7):(2'h2)];
        end
      if ((reg1428[(3'h4):(2'h3)] ?
          (^~$unsigned(reg1432[(5'h10):(1'h1)])) : reg1452))
        begin
          for (forvar1455 = (1'h0); (forvar1455 < (1'h0)); forvar1455 = (forvar1455 + (1'h1)))
            begin
              reg1456 <= {reg1444, $unsigned(reg1360)};
              reg1457 = forvar1444[(1'h1):(1'h1)];
            end
          reg1458 <= (^({(!(reg1442 ? reg1422 : (8'ha9))),
                  (~^reg1453[(4'hd):(2'h2)])} ?
              (reg1337[(4'ha):(4'ha)] | ($unsigned((8'hae)) ?
                  (reg1448 ? reg1417 : reg1431) : reg1446)) : {reg1454}));
          if (reg1348)
            begin
              reg1459 <= {(8'hb3),
                  (-(-(reg1348[(3'h4):(1'h1)] > (^~reg1395))))};
              reg1460 <= (&{$unsigned({reg1357, ((8'hbb) <<< reg1438)})});
              reg1461 <= (reg1438 * $unsigned(($signed((wire1390 | (7'h42))) ^ reg1385)));
              reg1462 <= reg1427[(2'h2):(1'h0)];
              reg1463 <= {(reg1453 ? reg1372[(3'h6):(1'h0)] : wire1321),
                  $unsigned(reg1433[(2'h2):(2'h2)])};
            end
          else
            begin
              reg1459 <= $signed($unsigned(reg1428[(3'h6):(3'h6)]));
              reg1464 = $signed({reg1340});
              reg1465 <= reg1434[(1'h1):(1'h0)];
              reg1466 <= reg1385[(2'h3):(1'h0)];
              reg1467 <= ($unsigned((reg1348 | (~|((8'ha8) < reg1403)))) <= (~^(((8'ha1) != {reg1454,
                      reg1386}) ?
                  (!(reg1348 ?
                      (8'hb3) : (7'h47))) : ($unsigned(reg1451) ^ ((8'ha5) ?
                      forvar1421 : reg1388)))));
            end
          for (forvar1468 = (1'h0); (forvar1468 < (3'h4)); forvar1468 = (forvar1468 + (1'h1)))
            begin
              reg1469 <= ((~|((7'h45) ?
                      $unsigned(reg1432) : $unsigned({reg1359, (8'ha1)}))) ?
                  {(8'h9d)} : (~(8'hb9)));
            end
          reg1470 <= $signed($unsigned($unsigned((^~(!reg1337)))));
        end
      else
        begin
          reg1455 = wire1390;
          for (forvar1456 = (1'h0); (forvar1456 < (2'h3)); forvar1456 = (forvar1456 + (1'h1)))
            begin
              reg1458 <= $signed(reg1401[(4'h9):(4'h9)]);
              reg1459 <= reg1348;
              reg1460 <= (~|reg1435);
              reg1464 = (~&($signed(reg1359) == $signed(reg1431)));
            end
          if (reg1454)
            begin
              reg1465 <= $signed($unsigned({$unsigned($unsigned(reg1389))}));
            end
          else
            begin
              reg1465 <= reg1420[(3'h7):(3'h6)];
              reg1466 <= ((8'hb7) >>> $unsigned($unsigned((8'ha0))));
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg1399[(3'h6):(1'h0)])
        begin
          if ((-(~$signed(reg1337))))
            begin
              reg1471 = $unsigned({$signed($signed((reg1399 ?
                      reg1454 : reg1357))),
                  reg1371});
              reg1472 <= ($signed($signed((reg1414 ~^ (~^reg1435)))) ?
                  $unsigned((^(reg1462 ?
                      (~&reg1465) : $signed(reg1386)))) : $signed(reg1442[(2'h3):(2'h2)]));
              reg1473 <= {reg1420};
              reg1474 <= $unsigned((reg1467 ?
                  (+(~|$unsigned(wire1318))) : reg1362));
              reg1475 = ($unsigned($signed({(reg1396 ? reg1435 : reg1371),
                      (-reg1469)})) ?
                  $unsigned($unsigned(((reg1357 < wire1325) ?
                      (reg1423 ^ reg1432) : (reg1343 ?
                          reg1343 : (8'ha7))))) : wire1333[(4'h8):(3'h7)]);
            end
          else
            begin
              reg1471 = $signed((~&{(-$unsigned(reg1399)),
                  $unsigned($unsigned((8'ha7)))}));
              reg1472 <= reg1469;
              reg1475 = reg1433[(1'h1):(1'h0)];
              reg1476 = $signed($signed((^~(7'h42))));
            end
          for (forvar1477 = (1'h0); (forvar1477 < (1'h0)); forvar1477 = (forvar1477 + (1'h1)))
            begin
              reg1478 <= $signed($signed(reg1441[(2'h2):(1'h0)]));
              reg1479 <= reg1467[(3'h4):(2'h2)];
              reg1480 <= ((~(({reg1423, wire1353} * (reg1452 ?
                          reg1474 : reg1465)) ?
                      ((reg1340 ? reg1448 : reg1474) ?
                          $signed(reg1458) : wire1353[(2'h2):(1'h0)]) : reg1478)) ?
                  $signed($signed(($signed(reg1472) <<< wire1319[(3'h4):(2'h3)]))) : (reg1474[(4'h8):(2'h2)] ?
                      reg1415[(2'h2):(1'h1)] : ({(~&reg1466)} <= reg1388)));
              reg1481 <= $signed((({reg1365} && (((7'h44) ?
                  (8'ha4) : wire1331) ^ {reg1444,
                  reg1452})) < reg1461[(1'h1):(1'h0)]));
              reg1482 <= $unsigned($unsigned((&$signed({reg1452, reg1448}))));
            end
          if ($unsigned((^~$unsigned((reg1471 ?
              $unsigned(reg1387) : $signed((7'h43)))))))
            begin
              reg1483 <= (^~((8'h9c) << ((8'hae) ?
                  (reg1371[(1'h0):(1'h0)] ?
                      (reg1478 & reg1459) : (^reg1360)) : $signed((reg1452 > reg1473)))));
              reg1484 <= (-$signed(wire1320));
              reg1485 <= (~&$unsigned($unsigned((reg1435 >= wire1353[(1'h1):(1'h1)]))));
              reg1486 = ($unsigned($signed(((wire1319 - reg1459) >> reg1336[(3'h5):(3'h5)]))) ^~ reg1459);
            end
          else
            begin
              reg1486 = $unsigned($signed(reg1369));
              reg1487 <= ((reg1429 ?
                      {(wire1373[(2'h2):(2'h2)] >> (wire1318 <<< reg1336))} : (^~{reg1414,
                          $signed(reg1460)})) ?
                  (!$signed($unsigned((reg1474 ?
                      wire1325 : (8'hbc))))) : $unsigned((^((forvar1477 ~^ wire1353) || reg1388))));
              reg1488 <= ((8'ha5) ?
                  ($unsigned($unsigned($signed(wire1320))) ?
                      $unsigned((reg1452[(2'h3):(1'h0)] - (reg1482 == (8'h9c)))) : wire1390) : $unsigned({reg1419}));
              reg1489 <= $signed($unsigned(((|(reg1450 ~^ reg1356)) ?
                  $unsigned((~^(8'h9c))) : (reg1461[(3'h4):(1'h1)] ~^ (~|reg1454)))));
              reg1490 <= (!(reg1336[(3'h4):(1'h1)] == (reg1465 ?
                  reg1479[(2'h2):(2'h2)] : ((reg1486 ? reg1442 : reg1460) ?
                      (~&reg1485) : $signed(reg1465)))));
            end
          reg1491 = $signed((reg1371[(3'h6):(2'h2)] * {$signed(reg1456[(3'h5):(3'h4)]),
              (reg1460 <= $unsigned((8'hbe)))}));
        end
      else
        begin
          for (forvar1471 = (1'h0); (forvar1471 < (1'h0)); forvar1471 = (forvar1471 + (1'h1)))
            begin
              reg1472 <= $unsigned($unsigned(($unsigned($signed(reg1366)) >> $signed(reg1419[(1'h1):(1'h0)]))));
              reg1475 = (($unsigned($signed($signed(reg1365))) ?
                      $unsigned(reg1372) : ($unsigned(wire1318[(4'hb):(4'h8)]) && reg1329[(3'h5):(1'h1)])) ?
                  reg1386 : $signed(($signed(reg1487) ~^ ((wire1333 || (8'hac)) ?
                      $unsigned(reg1472) : $signed(reg1469)))));
            end
          reg1477 <= (($unsigned(reg1415[(2'h3):(2'h3)]) - reg1329[(4'h8):(2'h3)]) ?
              reg1490 : (!$unsigned($unsigned((reg1459 ? reg1484 : reg1486)))));
        end
      reg1492 <= reg1433[(3'h5):(1'h0)];
      if ((({reg1460[(2'h3):(2'h3)],
              {(-reg1389)}} | (reg1343[(1'h0):(1'h0)] + ((reg1420 ?
              reg1359 : reg1454) == reg1417[(2'h3):(2'h3)]))) ?
          (reg1429[(1'h1):(1'h0)] && $unsigned(($signed(reg1371) ?
              $signed(reg1477) : (!reg1337)))) : reg1372[(4'h9):(3'h5)]))
        begin
          for (forvar1493 = (1'h0); (forvar1493 < (2'h2)); forvar1493 = (forvar1493 + (1'h1)))
            begin
              reg1494 = (+reg1484[(4'ha):(3'h4)]);
              reg1495 <= $unsigned(reg1483[(4'hd):(3'h4)]);
              reg1496 <= reg1460[(2'h2):(1'h1)];
              reg1497 <= $unsigned(((~((reg1450 ? reg1485 : reg1419) ?
                      (^(8'hbf)) : wire1334[(5'h14):(1'h1)])) ?
                  $unsigned({((8'ha2) ? reg1423 : reg1483),
                      (&reg1492)}) : reg1365));
            end
        end
      else
        begin
          for (forvar1493 = (1'h0); (forvar1493 < (2'h2)); forvar1493 = (forvar1493 + (1'h1)))
            begin
              reg1494 = reg1382[(3'h5):(1'h1)];
              reg1498 = reg1369[(1'h1):(1'h1)];
            end
          reg1499 <= reg1458[(4'hf):(4'he)];
          if ($signed(reg1417))
            begin
              reg1500 = (($unsigned(($signed(reg1491) ?
                  reg1419 : (reg1495 ~^ wire1321))) != {reg1492[(4'hf):(1'h0)]}) > $signed((^~wire1334[(4'hc):(4'h9)])));
            end
          else
            begin
              reg1500 = wire1320[(3'h4):(1'h1)];
              reg1501 <= (-(^~(|(wire1320 ?
                  reg1459[(2'h3):(2'h2)] : (reg1483 ? reg1492 : reg1357)))));
              reg1502 <= reg1472;
              reg1503 <= (&$unsigned(((wire1325 | $signed(reg1366)) ?
                  $unsigned(((7'h42) || reg1458)) : reg1448)));
            end
          reg1504 <= reg1428;
        end
    end
  always
    @(posedge clk) begin
      for (forvar1505 = (1'h0); (forvar1505 < (1'h1)); forvar1505 = (forvar1505 + (1'h1)))
        begin
          if ((&($unsigned($unsigned({(8'hbf)})) ?
              reg1419 : reg1454[(4'hc):(1'h1)])))
            begin
              reg1506 = reg1419;
              reg1507 <= $signed((&reg1424));
              reg1508 = $unsigned((~&(&{(reg1395 ? (8'hae) : reg1423),
                  (~|reg1433)})));
              reg1509 <= $signed($signed((8'hbd)));
            end
          else
            begin
              reg1507 <= reg1452;
              reg1509 <= reg1469;
            end
          for (forvar1510 = (1'h0); (forvar1510 < (2'h3)); forvar1510 = (forvar1510 + (1'h1)))
            begin
              reg1511 <= {$unsigned({{reg1340[(1'h0):(1'h0)],
                          $unsigned(reg1366)},
                      reg1463[(3'h7):(3'h4)]})};
              reg1512 = ($signed(reg1470) ?
                  $signed({reg1424[(4'h9):(4'h9)],
                      $signed(reg1499)}) : (8'h9d));
              reg1513 = (|{reg1484,
                  ($signed({reg1419, reg1439}) ?
                      (+reg1365) : reg1445[(4'ha):(4'h8)])});
            end
        end
      if ((~^(reg1467[(4'h9):(2'h2)] ~^ (&$unsigned(wire1334[(3'h6):(1'h1)])))))
        begin
          if (reg1507)
            begin
              reg1514 <= $unsigned((^reg1403[(4'h9):(1'h1)]));
              reg1515 <= (~&($unsigned({(reg1480 ?
                      reg1485 : reg1506)}) <= reg1482));
            end
          else
            begin
              reg1516 = reg1326[(1'h0):(1'h0)];
              reg1517 = (~^reg1324);
              reg1518 = reg1477[(2'h3):(2'h2)];
              reg1519 <= reg1445[(4'h8):(2'h3)];
            end
        end
      else
        begin
          reg1516 = reg1487[(4'h8):(1'h1)];
          if ((~^reg1360))
            begin
              reg1519 <= (^~((reg1488 ~^ reg1343[(2'h2):(1'h1)]) ?
                  (reg1422 && reg1401[(4'h9):(1'h0)]) : (-$unsigned(reg1458))));
              reg1520 = {reg1477[(4'hf):(4'hb)]};
              reg1521 = (-($signed(reg1520[(2'h2):(1'h1)]) ^~ reg1385[(4'hb):(3'h6)]));
              reg1522 = ((~^(((reg1441 >= reg1478) ?
                      $unsigned(reg1504) : reg1472) ?
                  reg1356[(1'h1):(1'h1)] : $unsigned(reg1458))) * ($unsigned($unsigned($signed(reg1470))) <<< reg1458[(4'h8):(4'h8)]));
            end
          else
            begin
              reg1519 <= ((reg1507 ?
                  reg1432[(5'h12):(3'h5)] : $unsigned(reg1492[(5'h12):(1'h0)])) << (8'ha1));
              reg1523 <= $signed((~^((!reg1483[(2'h2):(2'h2)]) != (reg1511 ?
                  (reg1513 & reg1336) : (wire1390 ^ reg1511)))));
              reg1524 = {($unsigned(((reg1492 ? (8'ha4) : reg1513) ?
                      ((7'h42) || (7'h46)) : wire1390[(4'hc):(1'h0)])) << reg1511),
                  (~^$unsigned((8'ha0)))};
            end
          for (forvar1525 = (1'h0); (forvar1525 < (1'h1)); forvar1525 = (forvar1525 + (1'h1)))
            begin
              reg1526 <= (-(~|(forvar1525[(4'hf):(4'h9)] ?
                  reg1497[(2'h2):(1'h0)] : ((reg1524 ? (8'ha8) : reg1485) ?
                      (+reg1461) : {reg1514}))));
              reg1527 <= (-{(($unsigned(reg1502) ?
                      (-reg1362) : (reg1483 | reg1360)) || {$unsigned(reg1512)}),
                  ($signed(reg1470) <<< $unsigned(reg1515))});
              reg1528 = ($signed(reg1504) ?
                  {reg1429[(3'h5):(2'h2)], reg1518} : {$signed(reg1387)});
            end
          for (forvar1529 = (1'h0); (forvar1529 < (2'h2)); forvar1529 = (forvar1529 + (1'h1)))
            begin
              reg1530 = $unsigned(reg1467[(3'h5):(2'h3)]);
              reg1531 <= reg1469[(3'h4):(1'h1)];
            end
          reg1532 <= ((^reg1518) ?
              reg1462 : ((~{(reg1422 ?
                      reg1524 : reg1366)}) - (reg1366 ~^ reg1435)));
        end
      reg1533 <= $signed(({(~{reg1337}), (-(reg1503 ~^ reg1516))} ?
          reg1375 : $signed({reg1497[(2'h3):(1'h0)]})));
    end
  assign wire1534 = (~^(reg1456[(3'h6):(1'h1)] == (reg1444[(3'h4):(1'h1)] - (^(-reg1408)))));
  assign wire1535 = (wire1390[(2'h3):(2'h3)] | reg1533[(3'h4):(3'h4)]);
  assign wire1536 = ($signed(((((8'hac) ? reg1515 : wire1325) ?
                        (reg1366 ?
                            (8'h9e) : reg1348) : (~|(8'hbb))) ~^ ($signed(reg1462) ?
                        (reg1365 ?
                            (7'h40) : reg1388) : {(8'hb3)}))) & ((reg1386 ?
                            reg1488 : $signed(reg1359)) ?
                        ({{wire1319}} ?
                            wire1534[(3'h4):(2'h3)] : wire1535) : reg1445[(4'hd):(2'h3)]));
  always
    @(posedge clk) begin
      for (forvar1537 = (1'h0); (forvar1537 < (3'h4)); forvar1537 = (forvar1537 + (1'h1)))
        begin
          reg1538 <= (7'h40);
          reg1539 = reg1360[(1'h0):(1'h0)];
          reg1540 <= (~|(~^$unsigned(($signed(reg1419) ~^ ((7'h43) ?
              reg1337 : reg1415)))));
          for (forvar1541 = (1'h0); (forvar1541 < (2'h2)); forvar1541 = (forvar1541 + (1'h1)))
            begin
              reg1542 <= ($signed(reg1533[(4'hb):(2'h3)]) + reg1375);
              reg1543 <= (~&{(&{$unsigned(reg1432)})});
              reg1544 = $signed((~^{((reg1456 != reg1514) > $unsigned((7'h44))),
                  $unsigned((~&reg1488))}));
              reg1545 = $unsigned(reg1488[(3'h6):(2'h3)]);
              reg1546 = $unsigned(((((+reg1470) ?
                          reg1482[(1'h0):(1'h0)] : (reg1443 ~^ reg1386)) ?
                      (((8'hbb) < reg1490) ?
                          {reg1444, reg1460} : $signed(reg1348)) : wire1319) ?
                  (|reg1415[(3'h6):(3'h4)]) : ((reg1533[(2'h3):(1'h1)] ?
                      {reg1467,
                          reg1474} : $unsigned(reg1443)) - {reg1336[(4'h8):(2'h3)],
                      (reg1442 <= reg1504)})));
            end
          reg1547 <= $unsigned(wire1334[(3'h7):(3'h5)]);
        end
      reg1548 <= reg1497[(2'h2):(2'h2)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1218
#(parameter param1289 = (!(8'hbf)))
(y, clk, wire1223, wire1222, wire1221, wire1220, wire1219);
  output wire [(32'h397):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire1223;
  input wire [(5'h18):(1'h0)] wire1222;
  input wire signed [(5'h16):(1'h0)] wire1221;
  input wire signed [(4'ha):(1'h0)] wire1220;
  input wire signed [(5'h12):(1'h0)] wire1219;
  wire [(5'h15):(1'h0)] wire1267;
  wire [(4'he):(1'h0)] wire1253;
  reg signed [(4'hb):(1'h0)] reg1286 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1285 = (1'h0);
  reg [(5'h11):(1'h0)] reg1284 = (1'h0);
  reg [(5'h16):(1'h0)] reg1283 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1281 = (1'h0);
  reg [(3'h6):(1'h0)] reg1279 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1277 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1276 = (1'h0);
  reg [(3'h7):(1'h0)] reg1273 = (1'h0);
  reg [(5'h12):(1'h0)] reg1272 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1271 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1270 = (1'h0);
  reg [(5'h15):(1'h0)] reg1266 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1265 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1255 = (1'h0);
  reg [(5'h11):(1'h0)] reg1264 = (1'h0);
  reg [(5'h13):(1'h0)] reg1263 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1262 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1258 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1257 = (1'h0);
  reg [(4'hc):(1'h0)] reg1246 = (1'h0);
  reg [(5'h15):(1'h0)] reg1249 = (1'h0);
  reg [(4'hf):(1'h0)] reg1248 = (1'h0);
  reg [(4'hc):(1'h0)] reg1247 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1245 = (1'h0);
  reg [(5'h11):(1'h0)] reg1244 = (1'h0);
  reg [(2'h2):(1'h0)] reg1241 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1235 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1230 = (1'h0);
  reg [(3'h6):(1'h0)] reg1228 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1226 = (1'h0);
  reg [(4'ha):(1'h0)] reg1288 = (1'h0);
  reg [(3'h7):(1'h0)] reg1287 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1282 = (1'h0);
  reg [(4'h9):(1'h0)] reg1280 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1282 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1280 = (1'h0);
  reg [(5'h16):(1'h0)] reg1278 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1275 = (1'h0);
  reg [(3'h6):(1'h0)] reg1274 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1269 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1268 = (1'h0);
  reg [(2'h3):(1'h0)] reg1261 = (1'h0);
  reg [(4'hf):(1'h0)] reg1260 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1259 = (1'h0);
  reg [(2'h3):(1'h0)] reg1256 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1255 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1254 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1252 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1251 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1250 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1246 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1243 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1242 = (1'h0);
  reg [(4'hb):(1'h0)] reg1240 = (1'h0);
  reg [(2'h3):(1'h0)] reg1239 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1238 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1237 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1236 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1234 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1233 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1232 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1231 = (1'h0);
  reg [(3'h7):(1'h0)] reg1229 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1224 = (1'h0);
  reg [(5'h18):(1'h0)] reg1227 = (1'h0);
  reg [(4'hd):(1'h0)] reg1225 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1224 = (1'h0);
  assign y = {wire1267,
                 wire1253,
                 reg1286,
                 reg1285,
                 reg1284,
                 reg1283,
                 reg1281,
                 reg1279,
                 reg1277,
                 reg1276,
                 reg1273,
                 reg1272,
                 reg1271,
                 reg1270,
                 reg1266,
                 reg1265,
                 reg1255,
                 reg1264,
                 reg1263,
                 reg1262,
                 reg1258,
                 reg1257,
                 reg1246,
                 reg1249,
                 reg1248,
                 reg1247,
                 reg1245,
                 reg1244,
                 reg1241,
                 reg1235,
                 reg1230,
                 reg1228,
                 reg1226,
                 reg1288,
                 reg1287,
                 forvar1282,
                 reg1280,
                 reg1282,
                 forvar1280,
                 reg1278,
                 reg1275,
                 reg1274,
                 forvar1269,
                 forvar1268,
                 reg1261,
                 reg1260,
                 forvar1259,
                 reg1256,
                 forvar1255,
                 reg1254,
                 reg1252,
                 reg1251,
                 reg1250,
                 forvar1246,
                 reg1243,
                 reg1242,
                 reg1240,
                 reg1239,
                 reg1238,
                 reg1237,
                 forvar1236,
                 reg1234,
                 forvar1233,
                 reg1232,
                 reg1231,
                 reg1229,
                 forvar1224,
                 reg1227,
                 reg1225,
                 reg1224,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (($signed($unsigned((~wire1221[(3'h7):(3'h7)]))) ?
          $signed(wire1223) : (|$unsigned(((wire1221 ? wire1221 : wire1221) ?
              wire1223[(3'h6):(1'h0)] : {wire1219})))))
        begin
          reg1224 = (!(wire1219 && wire1223[(4'hf):(4'ha)]));
          reg1225 = $unsigned(wire1221);
          reg1226 <= ($signed((wire1222[(1'h0):(1'h0)] <<< {(^(8'hb0))})) ^ (~|$unsigned((~&(reg1225 >>> wire1222)))));
          reg1227 = wire1221;
        end
      else
        begin
          for (forvar1224 = (1'h0); (forvar1224 < (2'h2)); forvar1224 = (forvar1224 + (1'h1)))
            begin
              reg1225 = (^wire1220[(4'h8):(2'h2)]);
            end
          reg1226 <= $signed($signed(($signed((reg1227 >> wire1223)) >> (wire1221 ?
              (&(8'hbd)) : reg1225[(1'h1):(1'h0)]))));
          if ($unsigned((wire1220[(1'h1):(1'h0)] <<< forvar1224)))
            begin
              reg1228 <= (-$signed(($unsigned(reg1225[(4'h8):(3'h6)]) ?
                  (wire1222[(5'h13):(3'h5)] ?
                      reg1224 : wire1220[(4'h8):(3'h6)]) : ((wire1223 | reg1225) ?
                      (wire1219 ? wire1220 : wire1223) : (wire1220 ?
                          wire1221 : wire1222)))));
            end
          else
            begin
              reg1228 <= $unsigned(reg1228[(3'h4):(2'h2)]);
              reg1229 = ($signed({reg1228}) ?
                  (!($signed($unsigned(wire1220)) ?
                      (!(~^wire1221)) : $unsigned($unsigned(forvar1224)))) : ((^~(reg1227[(5'h13):(2'h2)] ?
                      (reg1225 & (8'hb9)) : wire1219[(3'h4):(2'h2)])) << reg1228));
              reg1230 <= (~|($unsigned({$unsigned(reg1229),
                  {(8'ha0)}}) >= $signed({$signed(wire1219), (~reg1228)})));
              reg1231 = (($unsigned($unsigned((wire1220 ?
                      wire1223 : reg1229))) ?
                  wire1221 : reg1225) > (($unsigned((reg1225 ?
                          reg1224 : wire1220)) ?
                      $signed($signed((8'h9e))) : ($signed(wire1223) || (~^reg1225))) ?
                  $signed(reg1225[(4'hc):(4'hc)]) : $signed(wire1223)));
            end
          reg1232 = reg1230[(2'h2):(2'h2)];
          for (forvar1233 = (1'h0); (forvar1233 < (2'h2)); forvar1233 = (forvar1233 + (1'h1)))
            begin
              reg1234 = ($unsigned(reg1229) >> (~^{(8'ha7)}));
              reg1235 <= $signed($signed(({$unsigned(reg1231),
                  $signed(reg1227)} ^ (8'hb8))));
            end
        end
      for (forvar1236 = (1'h0); (forvar1236 < (1'h1)); forvar1236 = (forvar1236 + (1'h1)))
        begin
          reg1237 = (!(reg1234[(4'hb):(3'h7)] >>> (reg1225[(1'h1):(1'h1)] <<< ((-reg1235) ?
              (|wire1222) : (^~reg1231)))));
        end
      if ($signed(reg1237[(1'h1):(1'h1)]))
        begin
          if (($unsigned((&$signed((reg1224 ?
              reg1235 : (8'haf))))) | (+(8'haa))))
            begin
              reg1238 = reg1234[(4'h9):(4'h9)];
            end
          else
            begin
              reg1238 = {((((forvar1233 ?
                      wire1219 : wire1221) ~^ $signed(reg1225)) != wire1223) && (8'hbe)),
                  forvar1224};
              reg1239 = $signed(reg1237[(3'h4):(2'h3)]);
              reg1240 = forvar1224;
              reg1241 <= (8'ha5);
              reg1242 = reg1237;
            end
          reg1243 = ($unsigned((((|(8'ha2)) ?
                      $unsigned(wire1223) : {reg1226, reg1242}) ?
                  reg1240 : reg1230)) ?
              (~^(reg1242 ?
                  $unsigned((reg1237 - reg1237)) : (wire1222 ?
                      wire1219 : $unsigned(reg1239)))) : (forvar1236[(1'h0):(1'h0)] ?
                  (&wire1223[(1'h0):(1'h0)]) : $unsigned(reg1228[(2'h3):(2'h3)])));
        end
      else
        begin
          reg1238 = (((8'h9d) ?
                  $unsigned({$signed(reg1231),
                      reg1226[(3'h5):(2'h3)]}) : reg1238[(4'h8):(3'h4)]) ?
              $unsigned(reg1234[(2'h2):(2'h2)]) : (!$unsigned(({reg1238,
                      wire1220} ?
                  reg1239 : $signed(reg1224)))));
          reg1241 <= reg1234;
          reg1242 = (reg1235[(2'h3):(1'h1)] ?
              (wire1219[(4'ha):(1'h0)] ?
                  $signed(($unsigned(reg1241) + (-reg1225))) : (reg1241[(2'h2):(2'h2)] ?
                      (reg1226[(5'h13):(5'h13)] ~^ (reg1230 ?
                          wire1219 : reg1225)) : reg1232[(4'h8):(3'h7)])) : (8'h9d));
          reg1244 <= $unsigned(((forvar1224 ^ ((forvar1224 ?
              reg1243 : (8'h9f)) * {(8'haf), reg1228})) ~^ (reg1224 ?
              ($signed(forvar1236) ^ (reg1242 * reg1239)) : ($unsigned(reg1239) ?
                  $signed(reg1232) : {reg1239}))));
        end
      if (reg1244[(4'h9):(3'h4)])
        begin
          reg1245 <= $unsigned($unsigned(($unsigned($unsigned(wire1222)) ?
              (8'ha6) : ((reg1237 ? forvar1236 : forvar1224) ?
                  forvar1224 : (reg1242 ? reg1244 : (8'hbc))))));
          for (forvar1246 = (1'h0); (forvar1246 < (3'h4)); forvar1246 = (forvar1246 + (1'h1)))
            begin
              reg1247 <= $unsigned(forvar1236);
              reg1248 <= $unsigned(((($signed(reg1247) ?
                      (~|reg1244) : reg1229) <<< $signed((reg1245 ?
                      wire1221 : reg1238))) ?
                  (^~forvar1233[(3'h6):(1'h1)]) : reg1228));
            end
          reg1249 <= reg1237[(5'h12):(4'hf)];
        end
      else
        begin
          if (forvar1224[(2'h2):(2'h2)])
            begin
              reg1245 <= reg1227;
            end
          else
            begin
              reg1245 <= {forvar1233[(4'h8):(3'h6)],
                  (reg1234 ?
                      reg1248 : {forvar1246[(2'h2):(1'h1)],
                          ({(8'ha3)} ~^ (reg1231 ? forvar1233 : reg1242))})};
              reg1246 <= $signed($unsigned((-wire1219[(4'h9):(3'h6)])));
              reg1250 = (7'h42);
              reg1251 = $unsigned({(reg1231 ~^ reg1224),
                  $signed(reg1238[(3'h7):(1'h1)])});
              reg1252 = reg1241;
            end
        end
    end
  assign wire1253 = (~$signed({$unsigned($unsigned(reg1235))}));
  always
    @(posedge clk) begin
      reg1254 = ((8'hb5) <<< reg1244[(1'h0):(1'h0)]);
      if ((((reg1244[(1'h1):(1'h0)] | reg1247) == wire1222[(5'h18):(4'hf)]) ?
          wire1253[(4'he):(3'h4)] : reg1254))
        begin
          for (forvar1255 = (1'h0); (forvar1255 < (1'h0)); forvar1255 = (forvar1255 + (1'h1)))
            begin
              reg1256 = (+reg1248[(2'h3):(1'h0)]);
              reg1257 <= (wire1220[(3'h7):(2'h3)] ?
                  $unsigned((reg1230[(2'h2):(2'h2)] ?
                      ({reg1235} || {reg1228, wire1222}) : ($signed(wire1219) ?
                          wire1221 : reg1235[(3'h7):(3'h4)]))) : {{reg1254,
                          (reg1254[(5'h10):(4'h8)] * reg1248[(3'h5):(1'h1)])},
                      wire1222[(2'h3):(2'h2)]});
            end
          reg1258 <= $signed(reg1246);
          for (forvar1259 = (1'h0); (forvar1259 < (2'h3)); forvar1259 = (forvar1259 + (1'h1)))
            begin
              reg1260 = ((^(wire1220 || wire1219[(5'h10):(4'hb)])) + forvar1255);
              reg1261 = ($signed(reg1248) ? reg1257 : wire1220);
              reg1262 <= (8'hb7);
              reg1263 <= reg1228[(3'h4):(3'h4)];
            end
          reg1264 <= reg1248;
        end
      else
        begin
          reg1255 <= $unsigned(reg1264[(3'h6):(3'h5)]);
        end
      reg1265 <= reg1264;
      reg1266 <= (reg1245 | (7'h41));
    end
  assign wire1267 = (reg1266[(4'ha):(1'h0)] ~^ $signed({reg1241[(1'h0):(1'h0)],
                        ((~&reg1258) ? $unsigned(reg1246) : (+wire1220))}));
  always
    @(posedge clk) begin
      for (forvar1268 = (1'h0); (forvar1268 < (2'h3)); forvar1268 = (forvar1268 + (1'h1)))
        begin
          for (forvar1269 = (1'h0); (forvar1269 < (1'h1)); forvar1269 = (forvar1269 + (1'h1)))
            begin
              reg1270 <= $unsigned((8'hbf));
              reg1271 <= (reg1246 && $unsigned(reg1264));
            end
          if ($signed(reg1246[(3'h5):(2'h2)]))
            begin
              reg1272 <= reg1264;
            end
          else
            begin
              reg1272 <= (^~reg1262[(4'hd):(4'h8)]);
              reg1273 <= wire1253[(3'h6):(2'h3)];
              reg1274 = $unsigned($unsigned({reg1264[(1'h0):(1'h0)],
                  (((7'h49) >>> wire1267) ?
                      forvar1268[(4'hd):(2'h3)] : {(8'h9d), reg1263})}));
            end
          reg1275 = (~&$unsigned(wire1223[(4'hb):(3'h6)]));
          if ((wire1222 || (reg1246[(4'ha):(2'h2)] == (~^reg1264))))
            begin
              reg1276 <= reg1271[(3'h4):(3'h4)];
            end
          else
            begin
              reg1276 <= $signed({(^~reg1262),
                  (reg1241 ?
                      ((^~reg1226) ?
                          $unsigned((8'hb8)) : $signed((8'ha7))) : $signed($unsigned(reg1258)))});
              reg1277 <= $unsigned(wire1222);
              reg1278 = (wire1253 || $unsigned(reg1255));
            end
          reg1279 <= $signed((^~$signed(reg1255[(2'h3):(2'h2)])));
        end
      if ($unsigned($signed((reg1246[(3'h5):(2'h3)] ?
          ($signed(reg1245) ?
              (reg1264 >= (8'hb5)) : reg1273[(3'h5):(1'h1)]) : $unsigned((reg1246 ?
              reg1228 : reg1245))))))
        begin
          for (forvar1280 = (1'h0); (forvar1280 < (2'h3)); forvar1280 = (forvar1280 + (1'h1)))
            begin
              reg1281 <= $signed(reg1277);
              reg1282 = ((-{forvar1268[(5'h11):(2'h3)]}) - (8'hab));
            end
        end
      else
        begin
          if ($unsigned(reg1272))
            begin
              reg1280 = $unsigned(($unsigned($signed($signed(reg1258))) <= reg1282));
            end
          else
            begin
              reg1280 = ($signed((({reg1249, reg1280} >= $unsigned(reg1276)) ?
                  (((8'hb9) & wire1267) && $signed(reg1235)) : $signed($signed(wire1222)))) && $signed((&(&(reg1273 ?
                  reg1258 : wire1219)))));
              reg1281 <= $signed(forvar1269);
            end
          for (forvar1282 = (1'h0); (forvar1282 < (3'h4)); forvar1282 = (forvar1282 + (1'h1)))
            begin
              reg1283 <= reg1281;
              reg1284 <= {(reg1258 ?
                      {$unsigned(forvar1268), reg1272} : ((~(^~reg1247)) ?
                          (~(~&(7'h41))) : (wire1253[(4'h8):(2'h3)] && (~&(8'hb8))))),
                  (($signed($signed(reg1275)) >> ($unsigned(reg1274) ~^ (reg1273 ?
                      reg1281 : reg1246))) && (($unsigned((8'hbc)) <<< $unsigned(reg1235)) >>> (|(reg1273 ?
                      reg1244 : reg1282))))};
            end
          reg1285 <= ((7'h42) ? (~^forvar1280) : wire1222[(4'h8):(3'h5)]);
        end
      reg1286 <= reg1266;
      reg1287 = (8'hb4);
      reg1288 = (({reg1273,
              $unsigned((reg1265 <<< reg1281))} <= $unsigned($signed($unsigned(reg1274)))) ?
          (~((-reg1228[(1'h0):(1'h0)]) == {reg1241[(2'h2):(2'h2)]})) : (8'hb4));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module857
#(parameter param1056 = (^~((({(7'h40), (7'h43)} || {(8'haa), (8'hb8)}) ? ((+(8'hbd)) < {(8'hbb)}) : ({(8'h9f)} ? (|(8'hba)) : ((8'ha6) && (8'ha7)))) ? (^~({(8'hbb)} || ((8'ha8) >= (8'ha2)))) : (+{{(8'hab)}}))))
(y, clk, wire861, wire860, wire859, wire858);
  output wire [(32'ha0c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire861;
  input wire signed [(4'hb):(1'h0)] wire860;
  input wire [(3'h7):(1'h0)] wire859;
  input wire [(5'h17):(1'h0)] wire858;
  wire signed [(3'h6):(1'h0)] wire1055;
  wire [(3'h5):(1'h0)] wire1054;
  wire [(5'h10):(1'h0)] wire1053;
  wire [(2'h2):(1'h0)] wire1052;
  wire [(4'hc):(1'h0)] wire1051;
  wire signed [(5'h10):(1'h0)] wire1043;
  wire [(2'h2):(1'h0)] wire1036;
  wire signed [(4'hf):(1'h0)] wire1001;
  wire signed [(3'h7):(1'h0)] wire1000;
  wire signed [(3'h4):(1'h0)] wire982;
  wire signed [(5'h16):(1'h0)] wire951;
  wire signed [(5'h11):(1'h0)] wire863;
  wire signed [(5'h14):(1'h0)] wire862;
  reg signed [(3'h7):(1'h0)] reg1045 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1049 = (1'h0);
  reg [(3'h6):(1'h0)] reg1047 = (1'h0);
  reg [(4'h9):(1'h0)] reg1038 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1035 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1034 = (1'h0);
  reg [(5'h17):(1'h0)] reg1031 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1028 = (1'h0);
  reg [(3'h6):(1'h0)] reg1027 = (1'h0);
  reg [(3'h7):(1'h0)] reg1025 = (1'h0);
  reg [(5'h15):(1'h0)] reg1023 = (1'h0);
  reg [(5'h18):(1'h0)] reg1021 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1016 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1019 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1018 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1017 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1015 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1014 = (1'h0);
  reg [(3'h6):(1'h0)] reg1011 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1009 = (1'h0);
  reg [(3'h4):(1'h0)] reg1006 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1004 = (1'h0);
  reg [(5'h16):(1'h0)] reg998 = (1'h0);
  reg [(2'h3):(1'h0)] reg997 = (1'h0);
  reg [(5'h14):(1'h0)] reg995 = (1'h0);
  reg [(3'h5):(1'h0)] reg994 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg993 = (1'h0);
  reg [(5'h12):(1'h0)] reg991 = (1'h0);
  reg [(3'h4):(1'h0)] reg989 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg986 = (1'h0);
  reg [(5'h14):(1'h0)] reg984 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg983 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg979 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg978 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg977 = (1'h0);
  reg signed [(4'he):(1'h0)] reg974 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg973 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg968 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg966 = (1'h0);
  reg [(4'hd):(1'h0)] reg965 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg964 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg963 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg961 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg960 = (1'h0);
  reg [(2'h3):(1'h0)] reg959 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg957 = (1'h0);
  reg [(5'h15):(1'h0)] reg948 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg947 = (1'h0);
  reg [(5'h18):(1'h0)] reg946 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg945 = (1'h0);
  reg [(2'h2):(1'h0)] reg944 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg940 = (1'h0);
  reg [(5'h18):(1'h0)] reg938 = (1'h0);
  reg [(2'h2):(1'h0)] reg934 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg933 = (1'h0);
  reg [(2'h2):(1'h0)] reg930 = (1'h0);
  reg [(2'h3):(1'h0)] reg927 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg926 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg923 = (1'h0);
  reg [(4'hc):(1'h0)] reg922 = (1'h0);
  reg [(4'hc):(1'h0)] reg921 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg918 = (1'h0);
  reg [(4'hd):(1'h0)] reg917 = (1'h0);
  reg [(4'h9):(1'h0)] reg916 = (1'h0);
  reg [(3'h7):(1'h0)] reg914 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg911 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg907 = (1'h0);
  reg [(4'hd):(1'h0)] reg906 = (1'h0);
  reg [(4'hc):(1'h0)] reg903 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg901 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg899 = (1'h0);
  reg signed [(4'he):(1'h0)] reg898 = (1'h0);
  reg [(4'h9):(1'h0)] reg897 = (1'h0);
  reg [(4'hd):(1'h0)] reg892 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg891 = (1'h0);
  reg [(3'h6):(1'h0)] reg888 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg886 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg885 = (1'h0);
  reg [(3'h4):(1'h0)] reg883 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg882 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg879 = (1'h0);
  reg [(4'he):(1'h0)] reg878 = (1'h0);
  reg [(5'h12):(1'h0)] reg876 = (1'h0);
  reg [(5'h10):(1'h0)] reg875 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg872 = (1'h0);
  reg [(5'h16):(1'h0)] reg871 = (1'h0);
  reg [(4'hc):(1'h0)] reg869 = (1'h0);
  reg [(4'h9):(1'h0)] reg867 = (1'h0);
  reg [(4'hf):(1'h0)] reg864 = (1'h0);
  reg [(4'h9):(1'h0)] reg1048 = (1'h0);
  reg [(3'h7):(1'h0)] reg1050 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1048 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1046 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1045 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1044 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1042 = (1'h0);
  reg [(4'he):(1'h0)] reg1041 = (1'h0);
  reg [(5'h15):(1'h0)] reg1040 = (1'h0);
  reg [(4'hd):(1'h0)] reg1039 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1037 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1033 = (1'h0);
  reg [(5'h17):(1'h0)] reg1032 = (1'h0);
  reg [(4'hd):(1'h0)] reg1030 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1029 = (1'h0);
  reg [(3'h6):(1'h0)] reg1026 = (1'h0);
  reg [(4'hf):(1'h0)] reg1024 = (1'h0);
  reg [(4'he):(1'h0)] reg1022 = (1'h0);
  reg [(5'h18):(1'h0)] reg1020 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1016 = (1'h0);
  reg [(3'h5):(1'h0)] reg1013 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1012 = (1'h0);
  reg [(4'hf):(1'h0)] reg1010 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1008 = (1'h0);
  reg [(3'h7):(1'h0)] reg1007 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1005 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1003 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1002 = (1'h0);
  reg [(3'h4):(1'h0)] reg999 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg992 = (1'h0);
  reg [(4'he):(1'h0)] forvar991 = (1'h0);
  reg [(4'he):(1'h0)] reg996 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar992 = (1'h0);
  reg [(3'h6):(1'h0)] reg990 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar983 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg988 = (1'h0);
  reg [(4'h8):(1'h0)] reg987 = (1'h0);
  reg [(4'h8):(1'h0)] reg985 = (1'h0);
  reg [(5'h17):(1'h0)] reg981 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg980 = (1'h0);
  reg [(3'h6):(1'h0)] reg976 = (1'h0);
  reg [(5'h16):(1'h0)] reg975 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar969 = (1'h0);
  reg [(4'ha):(1'h0)] reg972 = (1'h0);
  reg [(5'h16):(1'h0)] reg971 = (1'h0);
  reg [(5'h14):(1'h0)] reg970 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg969 = (1'h0);
  reg [(5'h13):(1'h0)] reg967 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar962 = (1'h0);
  reg [(5'h13):(1'h0)] reg958 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg956 = (1'h0);
  reg [(4'hb):(1'h0)] reg955 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg954 = (1'h0);
  reg [(5'h13):(1'h0)] reg953 = (1'h0);
  reg [(5'h11):(1'h0)] forvar952 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg950 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg949 = (1'h0);
  reg [(4'he):(1'h0)] reg943 = (1'h0);
  reg [(5'h13):(1'h0)] forvar942 = (1'h0);
  reg [(2'h3):(1'h0)] forvar941 = (1'h0);
  reg [(3'h5):(1'h0)] reg939 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg937 = (1'h0);
  reg [(4'he):(1'h0)] reg936 = (1'h0);
  reg [(5'h13):(1'h0)] reg935 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar932 = (1'h0);
  reg [(5'h10):(1'h0)] forvar931 = (1'h0);
  reg [(4'h9):(1'h0)] reg929 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg928 = (1'h0);
  reg [(3'h4):(1'h0)] forvar925 = (1'h0);
  reg [(3'h5):(1'h0)] reg924 = (1'h0);
  reg [(5'h16):(1'h0)] reg920 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg919 = (1'h0);
  reg signed [(4'he):(1'h0)] reg915 = (1'h0);
  reg [(4'hb):(1'h0)] reg913 = (1'h0);
  reg [(5'h17):(1'h0)] reg912 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar910 = (1'h0);
  reg [(2'h3):(1'h0)] reg909 = (1'h0);
  reg [(5'h14):(1'h0)] forvar908 = (1'h0);
  reg [(5'h10):(1'h0)] reg905 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg904 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg902 = (1'h0);
  reg [(5'h12):(1'h0)] reg900 = (1'h0);
  reg [(5'h14):(1'h0)] reg896 = (1'h0);
  reg [(2'h2):(1'h0)] forvar895 = (1'h0);
  reg [(5'h17):(1'h0)] forvar894 = (1'h0);
  reg [(5'h12):(1'h0)] reg893 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg890 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg889 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg887 = (1'h0);
  reg [(3'h5):(1'h0)] reg884 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar881 = (1'h0);
  reg [(3'h6):(1'h0)] reg880 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg877 = (1'h0);
  reg [(4'he):(1'h0)] reg874 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg873 = (1'h0);
  reg [(5'h17):(1'h0)] reg870 = (1'h0);
  reg [(5'h15):(1'h0)] reg868 = (1'h0);
  reg [(4'he):(1'h0)] reg866 = (1'h0);
  reg [(4'h8):(1'h0)] reg865 = (1'h0);
  assign y = {wire1055,
                 wire1054,
                 wire1053,
                 wire1052,
                 wire1051,
                 wire1043,
                 wire1036,
                 wire1001,
                 wire1000,
                 wire982,
                 wire951,
                 wire863,
                 wire862,
                 reg1045,
                 reg1049,
                 reg1047,
                 reg1038,
                 reg1035,
                 reg1034,
                 reg1031,
                 reg1028,
                 reg1027,
                 reg1025,
                 reg1023,
                 reg1021,
                 reg1016,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1015,
                 reg1014,
                 reg1011,
                 reg1009,
                 reg1006,
                 reg1004,
                 reg998,
                 reg997,
                 reg995,
                 reg994,
                 reg993,
                 reg991,
                 reg989,
                 reg986,
                 reg984,
                 reg983,
                 reg979,
                 reg978,
                 reg977,
                 reg974,
                 reg973,
                 reg968,
                 reg966,
                 reg965,
                 reg964,
                 reg963,
                 reg961,
                 reg960,
                 reg959,
                 reg957,
                 reg948,
                 reg947,
                 reg946,
                 reg945,
                 reg944,
                 reg940,
                 reg938,
                 reg934,
                 reg933,
                 reg930,
                 reg927,
                 reg926,
                 reg923,
                 reg922,
                 reg921,
                 reg918,
                 reg917,
                 reg916,
                 reg914,
                 reg911,
                 reg907,
                 reg906,
                 reg903,
                 reg901,
                 reg899,
                 reg898,
                 reg897,
                 reg892,
                 reg891,
                 reg888,
                 reg886,
                 reg885,
                 reg883,
                 reg882,
                 reg879,
                 reg878,
                 reg876,
                 reg875,
                 reg872,
                 reg871,
                 reg869,
                 reg867,
                 reg864,
                 reg1048,
                 reg1050,
                 forvar1048,
                 reg1046,
                 forvar1045,
                 reg1044,
                 reg1042,
                 reg1041,
                 reg1040,
                 reg1039,
                 reg1037,
                 reg1033,
                 reg1032,
                 reg1030,
                 forvar1029,
                 reg1026,
                 reg1024,
                 reg1022,
                 reg1020,
                 forvar1016,
                 reg1013,
                 reg1012,
                 reg1010,
                 reg1008,
                 reg1007,
                 reg1005,
                 forvar1003,
                 forvar1002,
                 reg999,
                 reg992,
                 forvar991,
                 reg996,
                 forvar992,
                 reg990,
                 forvar983,
                 reg988,
                 reg987,
                 reg985,
                 reg981,
                 reg980,
                 reg976,
                 reg975,
                 forvar969,
                 reg972,
                 reg971,
                 reg970,
                 reg969,
                 reg967,
                 forvar962,
                 reg958,
                 reg956,
                 reg955,
                 reg954,
                 reg953,
                 forvar952,
                 reg950,
                 reg949,
                 reg943,
                 forvar942,
                 forvar941,
                 reg939,
                 reg937,
                 reg936,
                 reg935,
                 forvar932,
                 forvar931,
                 reg929,
                 reg928,
                 forvar925,
                 reg924,
                 reg920,
                 reg919,
                 reg915,
                 reg913,
                 reg912,
                 forvar910,
                 reg909,
                 forvar908,
                 reg905,
                 reg904,
                 reg902,
                 reg900,
                 reg896,
                 forvar895,
                 forvar894,
                 reg893,
                 reg890,
                 reg889,
                 reg887,
                 reg884,
                 forvar881,
                 reg880,
                 reg877,
                 reg874,
                 reg873,
                 reg870,
                 reg868,
                 reg866,
                 reg865,
                 (1'h0)};
  assign wire862 = wire860;
  assign wire863 = $unsigned((^({wire862,
                       $unsigned(wire859)} - $unsigned(wire861))));
  always
    @(posedge clk) begin
      if ((((((wire859 + wire863) ?
                  $unsigned(wire861) : $signed(wire861)) > wire863[(4'ha):(3'h7)]) ?
              $signed(wire861[(4'h9):(3'h5)]) : $signed({wire863})) ?
          {wire859[(2'h3):(2'h2)], wire862} : wire859[(3'h4):(2'h3)]))
        begin
          reg864 <= wire858[(4'he):(4'ha)];
          reg865 = (&wire863);
          if ($unsigned(($signed({((8'h9d) ? (8'hb2) : wire862)}) ?
              (|$signed((8'hb5))) : wire861[(4'he):(1'h0)])))
            begin
              reg866 = wire861[(3'h4):(2'h2)];
              reg867 <= ((reg865 ?
                      (^~$unsigned(reg866[(4'hb):(2'h3)])) : ($unsigned(wire862[(5'h10):(4'hc)]) >>> $unsigned((wire863 << (7'h45))))) ?
                  reg864 : wire859);
              reg868 = $unsigned($unsigned((+reg866)));
              reg869 <= ((~|(~|reg868[(2'h2):(1'h0)])) ?
                  (+$unsigned($signed(wire863))) : (-{reg868[(5'h13):(4'hb)],
                      {$unsigned(wire861)}}));
              reg870 = $unsigned({(reg866 ?
                      $signed(reg864) : $signed(reg868))});
            end
          else
            begin
              reg866 = $signed(reg864);
              reg867 <= (8'ha3);
            end
          if ($unsigned(((((reg864 || reg866) ?
                  {wire863,
                      wire863} : reg867[(1'h0):(1'h0)]) & $signed((!wire860))) ?
              (^(!reg870[(3'h4):(3'h4)])) : $unsigned(($unsigned(reg865) ?
                  reg866[(4'ha):(3'h6)] : $signed(reg865))))))
            begin
              reg871 <= (~&(wire861 > (($signed(wire863) ?
                  $signed(reg865) : reg865) || $unsigned((reg865 * wire858)))));
              reg872 <= $signed(reg866);
            end
          else
            begin
              reg871 <= (&$unsigned($signed(((reg872 * reg872) != wire860))));
            end
        end
      else
        begin
          reg864 <= ($unsigned((^~reg864)) < (reg867 ?
              (~|((reg868 ? reg869 : reg869) ?
                  $signed(reg872) : $signed(reg870))) : ($signed(((8'h9d) && wire861)) ?
                  (~^{reg865, reg871}) : $signed((wire861 ?
                      (8'hb6) : (7'h40))))));
          if (($signed(({((8'haa) ? reg872 : (8'hbb)), $unsigned(reg867)} ?
                  ($unsigned(reg865) ^ wire858[(4'hc):(4'hc)]) : $unsigned((wire859 ?
                      (7'h4a) : wire859)))) ?
              $signed($unsigned({(wire860 ?
                      reg867 : (8'hac))})) : ((((!reg871) ?
                  $signed(reg869) : wire858[(1'h0):(1'h0)]) ~^ ($signed(wire858) ?
                  $unsigned(reg872) : (reg865 - reg866))) && wire862[(2'h2):(2'h2)])))
            begin
              reg865 = $signed(((-((reg868 ?
                  wire860 : (8'hb7)) < reg867)) != ((reg869[(4'hb):(4'hb)] ?
                  (reg871 | reg872) : $unsigned((8'ha2))) == reg865[(2'h2):(1'h0)])));
              reg866 = (^(8'hba));
              reg868 = (reg872 >> reg871[(4'hf):(4'hc)]);
              reg869 <= (~&(((-$unsigned(wire861)) ?
                      reg867 : (wire860 - $unsigned(reg872))) ?
                  (|($signed(reg865) ?
                      $unsigned(reg872) : reg869[(3'h7):(1'h1)])) : $unsigned($unsigned((~^(8'ha0))))));
              reg870 = {reg867[(3'h4):(2'h3)],
                  $signed((wire861 & {(|wire859),
                      ((8'h9c) ? (8'hb9) : reg870)}))};
            end
          else
            begin
              reg865 = (((8'h9e) >= reg865) ?
                  (wire859 << reg865) : {reg865[(2'h3):(2'h3)],
                      (!$signed((wire860 ^ (8'ha5))))});
              reg867 <= (~&(-($unsigned($signed(reg867)) >= (reg872[(1'h0):(1'h0)] ?
                  (+(8'hae)) : (8'ha4)))));
            end
          reg873 = {(~&$signed($signed((reg870 ? reg870 : reg864)))), {reg870}};
          if (({$unsigned((+reg871)),
                  $signed(((wire858 | wire859) ?
                      (-reg864) : (reg866 > reg867)))} ?
              $signed((-{$unsigned(reg871),
                  ((8'had) ? reg870 : reg868)})) : (~&wire861[(1'h1):(1'h0)])))
            begin
              reg874 = (((~^{$unsigned(reg868), reg869}) ?
                      $unsigned((&reg865)) : $signed($unsigned((reg864 ?
                          wire862 : wire862)))) ?
                  $signed(wire863) : $signed(reg872));
              reg875 <= $unsigned($unsigned(reg871[(5'h13):(5'h13)]));
            end
          else
            begin
              reg875 <= $unsigned(reg872[(3'h4):(2'h2)]);
              reg876 <= (~^(~&{$signed((~|reg869))}));
              reg877 = (~&$unsigned(((-$unsigned(wire861)) ?
                  {(~|(8'ha1))} : $signed((reg873 ? wire862 : reg876)))));
              reg878 <= ($unsigned((^~(wire863 != $unsigned((8'hb7))))) == reg866);
            end
          reg879 <= (^~$signed(wire861));
        end
      reg880 = ($unsigned(((-(reg878 <<< reg875)) ~^ ({(8'ha7)} ?
              (~^(8'ha9)) : reg868))) ?
          $signed(reg864[(3'h4):(3'h4)]) : reg870[(5'h15):(3'h5)]);
    end
  always
    @(posedge clk) begin
      for (forvar881 = (1'h0); (forvar881 < (3'h4)); forvar881 = (forvar881 + (1'h1)))
        begin
          if ((^~$unsigned((~^$unsigned((wire863 >> reg871))))))
            begin
              reg882 <= (!$signed($unsigned(((~|reg872) ~^ (^~wire861)))));
              reg883 <= (8'hb4);
            end
          else
            begin
              reg884 = (^~(reg879[(1'h0):(1'h0)] ?
                  reg876[(3'h4):(2'h3)] : reg875));
              reg885 <= {(~^$unsigned($signed((reg867 & reg878))))};
              reg886 <= (+wire862[(4'ha):(4'h8)]);
              reg887 = reg876[(4'ha):(4'h8)];
              reg888 <= $unsigned((reg871[(3'h6):(2'h2)] <= ((wire859 ^ (~^(8'ha3))) ?
                  reg864[(4'hd):(4'h8)] : wire858)));
            end
          reg889 = (-reg869);
          reg890 = (($signed(forvar881) && $signed($signed((!(8'ha6))))) == (+$signed(wire863[(4'ha):(2'h2)])));
          reg891 <= reg886;
        end
    end
  always
    @(posedge clk) begin
      reg892 <= {reg867[(4'h9):(3'h4)]};
      reg893 = $signed({reg883});
      for (forvar894 = (1'h0); (forvar894 < (3'h4)); forvar894 = (forvar894 + (1'h1)))
        begin
          for (forvar895 = (1'h0); (forvar895 < (2'h2)); forvar895 = (forvar895 + (1'h1)))
            begin
              reg896 = {((~$signed((wire860 && forvar895))) ?
                      $signed(reg869) : {$unsigned((reg879 ?
                              (8'hb2) : (8'ha4)))}),
                  ($unsigned($signed((reg864 ?
                      (7'h49) : reg891))) || wire862[(3'h4):(2'h3)])};
              reg897 <= $unsigned((!$signed($unsigned((&reg876)))));
              reg898 <= $signed($unsigned(wire863[(4'hc):(4'h8)]));
              reg899 <= ({wire860} ?
                  (&$signed(((~&reg875) & $unsigned(reg879)))) : (-reg888));
              reg900 = reg882;
            end
          if ($unsigned((({$signed(reg892), reg867[(3'h5):(2'h3)]} ?
                  {$signed((7'h46))} : reg897) ?
              $signed($unsigned(reg875[(5'h10):(1'h1)])) : reg879[(2'h3):(1'h0)])))
            begin
              reg901 <= $signed(($signed(({reg888, forvar894} ?
                      (reg886 ? (8'ha5) : wire859) : (~&reg864))) ?
                  (~|(reg893[(5'h11):(4'hd)] ?
                      (&reg875) : ((7'h46) ?
                          reg864 : reg871))) : reg898[(2'h3):(1'h1)]));
              reg902 = reg891[(3'h4):(3'h4)];
            end
          else
            begin
              reg902 = $signed({wire860,
                  (reg871 == (((7'h43) ? wire858 : reg902) ?
                      ((8'hb9) ? reg900 : reg864) : (8'ha5)))});
            end
          reg903 <= $signed($signed($signed(((wire858 << reg898) ?
              (^reg898) : (reg864 ? reg891 : (8'hba))))));
          if (reg876[(5'h12):(2'h3)])
            begin
              reg904 = {reg897};
              reg905 = (8'hac);
              reg906 <= $unsigned($signed($unsigned((reg888 ?
                  (~reg878) : (reg883 ? reg872 : reg901)))));
            end
          else
            begin
              reg904 = $signed(wire862);
              reg905 = $unsigned($unsigned(((forvar894[(5'h11):(3'h7)] >> reg867[(2'h3):(2'h3)]) >> ($unsigned(wire860) >> $unsigned(forvar895)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg907 <= $signed((reg882 >> wire859[(2'h3):(1'h0)]));
      for (forvar908 = (1'h0); (forvar908 < (1'h1)); forvar908 = (forvar908 + (1'h1)))
        begin
          reg909 = $unsigned(forvar908[(4'hf):(3'h7)]);
          for (forvar910 = (1'h0); (forvar910 < (2'h3)); forvar910 = (forvar910 + (1'h1)))
            begin
              reg911 <= reg882;
              reg912 = wire862;
              reg913 = (&reg903[(1'h0):(1'h0)]);
              reg914 <= $unsigned(reg909);
              reg915 = ({$unsigned((wire858 & (8'ha3))),
                  ($unsigned(wire863[(1'h0):(1'h0)]) >>> ((~^wire861) <= reg891[(2'h2):(1'h0)]))} ^~ $signed((+(wire860[(4'h9):(3'h7)] - (reg911 >> reg871)))));
            end
          reg916 <= reg909[(2'h2):(2'h2)];
          if (wire859)
            begin
              reg917 <= $signed(forvar908);
              reg918 <= $unsigned(reg879[(1'h0):(1'h0)]);
              reg919 = $signed($unsigned(reg918));
              reg920 = (reg915 == (+reg911));
              reg921 <= (!(!{$unsigned({reg907}), (&((8'h9d) * reg918))}));
            end
          else
            begin
              reg919 = ((wire861[(3'h6):(1'h1)] ?
                      (reg916 ^~ (^~(reg916 ?
                          reg878 : reg872))) : reg909[(2'h3):(1'h0)]) ?
                  reg898[(1'h1):(1'h0)] : $signed(reg869));
              reg921 <= (({$unsigned((wire861 ~^ (8'hae))),
                      ($signed(reg879) >= reg876)} ?
                  reg897[(3'h6):(1'h1)] : (~&$unsigned($signed((8'had))))) * reg891[(3'h5):(1'h1)]);
              reg922 <= reg872[(4'h8):(3'h6)];
              reg923 <= $signed((reg922[(2'h2):(1'h0)] ?
                  ((~&reg897) ?
                      reg892 : ((!reg883) ?
                          (8'ha3) : wire861[(1'h0):(1'h0)])) : $unsigned($unsigned((reg897 & (8'hae))))));
              reg924 = wire862[(4'hd):(3'h6)];
            end
          for (forvar925 = (1'h0); (forvar925 < (2'h3)); forvar925 = (forvar925 + (1'h1)))
            begin
              reg926 <= wire861[(3'h4):(3'h4)];
              reg927 <= (($unsigned(((~&forvar908) ?
                  {reg911,
                      reg883} : reg924[(1'h1):(1'h0)])) * $unsigned({reg891[(3'h7):(2'h2)]})) != (+(forvar925[(1'h0):(1'h0)] ?
                  $unsigned((wire863 ? (7'h41) : reg882)) : reg915)));
              reg928 = {(&(reg869[(3'h4):(3'h4)] ~^ reg888[(2'h3):(2'h2)]))};
              reg929 = $signed(((($unsigned(reg903) ?
                  (forvar908 ?
                      reg886 : reg920) : reg875[(4'hf):(1'h1)]) * ($signed(reg921) | $signed(reg907))) || reg882[(2'h3):(2'h3)]));
              reg930 <= reg928;
            end
        end
      for (forvar931 = (1'h0); (forvar931 < (2'h3)); forvar931 = (forvar931 + (1'h1)))
        begin
          for (forvar932 = (1'h0); (forvar932 < (2'h2)); forvar932 = (forvar932 + (1'h1)))
            begin
              reg933 <= (+((~^reg917[(3'h4):(3'h4)]) <<< reg920[(3'h5):(1'h0)]));
              reg934 <= (-{$unsigned($unsigned((reg917 ? (8'had) : (7'h49))))});
              reg935 = (-forvar910);
            end
          reg936 = (reg906[(4'hc):(3'h5)] ?
              (((+((7'h41) - reg924)) ?
                      reg888[(2'h3):(1'h1)] : $signed($unsigned(reg867))) ?
                  reg897[(3'h5):(2'h3)] : ({{(8'h9c)}} ?
                      ($signed(reg934) ?
                          $unsigned(reg875) : $signed(reg923)) : ((+reg871) ?
                          reg922[(1'h0):(1'h0)] : forvar931))) : $unsigned({reg916,
                  wire862}));
          if ($signed($unsigned($signed(($signed(reg913) ?
              $unsigned(reg914) : reg876[(4'hc):(3'h7)])))))
            begin
              reg937 = reg875[(3'h4):(3'h4)];
            end
          else
            begin
              reg938 <= reg867[(3'h4):(3'h4)];
              reg939 = (reg888 < (~reg935[(5'h13):(2'h2)]));
            end
          reg940 <= ((forvar910[(5'h10):(3'h5)] ?
              $signed((reg928[(2'h3):(1'h0)] ?
                  reg879[(3'h4):(3'h4)] : ((8'hbe) <= reg885))) : reg888) & reg914);
        end
      for (forvar941 = (1'h0); (forvar941 < (3'h4)); forvar941 = (forvar941 + (1'h1)))
        begin
          for (forvar942 = (1'h0); (forvar942 < (2'h3)); forvar942 = (forvar942 + (1'h1)))
            begin
              reg943 = $unsigned($signed((reg909[(2'h3):(2'h3)] + $signed($signed(reg916)))));
            end
          reg944 <= reg886;
          reg945 <= $signed(reg892);
          if (reg888[(2'h3):(2'h2)])
            begin
              reg946 <= $signed($unsigned($unsigned((^(reg883 <= (7'h40))))));
              reg947 <= {$unsigned((reg917[(3'h4):(3'h4)] <<< (~|$signed(reg897))))};
              reg948 <= ((reg913[(2'h3):(1'h0)] ?
                  $signed({reg869, {reg885}}) : (forvar942[(2'h3):(1'h0)] ?
                      wire860 : $signed(((8'ha4) ?
                          (8'h9e) : reg906)))) >>> $signed(reg916));
            end
          else
            begin
              reg946 <= ($unsigned(($signed((reg906 ?
                      reg934 : reg911)) >> {{(8'ha3)}, $signed(reg933)})) ?
                  reg943 : ((~&{$signed(reg936)}) ~^ ($unsigned($signed(reg919)) ^ (^~(-reg864)))));
              reg947 <= reg922[(3'h7):(3'h7)];
              reg948 <= (!({reg913,
                      ((reg934 ? reg916 : (7'h46)) != (reg912 ^ reg885))} ?
                  reg869 : ((reg899[(3'h6):(1'h1)] || $unsigned(reg879)) ?
                      (~&$unsigned(reg907)) : $signed(((8'hac) == reg883)))));
              reg949 = reg918[(4'hc):(4'hc)];
            end
        end
      reg950 = $unsigned($signed((forvar942[(4'h9):(2'h3)] - ($unsigned(wire858) ?
          (forvar925 ? reg918 : (8'h9d)) : reg886[(4'h9):(3'h6)]))));
    end
  assign wire951 = reg930[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar952 = (1'h0); (forvar952 < (2'h3)); forvar952 = (forvar952 + (1'h1)))
        begin
          if ($signed($signed(((((7'h40) ? reg947 : (8'h9e)) ?
              $unsigned(forvar952) : wire951) | ((-(8'ha8)) + {reg892})))))
            begin
              reg953 = ((reg898 >>> (^$unsigned(reg911))) ?
                  {$unsigned(({wire951} || (!reg875)))} : reg930[(1'h0):(1'h0)]);
              reg954 = $signed(reg903[(4'hb):(4'h8)]);
              reg955 = $unsigned($signed((7'h49)));
              reg956 = $unsigned({reg938[(5'h13):(4'h9)]});
            end
          else
            begin
              reg957 <= $signed(($signed(reg940) ?
                  reg914 : {((8'ha9) * $unsigned(reg914)),
                      $unsigned((reg954 ^ reg897))}));
              reg958 = ((^~(+(reg869 ? ((8'h9d) > wire951) : (8'hbe)))) ?
                  $signed((reg955 >>> $unsigned(wire863))) : $signed(($unsigned($signed(reg883)) ?
                      $signed((reg867 < reg930)) : (+reg872[(2'h3):(1'h0)]))));
              reg959 <= {$signed((~((wire951 != (8'ha6)) == wire861[(4'hd):(4'ha)]))),
                  ($unsigned(((reg867 ?
                      reg867 : (8'ha6)) > (7'h49))) & $signed(reg934[(1'h0):(1'h0)]))};
              reg960 <= {({((wire860 < reg933) ?
                          $signed(reg879) : reg944)} || $unsigned(((reg891 <<< reg882) & $unsigned(reg934))))};
              reg961 <= {$unsigned(($signed((8'haf)) ?
                      reg922 : ((reg878 ? reg955 : reg869) ?
                          (reg960 ^~ reg907) : $signed(reg879)))),
                  ($unsigned((~&reg892[(3'h4):(1'h1)])) ?
                      (!{{reg886}}) : (-reg888))};
            end
          for (forvar962 = (1'h0); (forvar962 < (1'h0)); forvar962 = (forvar962 + (1'h1)))
            begin
              reg963 <= $signed(reg959[(2'h2):(1'h0)]);
              reg964 <= reg867[(1'h0):(1'h0)];
              reg965 <= $unsigned(forvar952);
              reg966 <= $signed({reg958[(1'h1):(1'h0)], reg883[(2'h3):(1'h1)]});
            end
        end
      reg967 = $unsigned(reg879[(2'h2):(2'h2)]);
      reg968 <= $signed(reg921[(1'h1):(1'h1)]);
      if (((~^((^~(reg960 ? reg954 : reg946)) + wire859[(3'h6):(1'h1)])) ?
          reg872[(3'h6):(3'h4)] : $unsigned($signed(reg961[(4'h8):(3'h7)]))))
        begin
          if ((({(reg930 ?
                      {reg957,
                          reg923} : reg906[(2'h3):(1'h1)])} <= $signed(({reg938} ?
                  wire858[(5'h13):(5'h13)] : $signed(reg911)))) ?
              reg922[(3'h6):(1'h1)] : $unsigned($unsigned($unsigned((reg883 ?
                  reg965 : reg882))))))
            begin
              reg969 = (reg933 != $unsigned(((~|(~&forvar962)) <= reg916)));
              reg970 = reg969[(2'h2):(1'h0)];
              reg971 = (-reg970[(4'h8):(2'h2)]);
              reg972 = wire859;
            end
          else
            begin
              reg969 = ({reg965[(2'h3):(1'h1)]} ?
                  {{(~|$unsigned(wire860)),
                          {(reg926 >>> reg914)}}} : ($signed(wire859[(2'h2):(2'h2)]) ?
                      {reg888[(3'h5):(3'h4)]} : $unsigned({$signed(reg944),
                          {reg885}})));
            end
          reg973 <= (|(|($signed((~&reg885)) ?
              ((reg901 ?
                  reg879 : reg882) ^ (reg927 >= reg885)) : (forvar962[(4'ha):(4'h9)] + $unsigned(reg947)))));
        end
      else
        begin
          for (forvar969 = (1'h0); (forvar969 < (3'h4)); forvar969 = (forvar969 + (1'h1)))
            begin
              reg970 = reg948;
              reg973 <= ($unsigned($unsigned(($signed(reg879) ^ reg955[(1'h1):(1'h1)]))) ?
                  (8'ha3) : $signed({(+$unsigned((8'hbd)))}));
              reg974 <= reg958;
              reg975 = forvar969;
            end
          reg976 = $unsigned(reg872[(3'h4):(2'h3)]);
        end
      reg977 <= reg867;
    end
  always
    @(posedge clk) begin
      reg978 <= (($unsigned((~&(reg960 << reg968))) ?
              (-$unsigned((^~reg922))) : ({{(8'ha6)}} ?
                  ((reg938 ? reg940 : reg922) ?
                      $signed(reg948) : $unsigned((8'hab))) : $signed($unsigned((8'h9f))))) ?
          ($signed($signed({(8'hac),
              reg898})) != reg938[(4'he):(2'h3)]) : $signed((((reg964 || reg947) ?
              reg886 : (reg966 > reg876)) == $signed(reg921[(3'h5):(3'h4)]))));
      reg979 <= reg926[(5'h10):(4'hd)];
      reg980 = ($signed(((+(reg871 - reg875)) ?
          reg963[(3'h6):(1'h0)] : {(reg978 ? (8'hb9) : reg914),
              (~|reg968)})) << $signed({($unsigned((8'ha7)) - (~&(8'hb6))),
          reg948[(4'hc):(4'h8)]}));
      reg981 = (-wire951);
    end
  assign wire982 = $unsigned(reg876[(3'h7):(3'h6)]);
  always
    @(posedge clk) begin
      if ((reg947 | ((reg957[(1'h0):(1'h0)] ? $signed(reg926) : {(|reg871)}) ?
          reg882 : (wire858 >> ((reg888 | reg885) ?
              reg916 : $signed(wire859))))))
        begin
          if (reg879[(2'h3):(2'h3)])
            begin
              reg983 <= reg979[(4'h9):(1'h0)];
              reg984 <= $signed(wire982);
              reg985 = reg891[(4'hc):(2'h3)];
              reg986 <= ($signed(reg897[(3'h5):(2'h2)]) >>> {reg871});
            end
          else
            begin
              reg983 <= (~&$unsigned(((^$unsigned(wire860)) ?
                  (reg974 ^~ ((8'hba) ?
                      (8'ha8) : reg973)) : $unsigned(reg965[(4'ha):(4'h9)]))));
              reg985 = reg876[(4'hc):(3'h5)];
              reg986 <= (!((wire861 <= $signed({reg907})) ?
                  (($unsigned((8'hb5)) >> reg882[(3'h5):(1'h1)]) ?
                      {$unsigned(reg906)} : wire863) : wire951));
              reg987 = (~|(~reg876));
            end
          reg988 = reg984;
        end
      else
        begin
          for (forvar983 = (1'h0); (forvar983 < (2'h2)); forvar983 = (forvar983 + (1'h1)))
            begin
              reg985 = {$signed({$unsigned(reg930), $unsigned({reg944})}),
                  (+({(wire863 ? reg960 : reg891)} ^ ((wire860 || reg882) ?
                      {reg977} : $signed(reg899))))};
              reg987 = forvar983[(3'h5):(1'h0)];
              reg989 <= (!(+(^({wire858} ?
                  $unsigned(reg901) : (reg957 >> reg917)))));
              reg990 = $signed((reg973 ?
                  (((reg944 & reg938) ?
                      reg911[(4'ha):(2'h3)] : reg918[(4'hb):(2'h2)]) && $unsigned((^~(8'hb0)))) : $unsigned(((^~reg966) ?
                      $unsigned((8'hb2)) : (reg978 ? reg879 : reg968)))));
            end
        end
      if ((^reg922[(2'h2):(2'h2)]))
        begin
          reg991 <= ({(^$unsigned((^~reg968))),
              ($signed($unsigned(reg990)) ?
                  (~$signed((7'h49))) : (reg869[(3'h5):(1'h1)] ?
                      {reg959,
                          (8'hbe)} : $unsigned(reg891)))} & $signed(reg901[(3'h7):(1'h0)]));
          for (forvar992 = (1'h0); (forvar992 < (3'h4)); forvar992 = (forvar992 + (1'h1)))
            begin
              reg993 <= $unsigned(reg933);
              reg994 <= ($signed(reg933) ?
                  ((reg940[(2'h2):(1'h1)] ?
                          ($signed(wire863) ^ (^reg916)) : (reg945 ?
                              (reg963 > reg918) : (~wire861))) ?
                      $unsigned(reg977[(2'h3):(2'h2)]) : {({reg989} ?
                              ((8'hbd) << reg879) : (reg878 << reg892))}) : ($unsigned(reg987) + (-((reg965 <= wire859) ?
                      reg960[(4'h8):(3'h4)] : (reg946 ? reg886 : reg944)))));
              reg995 <= reg979[(4'hc):(3'h7)];
              reg996 = (reg959[(2'h2):(2'h2)] ?
                  (({(reg966 ?
                          reg899 : wire859)} + $signed($signed(wire861))) | (reg974 ?
                      $signed((8'h9f)) : (|$unsigned(reg891)))) : (&reg875));
              reg997 <= (|{$signed($unsigned(reg983))});
            end
        end
      else
        begin
          for (forvar991 = (1'h0); (forvar991 < (1'h1)); forvar991 = (forvar991 + (1'h1)))
            begin
              reg992 = (((^(((8'hb5) ? wire860 : (8'hbd)) ?
                  $unsigned(reg964) : forvar992)) - reg879) >= (({$unsigned(reg940),
                      $signed(reg984)} != ((+reg907) > (wire858 ~^ reg906))) ?
                  reg930 : wire861[(4'hd):(1'h1)]));
            end
          reg993 <= reg991;
        end
      reg998 <= (^~reg864[(1'h0):(1'h0)]);
      reg999 = $unsigned($unsigned(($signed({wire863}) >> (reg986[(4'h8):(4'h8)] ?
          (reg875 ? reg879 : reg923) : ((7'h42) || (8'ha3))))));
    end
  assign wire1000 = $unsigned((^~(&reg923)));
  assign wire1001 = $unsigned(reg882[(4'hb):(3'h5)]);
  always
    @(posedge clk) begin
      for (forvar1002 = (1'h0); (forvar1002 < (2'h2)); forvar1002 = (forvar1002 + (1'h1)))
        begin
          for (forvar1003 = (1'h0); (forvar1003 < (3'h4)); forvar1003 = (forvar1003 + (1'h1)))
            begin
              reg1004 <= reg938;
              reg1005 = ((reg978 - (|$signed((reg923 ? reg906 : reg901)))) ?
                  (reg871 ?
                      ({(reg979 & reg959)} <= ($signed(reg922) ?
                          wire863 : {(8'ha8),
                              reg892})) : wire861) : ((reg892 < (reg901 ?
                          (+reg965) : (reg998 > wire858))) ?
                      reg991[(3'h6):(3'h6)] : (~|(~(reg879 ?
                          reg921 : reg903)))));
              reg1006 <= {$signed((forvar1002 >= $signed(reg960[(5'h10):(1'h1)])))};
            end
          if ($signed((+reg938)))
            begin
              reg1007 = reg945[(1'h0):(1'h0)];
              reg1008 = $unsigned(reg945[(2'h2):(1'h0)]);
              reg1009 <= ((|reg989[(2'h2):(2'h2)]) ?
                  reg948 : $unsigned(reg885[(4'he):(1'h1)]));
            end
          else
            begin
              reg1009 <= (reg977[(2'h3):(2'h3)] ?
                  ($unsigned($unsigned((-reg991))) ~^ (^{$unsigned(reg1008),
                      (reg918 ? reg901 : forvar1002)})) : (!reg974));
              reg1010 = {($unsigned({$unsigned(reg945),
                          reg979[(3'h5):(1'h1)]}) ?
                      (((reg1006 ? reg977 : reg892) ?
                          (reg991 > reg885) : reg891) & $unsigned($unsigned(reg879))) : {(reg886 + $unsigned(reg871)),
                          {$unsigned((8'haa)), $unsigned(forvar1002)}})};
              reg1011 <= ($signed(reg864) ?
                  reg927[(2'h2):(2'h2)] : reg989[(3'h4):(1'h1)]);
              reg1012 = (!reg983);
              reg1013 = reg875;
            end
        end
      if ((reg883 < reg991[(4'hd):(4'h8)]))
        begin
          reg1014 <= {(^~reg940[(2'h3):(2'h2)])};
          reg1015 <= reg998[(5'h10):(4'hd)];
          for (forvar1016 = (1'h0); (forvar1016 < (3'h4)); forvar1016 = (forvar1016 + (1'h1)))
            begin
              reg1017 <= reg977[(2'h3):(2'h3)];
              reg1018 <= $signed(wire861[(1'h1):(1'h0)]);
              reg1019 <= $signed($unsigned((-reg1017)));
            end
          reg1020 = (~&$signed(($signed($unsigned(reg922)) || (8'hb5))));
        end
      else
        begin
          reg1014 <= (((reg960[(2'h3):(2'h3)] ?
                  reg886 : $unsigned(((8'ha5) ?
                      reg1015 : (7'h47)))) == $signed((^~((8'hba) ^~ (7'h46))))) ?
              (~^$unsigned(reg961)) : (($signed({reg979,
                  reg918}) >= reg978[(4'ha):(4'h8)]) && $signed(((reg867 ?
                  reg898 : (7'h43)) == {reg995}))));
          reg1015 <= ((reg921 + (-$signed({reg940, reg986}))) <<< (reg963 ?
              $unsigned($signed({reg964,
                  reg869})) : ($signed((reg995 != reg998)) ?
                  $signed($signed(reg963)) : reg933)));
          if (reg891[(4'hc):(1'h0)])
            begin
              reg1016 <= {{$unsigned(reg986[(2'h3):(2'h2)]),
                      (((!reg914) ? ((8'hab) * wire1000) : $unsigned(reg984)) ?
                          $signed($unsigned(wire859)) : (reg933 >> (reg946 >>> reg1007)))},
                  reg883[(1'h1):(1'h1)]};
              reg1020 = reg899;
              reg1021 <= ((8'hae) ? ((8'hb3) >> reg986) : (~&reg1017));
              reg1022 = $signed(($unsigned((^~$unsigned((8'hae)))) >= reg926[(4'ha):(1'h0)]));
              reg1023 <= $signed((!reg998[(3'h5):(2'h3)]));
            end
          else
            begin
              reg1020 = (!(reg966[(1'h0):(1'h0)] <<< $signed($signed($unsigned(wire858)))));
            end
          if ((($unsigned({reg998[(4'hc):(4'h9)]}) ?
              reg998 : $unsigned({reg948, (7'h47)})) - reg1012[(1'h1):(1'h1)]))
            begin
              reg1024 = reg977;
              reg1025 <= wire1000;
              reg1026 = reg946[(1'h0):(1'h0)];
              reg1027 <= (!(-{$unsigned($unsigned(reg1014))}));
            end
          else
            begin
              reg1025 <= (8'ha5);
              reg1027 <= ($signed({{(reg885 & wire1001), reg926},
                  $signed(reg1007)}) ~^ {{reg1006}, (^(!$signed(reg938)))});
              reg1028 <= (reg891 ?
                  {(&reg882[(4'hb):(4'h8)])} : {(reg1026[(2'h3):(2'h2)] ?
                          $signed((~&reg903)) : ((8'ha2) >> reg886))});
            end
          for (forvar1029 = (1'h0); (forvar1029 < (1'h0)); forvar1029 = (forvar1029 + (1'h1)))
            begin
              reg1030 = reg984;
              reg1031 <= (-(reg886[(5'h18):(3'h4)] > {(((8'hb3) ?
                          reg875 : reg994) ?
                      (reg968 ^~ reg993) : (reg1020 != reg872)),
                  reg917[(4'h9):(3'h7)]}));
              reg1032 = (reg940 - $unsigned(((reg911 ?
                  $unsigned(reg869) : ((8'h9d) << wire863)) <= reg968)));
            end
        end
      reg1033 = $signed(forvar1003[(3'h6):(1'h0)]);
      reg1034 <= (~|$unsigned((((wire1001 | forvar1016) ?
              (reg911 << (8'hb8)) : reg1004) ?
          $unsigned((!reg946)) : {(8'hb9)})));
      reg1035 <= (-($signed((wire951[(3'h7):(2'h3)] ?
              $unsigned(reg978) : (reg964 || reg933))) ?
          reg948[(5'h14):(4'h8)] : reg1011));
    end
  assign wire1036 = (&{{reg1009, $unsigned(wire859)},
                        {((~wire863) & $unsigned(reg957)),
                            reg938[(2'h2):(2'h2)]}});
  always
    @(posedge clk) begin
      reg1037 = $signed($signed(reg961[(2'h2):(2'h2)]));
      reg1038 <= ((reg916 >> ($signed((~^reg968)) ?
              ((reg968 ? reg973 : reg914) ?
                  {reg961} : {reg926}) : reg892[(3'h6):(1'h0)])) ?
          (&$unsigned(reg948)) : ($unsigned((reg918 || reg891)) != {$unsigned($unsigned(reg1017)),
              (8'hbb)}));
      reg1039 = ((+reg947[(3'h6):(3'h5)]) ?
          ($unsigned($signed(reg871[(5'h11):(4'hf)])) ?
              $unsigned(($unsigned(reg1027) ?
                  $unsigned(wire862) : $unsigned(wire863))) : wire1036) : wire951);
    end
  always
    @(posedge clk) begin
      reg1040 = {reg978[(3'h5):(1'h0)],
          ($unsigned($unsigned($signed(reg933))) + $unsigned(wire860))};
      reg1041 = wire982[(1'h1):(1'h0)];
      reg1042 = $signed((reg871[(5'h10):(1'h1)] ?
          $signed(reg973[(4'he):(4'he)]) : wire982));
    end
  assign wire1043 = (^(+reg933));
  always
    @(posedge clk) begin
      if ((7'h44))
        begin
          reg1044 = (reg1019[(4'h8):(4'h8)] ?
              reg965[(4'ha):(3'h5)] : (^~reg979[(3'h5):(2'h2)]));
          for (forvar1045 = (1'h0); (forvar1045 < (1'h0)); forvar1045 = (forvar1045 + (1'h1)))
            begin
              reg1046 = ((~|$unsigned(reg960)) + ($unsigned((reg906[(4'ha):(4'h9)] ?
                  reg933[(1'h0):(1'h0)] : $unsigned((8'ha3)))) >> $signed({(^~(8'ha0))})));
              reg1047 <= $unsigned(($signed($unsigned(forvar1045)) != $unsigned((wire858 < reg906))));
            end
          for (forvar1048 = (1'h0); (forvar1048 < (1'h0)); forvar1048 = (forvar1048 + (1'h1)))
            begin
              reg1049 <= reg944;
            end
          reg1050 = reg1021;
        end
      else
        begin
          reg1045 <= (forvar1048[(5'h18):(4'hf)] ~^ reg926[(1'h1):(1'h1)]);
          if (($unsigned(reg968[(4'hd):(4'h9)]) - $unsigned((($unsigned((8'had)) ?
              {reg901, reg959} : (~reg1046)) & $unsigned((reg891 ?
              (8'had) : (8'haa)))))))
            begin
              reg1047 <= {((8'hb5) ^ (~|(-(reg979 ? (7'h40) : (8'hb0)))))};
              reg1048 = (reg940 == $signed($unsigned($signed($unsigned(reg991)))));
            end
          else
            begin
              reg1046 = $unsigned($signed((reg945 >= reg903[(2'h3):(2'h3)])));
            end
        end
    end
  assign wire1051 = $signed(reg926[(4'hf):(3'h4)]);
  assign wire1052 = reg957;
  assign wire1053 = (((~^$signed($signed(wire1043))) <= $signed($unsigned(reg986))) ^ ($unsigned($unsigned({(7'h48),
                            reg930})) ?
                        reg986 : $unsigned((~(reg938 ? (7'h48) : reg964)))));
  assign wire1054 = $signed(reg891);
  assign wire1055 = reg984[(3'h6):(3'h6)];
endmodule