(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param765 = (^~(!(~^(~&(8'hab))))))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h7b8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire0;
  input wire signed [(5'h14):(1'h0)] wire1;
  input wire signed [(5'h11):(1'h0)] wire2;
  input wire signed [(5'h11):(1'h0)] wire3;
  wire signed [(4'h8):(1'h0)] wire764;
  wire signed [(4'h9):(1'h0)] wire708;
  wire signed [(5'h12):(1'h0)] wire707;
  wire signed [(4'h8):(1'h0)] wire706;
  wire [(4'h9):(1'h0)] wire705;
  wire signed [(5'h10):(1'h0)] wire704;
  wire signed [(4'ha):(1'h0)] wire653;
  wire signed [(3'h7):(1'h0)] wire618;
  wire signed [(5'h12):(1'h0)] wire17;
  wire [(4'hc):(1'h0)] wire356;
  wire [(4'hf):(1'h0)] wire616;
  reg signed [(4'h8):(1'h0)] reg763 = (1'h0);
  reg [(5'h14):(1'h0)] reg758 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg757 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg754 = (1'h0);
  reg [(4'hf):(1'h0)] reg753 = (1'h0);
  reg [(2'h3):(1'h0)] reg751 = (1'h0);
  reg [(2'h2):(1'h0)] reg750 = (1'h0);
  reg [(3'h7):(1'h0)] reg749 = (1'h0);
  reg [(3'h6):(1'h0)] reg748 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg747 = (1'h0);
  reg [(4'hc):(1'h0)] reg745 = (1'h0);
  reg [(5'h15):(1'h0)] reg744 = (1'h0);
  reg [(4'h9):(1'h0)] reg742 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg741 = (1'h0);
  reg [(5'h11):(1'h0)] reg739 = (1'h0);
  reg signed [(4'he):(1'h0)] reg738 = (1'h0);
  reg [(4'hb):(1'h0)] reg737 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg736 = (1'h0);
  reg [(5'h14):(1'h0)] reg734 = (1'h0);
  reg [(4'hc):(1'h0)] reg732 = (1'h0);
  reg [(5'h14):(1'h0)] reg729 = (1'h0);
  reg [(4'hf):(1'h0)] reg726 = (1'h0);
  reg [(5'h11):(1'h0)] reg725 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg722 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg721 = (1'h0);
  reg [(5'h11):(1'h0)] reg718 = (1'h0);
  reg [(5'h10):(1'h0)] reg717 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg713 = (1'h0);
  reg [(4'ha):(1'h0)] reg712 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg711 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg710 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg703 = (1'h0);
  reg [(4'he):(1'h0)] reg702 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg701 = (1'h0);
  reg signed [(4'he):(1'h0)] reg699 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg697 = (1'h0);
  reg [(3'h4):(1'h0)] reg696 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg694 = (1'h0);
  reg [(5'h13):(1'h0)] reg691 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg689 = (1'h0);
  reg [(4'h8):(1'h0)] reg684 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg681 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg679 = (1'h0);
  reg [(5'h12):(1'h0)] reg678 = (1'h0);
  reg [(4'hf):(1'h0)] reg677 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg673 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg672 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg670 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg669 = (1'h0);
  reg [(4'hd):(1'h0)] reg668 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg666 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg663 = (1'h0);
  reg [(5'h12):(1'h0)] reg661 = (1'h0);
  reg [(5'h15):(1'h0)] reg659 = (1'h0);
  reg [(5'h15):(1'h0)] reg656 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg655 = (1'h0);
  reg [(4'hb):(1'h0)] reg654 = (1'h0);
  reg [(4'hd):(1'h0)] reg652 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg650 = (1'h0);
  reg [(5'h11):(1'h0)] reg648 = (1'h0);
  reg [(5'h15):(1'h0)] reg646 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg643 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg642 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg636 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg634 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg633 = (1'h0);
  reg [(5'h10):(1'h0)] reg622 = (1'h0);
  reg [(3'h7):(1'h0)] reg631 = (1'h0);
  reg [(4'ha):(1'h0)] reg630 = (1'h0);
  reg [(2'h2):(1'h0)] reg629 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg627 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg621 = (1'h0);
  reg [(5'h12):(1'h0)] reg619 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar762 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg759 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg761 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg760 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar759 = (1'h0);
  reg signed [(4'he):(1'h0)] reg756 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg755 = (1'h0);
  reg [(5'h14):(1'h0)] reg752 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg746 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg743 = (1'h0);
  reg signed [(4'he):(1'h0)] reg740 = (1'h0);
  reg signed [(4'he):(1'h0)] reg735 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar733 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg730 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar728 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar727 = (1'h0);
  reg [(4'h9):(1'h0)] reg724 = (1'h0);
  reg [(3'h5):(1'h0)] forvar723 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg720 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg719 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar716 = (1'h0);
  reg [(5'h13):(1'h0)] reg715 = (1'h0);
  reg [(5'h12):(1'h0)] reg714 = (1'h0);
  reg [(4'h8):(1'h0)] forvar709 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg700 = (1'h0);
  reg [(4'h9):(1'h0)] reg698 = (1'h0);
  reg [(2'h2):(1'h0)] reg692 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg695 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg693 = (1'h0);
  reg [(4'h9):(1'h0)] forvar692 = (1'h0);
  reg [(5'h13):(1'h0)] reg690 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg688 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg687 = (1'h0);
  reg [(4'ha):(1'h0)] reg686 = (1'h0);
  reg [(5'h14):(1'h0)] reg685 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg683 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg682 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg680 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar673 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg676 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg675 = (1'h0);
  reg [(5'h12):(1'h0)] reg674 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg671 = (1'h0);
  reg [(5'h13):(1'h0)] reg667 = (1'h0);
  reg [(4'hd):(1'h0)] reg665 = (1'h0);
  reg [(3'h4):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg662 = (1'h0);
  reg [(2'h3):(1'h0)] forvar654 = (1'h0);
  reg signed [(4'he):(1'h0)] reg660 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg658 = (1'h0);
  reg [(4'ha):(1'h0)] reg657 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg651 = (1'h0);
  reg [(5'h14):(1'h0)] reg649 = (1'h0);
  reg [(5'h10):(1'h0)] forvar647 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg645 = (1'h0);
  reg [(4'hc):(1'h0)] forvar644 = (1'h0);
  reg [(4'hc):(1'h0)] reg641 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg640 = (1'h0);
  reg [(5'h12):(1'h0)] reg639 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg637 = (1'h0);
  reg [(4'hd):(1'h0)] reg635 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar632 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg624 = (1'h0);
  reg [(4'h9):(1'h0)] forvar620 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg628 = (1'h0);
  reg signed [(4'he):(1'h0)] reg626 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg625 = (1'h0);
  reg [(4'hd):(1'h0)] forvar624 = (1'h0);
  reg [(4'hd):(1'h0)] forvar622 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg620 = (1'h0);
  assign y = {wire764,
                 wire708,
                 wire707,
                 wire706,
                 wire705,
                 wire704,
                 wire653,
                 wire618,
                 wire17,
                 wire356,
                 wire616,
                 reg763,
                 reg758,
                 reg757,
                 reg754,
                 reg753,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg747,
                 reg745,
                 reg744,
                 reg742,
                 reg741,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg734,
                 reg732,
                 reg729,
                 reg726,
                 reg725,
                 reg722,
                 reg721,
                 reg718,
                 reg717,
                 reg713,
                 reg712,
                 reg711,
                 reg710,
                 reg703,
                 reg702,
                 reg701,
                 reg699,
                 reg697,
                 reg696,
                 reg694,
                 reg691,
                 reg689,
                 reg684,
                 reg681,
                 reg679,
                 reg678,
                 reg677,
                 reg673,
                 reg672,
                 reg670,
                 reg669,
                 reg668,
                 reg666,
                 reg663,
                 reg661,
                 reg659,
                 reg656,
                 reg655,
                 reg654,
                 reg652,
                 reg650,
                 reg648,
                 reg646,
                 reg643,
                 reg642,
                 reg638,
                 reg636,
                 reg634,
                 reg633,
                 reg622,
                 reg631,
                 reg630,
                 reg629,
                 reg627,
                 reg623,
                 reg621,
                 reg619,
                 forvar762,
                 reg759,
                 reg761,
                 reg760,
                 forvar759,
                 reg756,
                 reg755,
                 reg752,
                 reg746,
                 reg743,
                 reg740,
                 reg735,
                 forvar733,
                 reg731,
                 reg730,
                 forvar728,
                 forvar727,
                 reg724,
                 forvar723,
                 reg720,
                 reg719,
                 forvar716,
                 reg715,
                 reg714,
                 forvar709,
                 reg700,
                 reg698,
                 reg692,
                 reg695,
                 reg693,
                 forvar692,
                 reg690,
                 reg688,
                 reg687,
                 reg686,
                 reg685,
                 reg683,
                 reg682,
                 reg680,
                 forvar673,
                 reg676,
                 reg675,
                 reg674,
                 reg671,
                 reg667,
                 reg665,
                 reg664,
                 reg662,
                 forvar654,
                 reg660,
                 reg658,
                 reg657,
                 reg651,
                 reg649,
                 forvar647,
                 reg645,
                 forvar644,
                 reg641,
                 reg640,
                 reg639,
                 reg637,
                 reg635,
                 forvar632,
                 reg624,
                 forvar620,
                 reg628,
                 reg626,
                 reg625,
                 forvar624,
                 forvar622,
                 reg620,
                 (1'h0)};
  module4 #() modinst18 (wire17, clk, wire0, wire2, wire3, wire1, (8'hac));
  module19 #() modinst357 (wire356, clk, wire0, wire1, wire3, wire17);
  module358 #() modinst617 (wire616, clk, wire1, wire2, wire0, wire356, wire17);
  assign wire618 = wire616[(4'hd):(4'h8)];
  always
    @(posedge clk) begin
      reg619 <= (wire2[(2'h3):(1'h0)] >> (^wire2[(1'h0):(1'h0)]));
      if ((wire616[(3'h5):(3'h4)] <= {((|wire616[(4'hd):(4'hd)]) && (((8'ha3) >= wire1) + (|(8'ha4)))),
          wire616}))
        begin
          reg620 = $unsigned((^~(wire618[(3'h7):(1'h1)] == (((8'hbd) ?
                  wire616 : (8'hb5)) ?
              $signed(wire0) : $signed(wire356)))));
          reg621 <= {$signed(wire3[(3'h6):(2'h2)])};
          for (forvar622 = (1'h0); (forvar622 < (2'h2)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 <= wire17[(4'hf):(4'hf)];
            end
          for (forvar624 = (1'h0); (forvar624 < (2'h2)); forvar624 = (forvar624 + (1'h1)))
            begin
              reg625 = forvar624[(4'ha):(2'h2)];
              reg626 = $signed((&$unsigned($signed($unsigned(wire356)))));
              reg627 <= (8'ha6);
              reg628 = (~|((^wire616) << $unsigned(((reg627 - wire616) >> wire356[(3'h4):(1'h0)]))));
              reg629 <= (reg620[(2'h3):(2'h3)] ~^ $unsigned(reg626[(2'h2):(1'h1)]));
            end
          if ((8'h9c))
            begin
              reg630 <= reg628[(2'h2):(1'h1)];
              reg631 <= $signed(($unsigned($signed(reg619)) < wire616));
            end
          else
            begin
              reg630 <= (((^~reg627) ?
                      (reg619 & (wire2[(5'h11):(4'hf)] ?
                          $unsigned(forvar624) : $unsigned(forvar624))) : {$signed((~&(8'hbc))),
                          $signed((!wire356))}) ?
                  reg620 : ($signed((8'ha0)) ^ (reg625 ?
                      ((reg619 ?
                          wire3 : reg628) != $unsigned(reg631)) : wire2)));
            end
        end
      else
        begin
          for (forvar620 = (1'h0); (forvar620 < (2'h2)); forvar620 = (forvar620 + (1'h1)))
            begin
              reg621 <= $signed(wire616[(4'hc):(4'hb)]);
              reg622 <= (wire17 >= $unsigned($unsigned($unsigned($signed(forvar624)))));
              reg623 <= (&(reg621[(5'h11):(3'h7)] >= (reg623[(1'h0):(1'h0)] <<< wire616[(4'hc):(4'ha)])));
            end
          reg624 = {$unsigned(($unsigned($signed(reg621)) ?
                  $signed($signed(wire356)) : (8'had))),
              (~&(wire356 ?
                  {reg619} : ($unsigned(forvar620) ?
                      $signed(wire618) : reg626[(3'h7):(3'h5)])))};
        end
      for (forvar632 = (1'h0); (forvar632 < (2'h3)); forvar632 = (forvar632 + (1'h1)))
        begin
          if (reg623[(1'h0):(1'h0)])
            begin
              reg633 <= reg626[(3'h4):(1'h0)];
              reg634 <= $unsigned(wire2[(3'h5):(3'h5)]);
            end
          else
            begin
              reg635 = {reg626};
            end
          if ((($signed({$unsigned(forvar620), $unsigned(reg622)}) ?
              $unsigned((~|reg635[(4'ha):(4'h8)])) : (reg630 ?
                  ($signed(wire1) ?
                      (reg629 ?
                          reg634 : (8'hb9)) : (~&reg628)) : ({wire17} <<< $signed(wire0)))) <<< (|reg622)))
            begin
              reg636 <= $signed((8'hb1));
              reg637 = $unsigned(((|(reg634 ?
                      (reg629 | (8'hbf)) : wire0[(2'h3):(2'h3)])) ?
                  wire17 : (&$signed((reg625 ? reg635 : reg633)))));
              reg638 <= ((({$unsigned(forvar632),
                      $unsigned(reg619)} * (~(wire0 >>> reg619))) == reg623) ?
                  $signed(((forvar622[(3'h6):(3'h6)] <= $unsigned(reg636)) == wire3[(5'h11):(1'h0)])) : $signed((reg636 ?
                      $signed(reg621) : ($unsigned(wire0) ?
                          $unsigned(reg625) : wire0))));
              reg639 = {$signed($unsigned(reg627[(5'h11):(4'hd)]))};
            end
          else
            begin
              reg636 <= (-$signed(wire3[(4'he):(4'h9)]));
            end
          if ((($signed($signed((reg625 != wire356))) ^~ reg622) ?
              $signed((~|wire17)) : ((((reg635 ? wire3 : wire356) ?
                      reg619[(5'h11):(5'h11)] : (+forvar622)) > $signed($unsigned(reg636))) ?
                  ($unsigned((reg630 ? reg635 : reg637)) | (^~{reg621,
                      reg630})) : (&({(8'ha5), wire356} ?
                      reg634 : wire17[(4'ha):(3'h4)])))))
            begin
              reg640 = (wire17[(4'h8):(3'h5)] ?
                  $unsigned((wire618[(3'h4):(1'h1)] ~^ (forvar632[(1'h0):(1'h0)] ?
                      (wire17 <= wire356) : (|wire618)))) : wire618);
              reg641 = (~wire1[(2'h3):(1'h1)]);
              reg642 <= wire1[(1'h1):(1'h0)];
            end
          else
            begin
              reg642 <= reg630;
            end
          reg643 <= ((8'h9c) < reg638);
          for (forvar644 = (1'h0); (forvar644 < (1'h1)); forvar644 = (forvar644 + (1'h1)))
            begin
              reg645 = reg638;
              reg646 <= (($unsigned(reg630) ?
                  $unsigned($unsigned((reg624 ?
                      wire616 : wire356))) : reg627[(3'h5):(3'h4)]) + (+$unsigned((&(8'ha9)))));
            end
        end
      if ($unsigned({$unsigned(reg627[(5'h10):(5'h10)]),
          reg642[(2'h3):(2'h3)]}))
        begin
          for (forvar647 = (1'h0); (forvar647 < (1'h1)); forvar647 = (forvar647 + (1'h1)))
            begin
              reg648 <= ((($unsigned((~(8'ha0))) ?
                      (^$signed(forvar620)) : ((+reg628) >> (reg641 || reg645))) & ((~&{wire356,
                      wire17}) == {$unsigned((8'h9e)), $signed(reg624)})) ?
                  $unsigned((((reg619 ?
                      forvar622 : forvar632) * $signed(forvar647)) - $signed((~&reg621)))) : $signed(reg628));
              reg649 = (-(reg635[(4'hb):(1'h0)] ?
                  reg639[(3'h7):(2'h2)] : (reg636[(4'he):(3'h6)] ?
                      (8'hb5) : $signed($unsigned(reg642)))));
              reg650 <= $signed($unsigned(forvar647));
            end
          reg651 = {($signed($unsigned($signed(forvar624))) ?
                  wire0[(5'h11):(3'h5)] : reg623[(4'h9):(3'h7)]),
              (~^(reg650[(4'h9):(1'h1)] + (~^(reg624 <<< (8'hb6)))))};
        end
      else
        begin
          for (forvar647 = (1'h0); (forvar647 < (2'h2)); forvar647 = (forvar647 + (1'h1)))
            begin
              reg648 <= $signed((~^$unsigned(reg626)));
            end
          reg650 <= {$unsigned(reg623),
              ((reg620 ? {(~^reg631)} : (~|{wire17, (8'had)})) ?
                  wire2 : reg621)};
        end
      reg652 <= ((!(wire0[(5'h12):(1'h0)] ?
          $unsigned((wire0 >> reg619)) : (reg642[(1'h1):(1'h1)] != (~reg636)))) >> reg628);
    end
  assign wire653 = wire2;
  always
    @(posedge clk) begin
      if (wire356)
        begin
          if (($signed({reg622[(1'h1):(1'h1)], $signed($signed((8'ha2)))}) ?
              ((~&reg650[(2'h2):(1'h1)]) ?
                  (8'hbd) : ($unsigned($signed((8'haf))) ?
                      (reg652 ?
                          wire17[(3'h7):(1'h1)] : wire3[(4'hc):(1'h0)]) : ((-reg636) ?
                          (wire1 ?
                              wire3 : (7'h44)) : (~(8'ha6))))) : (~&(^~reg630[(2'h3):(1'h1)]))))
            begin
              reg654 <= $signed(((^$signed($unsigned(reg642))) ?
                  $signed($unsigned((wire2 ?
                      reg636 : reg642))) : {$unsigned((^reg642)),
                      reg631[(1'h1):(1'h0)]}));
              reg655 <= {((~wire2[(3'h6):(3'h5)]) >> (-$signed($unsigned(reg648)))),
                  ((reg643[(1'h0):(1'h0)] >= (8'h9e)) ?
                      wire0[(4'he):(4'h8)] : reg646)};
              reg656 <= reg646[(4'hd):(1'h0)];
              reg657 = $signed(reg630[(4'h8):(1'h1)]);
              reg658 = (+reg646);
            end
          else
            begin
              reg654 <= $unsigned((8'hb8));
              reg657 = reg623;
              reg658 = wire616[(1'h1):(1'h1)];
              reg659 <= (reg621 ?
                  reg627[(3'h6):(2'h3)] : $unsigned($signed(($signed(wire653) ~^ (8'hbf)))));
              reg660 = ($signed(reg636[(3'h4):(2'h3)]) == $signed((reg654[(4'ha):(1'h1)] ?
                  {$unsigned(reg657), reg643} : (8'hb6))));
            end
        end
      else
        begin
          for (forvar654 = (1'h0); (forvar654 < (1'h0)); forvar654 = (forvar654 + (1'h1)))
            begin
              reg655 <= $signed(wire1[(1'h1):(1'h0)]);
              reg656 <= ({wire3[(4'he):(1'h0)], reg648[(4'hf):(4'hc)]} ?
                  {(({forvar654} ~^ ((7'h40) ?
                          reg631 : reg660)) ^ $signed((7'h43))),
                      reg646} : {reg659[(5'h12):(1'h0)], $signed(reg646)});
            end
          if (((reg630[(1'h1):(1'h1)] ?
              reg657 : (wire616 > ((wire653 ? reg658 : reg655) ?
                  $unsigned(reg623) : (reg659 ?
                      wire2 : (8'hab))))) == ($unsigned($signed((-reg658))) ?
              reg621[(4'hc):(1'h1)] : reg654)))
            begin
              reg659 <= (&reg634);
              reg661 <= ((((((8'ha8) ? reg642 : reg654) || {reg638}) ?
                      $signed(wire1) : (-(8'hab))) < ((forvar654[(2'h2):(2'h2)] ?
                          $unsigned(reg652) : $signed(reg650)) ?
                      $unsigned(((8'hae) + reg642)) : ($unsigned(wire356) >>> reg629[(1'h1):(1'h0)]))) ?
                  reg643[(3'h5):(2'h3)] : ({$signed((|wire2))} | ($signed((reg633 >> wire1)) ?
                      $signed((~|reg622)) : (+reg646))));
              reg662 = $unsigned((~^$signed(($signed(reg658) >> (~&wire17)))));
              reg663 <= {$signed((reg621 ? reg634 : (~(reg652 ~^ wire1))))};
              reg664 = $signed((+$signed($signed(reg658))));
            end
          else
            begin
              reg659 <= reg638;
              reg660 = ((((reg650[(3'h5):(3'h5)] > ((8'ha9) << reg622)) ?
                  $unsigned(reg655[(4'ha):(3'h7)]) : reg629[(2'h2):(1'h0)]) == (^~($unsigned(reg642) >>> wire3))) | ((((reg663 <= (8'ha2)) <= (reg629 - wire356)) ?
                      ($unsigned((8'hb9)) - $signed(reg629)) : ({reg652,
                              wire0} ?
                          $unsigned(reg664) : $signed(forvar654))) ?
                  {forvar654[(1'h1):(1'h1)],
                      $unsigned((~|reg664))} : ((^~(reg643 ?
                          reg623 : (8'hb1))) ?
                      ($signed(reg622) & (reg627 ?
                          reg652 : reg652)) : $signed({reg661}))));
            end
        end
      if ($unsigned({($signed($signed(reg654)) != reg633)}))
        begin
          if ($unsigned(reg622))
            begin
              reg665 = (~$signed(reg638));
              reg666 <= reg658[(2'h3):(1'h1)];
              reg667 = (reg638[(2'h3):(1'h0)] == forvar654);
              reg668 <= ({$signed((+$signed(reg660))), reg619} ?
                  (|($unsigned(reg665[(4'hb):(4'h8)]) >>> {reg646})) : $unsigned($signed($signed({reg665,
                      reg648}))));
              reg669 <= (&({reg621[(4'hd):(1'h0)], (8'had)} ?
                  $signed(({reg663} <= (8'hbe))) : $unsigned(wire17)));
            end
          else
            begin
              reg666 <= (+((+reg633[(1'h1):(1'h0)]) ?
                  wire1[(4'hf):(4'he)] : ($signed($signed(reg660)) ?
                      $signed((reg629 ? (8'ha3) : reg629)) : reg627)));
              reg668 <= (~^{{reg661, {$unsigned(reg656), wire17}}});
            end
          reg670 <= reg664;
          if ($unsigned((8'hb1)))
            begin
              reg671 = (((((reg636 ? reg646 : wire17) ?
                          (reg656 && reg655) : (reg661 ? reg622 : reg619)) ?
                      (-forvar654) : (wire17 ?
                          reg643 : reg621[(5'h11):(3'h4)])) >> $unsigned($unsigned(((8'hb5) <<< reg650)))) ?
                  (8'hbd) : (~^(reg656 ? wire3 : $signed((+reg666)))));
              reg672 <= ($signed({$signed(wire653)}) && (((reg665[(4'hb):(4'h8)] <<< (+reg658)) ?
                  $unsigned({(8'ha5),
                      forvar654}) : ($signed(wire17) ~^ (-wire616))) << $unsigned((reg670[(2'h3):(2'h3)] != $signed(reg633)))));
              reg673 <= reg670[(1'h0):(1'h0)];
              reg674 = {{(8'hbc),
                      ($unsigned((reg631 & reg629)) ?
                          reg654[(3'h4):(2'h3)] : (reg669[(1'h1):(1'h1)] != $unsigned(forvar654)))}};
              reg675 = $unsigned((wire2 ? reg636[(2'h3):(1'h1)] : reg650));
            end
          else
            begin
              reg672 <= (reg663 && reg642);
              reg674 = {wire356};
              reg675 = $signed(((wire1[(4'ha):(1'h1)] >>> $unsigned((reg672 >= reg657))) ?
                  $unsigned(reg662[(1'h1):(1'h0)]) : (8'ha5)));
              reg676 = ($unsigned(reg661[(1'h0):(1'h0)]) == reg648);
              reg677 <= $unsigned((~|reg631[(3'h6):(1'h0)]));
            end
          reg678 <= $signed($signed((!$signed(reg666[(3'h5):(3'h5)]))));
          reg679 <= (reg646 ?
              reg631[(3'h5):(2'h2)] : $signed($unsigned(reg666[(4'h8):(3'h6)])));
        end
      else
        begin
          if (reg671[(3'h7):(3'h4)])
            begin
              reg666 <= ({$unsigned((~&$unsigned(reg672)))} ?
                  $signed((|$signed((~reg664)))) : (~&reg643[(3'h6):(3'h6)]));
              reg668 <= (~&reg655);
              reg669 <= {$unsigned(($signed(reg677) ^~ {$unsigned(reg636)})),
                  (~&($unsigned($signed((8'h9c))) ~^ (^~$signed(reg673))))};
              reg670 <= $signed((reg666 ~^ (reg659[(4'hf):(1'h0)] ~^ (!{reg629,
                  reg648}))));
              reg672 <= reg650;
            end
          else
            begin
              reg665 = wire3;
              reg667 = {($signed($unsigned($unsigned(reg666))) ?
                      $unsigned(reg643) : reg633[(1'h0):(1'h0)])};
              reg668 <= (~&$signed({$signed(forvar654[(2'h2):(2'h2)])}));
              reg669 <= ($unsigned((((~|reg634) & $unsigned((7'h44))) >> $unsigned(((8'hba) ?
                      reg671 : reg677)))) ?
                  $unsigned((8'ha6)) : (reg638[(3'h4):(2'h3)] != (reg619[(3'h7):(3'h6)] ?
                      $unsigned($signed(reg674)) : ($unsigned((8'ha2)) > ((8'ha7) << wire616)))));
              reg671 = wire653;
            end
          for (forvar673 = (1'h0); (forvar673 < (2'h3)); forvar673 = (forvar673 + (1'h1)))
            begin
              reg674 = ($unsigned({((forvar673 | reg671) <= $signed(reg654)),
                  ((reg659 ?
                      wire616 : (8'hb7)) ^~ (~reg623))}) <<< $signed((&reg648[(3'h4):(2'h3)])));
              reg677 <= $unsigned(({$unsigned((~&reg634))} ?
                  reg657[(3'h7):(2'h2)] : $signed(reg646[(5'h15):(2'h2)])));
              reg680 = reg664;
              reg681 <= {$unsigned((~^(reg642[(3'h4):(1'h1)] & (8'ha3))))};
            end
          reg682 = {(reg680 <= (((^reg667) ? (~&reg667) : $unsigned(wire653)) ?
                  (^~(wire17 || reg661)) : (~^$signed((8'hbe)))))};
        end
      if ({(((reg655[(4'hd):(4'h8)] ?
              (~|reg672) : reg667[(3'h6):(3'h4)]) == $unsigned({reg657,
              reg648})) >>> ((reg665[(4'h8):(3'h5)] ?
              (reg678 | (7'h43)) : {reg680, reg631}) >= (-(reg658 ?
              (7'h40) : (8'hb0))))),
          (~$unsigned(((reg672 ^ reg664) ?
              $unsigned(reg652) : (reg619 ? reg623 : reg670))))})
        begin
          reg683 = $signed(reg636[(4'hf):(2'h2)]);
        end
      else
        begin
          if ((($unsigned((wire17[(4'ha):(2'h3)] ^ reg648[(2'h3):(2'h3)])) << (($signed(reg646) >> $signed(forvar673)) ?
              ((+reg680) > reg674[(4'h8):(3'h6)]) : ({(8'ha4), reg655} ?
                  ((8'ha1) > reg634) : $unsigned(reg658)))) < $unsigned(reg666)))
            begin
              reg683 = (^reg631[(3'h5):(1'h1)]);
              reg684 <= ((8'ha5) | $unsigned((|$signed($signed(reg680)))));
              reg685 = $unsigned({($signed(wire17[(3'h6):(1'h0)]) ?
                      (^reg678[(3'h6):(2'h3)]) : $unsigned($signed(reg631)))});
            end
          else
            begin
              reg683 = $unsigned(reg684[(3'h6):(3'h6)]);
              reg684 <= reg670;
              reg685 = reg660;
              reg686 = $unsigned({$unsigned((~(wire616 ? reg652 : reg660))),
                  $unsigned(($unsigned((8'hac)) || $unsigned(reg631)))});
            end
        end
      if ($unsigned($unsigned(reg657)))
        begin
          if ((^reg664[(1'h1):(1'h1)]))
            begin
              reg687 = $unsigned(((($signed(reg664) ?
                      reg623[(1'h0):(1'h0)] : $signed(reg643)) ?
                  {reg648[(5'h11):(1'h1)]} : {reg652[(4'ha):(4'h8)],
                      (reg627 ? reg654 : reg668)}) <= wire356));
              reg688 = reg670[(4'hf):(2'h3)];
              reg689 <= reg657;
              reg690 = $unsigned($unsigned(reg668));
              reg691 <= (((^((reg690 <= reg646) + (reg660 <= reg665))) < reg627) * $unsigned(reg680[(4'h9):(3'h4)]));
            end
          else
            begin
              reg687 = ((((-{(7'h43)}) * (~|forvar673)) == ((~&$unsigned(reg634)) ?
                      ($unsigned(wire3) ?
                          $signed(reg672) : (^~reg664)) : wire616)) ?
                  ((^$unsigned((reg667 & forvar654))) ?
                      reg671[(4'h8):(3'h6)] : {(~&$unsigned(reg631))}) : (((reg667[(2'h3):(1'h0)] ?
                          forvar654 : (^reg663)) ?
                      (8'hae) : ($unsigned(reg630) ?
                          (reg662 + reg658) : {reg636})) >= reg665[(3'h6):(3'h4)]));
              reg688 = reg648[(4'hb):(3'h7)];
              reg690 = $unsigned((wire3 ? wire1 : $signed(wire17)));
              reg691 <= reg622;
            end
          for (forvar692 = (1'h0); (forvar692 < (3'h4)); forvar692 = (forvar692 + (1'h1)))
            begin
              reg693 = $signed($unsigned((&(~(~^(8'h9d))))));
              reg694 <= (8'h9c);
              reg695 = $signed(((reg646[(2'h3):(1'h0)] ?
                      reg672[(1'h0):(1'h0)] : wire0[(4'h9):(4'h8)]) ?
                  $signed(((reg681 == (7'h40)) ?
                      reg667 : $unsigned(reg668))) : $signed($signed((^reg646)))));
              reg696 <= $unsigned($unsigned((^((^reg664) ~^ (reg660 * reg661)))));
            end
          reg697 <= $signed(reg664[(1'h0):(1'h0)]);
        end
      else
        begin
          if ((reg661 >= (((^~{reg688, reg676}) ?
              (((8'hbd) ? reg634 : reg633) ?
                  $unsigned(reg643) : (+(8'ha7))) : reg638[(3'h5):(1'h0)]) || $signed({$unsigned((8'ha9)),
              $unsigned(wire618)}))))
            begin
              reg687 = ($signed($signed((8'hb8))) < $signed({$signed(reg671)}));
              reg688 = (((((~^reg691) ^~ reg662) || ($signed(reg682) * (^~reg622))) ?
                  reg636[(4'hf):(1'h1)] : reg676[(4'hc):(3'h6)]) || $unsigned($unsigned(((-reg682) <= (wire1 << forvar692)))));
              reg689 <= ($signed(({reg693[(2'h2):(1'h0)]} >= (8'ha8))) || ($signed(reg674[(4'ha):(2'h2)]) <= (8'hbc)));
            end
          else
            begin
              reg689 <= forvar673[(5'h12):(5'h12)];
              reg691 <= ((&$signed({$signed(wire0)})) ?
                  ($signed(wire3) <= reg688[(3'h7):(1'h0)]) : (~|$unsigned(reg629)));
              reg692 = (($signed(({reg675} ?
                      $unsigned((8'ha5)) : (8'had))) && wire0) ?
                  ($unsigned($signed($signed(reg665))) + (+(^~$unsigned(reg623)))) : $unsigned((~reg638[(1'h1):(1'h0)])));
              reg694 <= ($unsigned(($signed($unsigned(reg692)) ?
                  $unsigned({reg642}) : reg621)) <= (+((~^(&(8'ha9))) << (^reg636[(4'hb):(1'h1)]))));
              reg696 <= (+(7'h41));
            end
          if (((^~(+reg680)) ? (&reg671) : reg692))
            begin
              reg698 = $signed(((|((forvar654 ? reg664 : reg621) ?
                      (reg664 < reg630) : reg654)) ?
                  (+($unsigned(reg629) ^ (reg673 - forvar654))) : reg648));
              reg699 <= (|(~|reg696[(3'h4):(2'h3)]));
            end
          else
            begin
              reg698 = (forvar673[(1'h0):(1'h0)] ?
                  ((($unsigned(reg668) ?
                          ((8'hae) ? reg699 : reg654) : (reg657 ?
                              reg670 : reg665)) && ($unsigned(wire356) && ((8'hb1) ?
                          reg658 : reg662))) ?
                      $unsigned(({reg675} ?
                          ((8'hb1) && reg656) : $unsigned(reg676))) : (($unsigned((8'h9e)) <= $unsigned((7'h42))) ?
                          (reg629 & $unsigned(wire616)) : $signed($unsigned((8'h9c))))) : {$unsigned((^{reg680,
                          reg692})),
                      $signed({(reg679 + reg670)})});
              reg700 = reg648;
              reg701 <= reg638;
              reg702 <= $signed($signed((reg652 + reg684[(1'h1):(1'h1)])));
            end
        end
      reg703 <= (^~(($signed($signed(reg631)) ^ ((~&reg622) ?
          ((8'ha0) ? (8'hb6) : reg659) : (reg698 + wire17))) > reg671));
    end
  assign wire704 = ($unsigned(($unsigned($signed(reg627)) | ({reg697, reg672} ?
                       {reg630,
                           reg679} : $unsigned(wire3)))) & (reg659[(4'hb):(4'h9)] ?
                       $signed(((reg703 ?
                           (8'hbf) : reg655) << reg633[(2'h2):(2'h2)])) : {$unsigned(reg670),
                           $unsigned((reg633 ? reg691 : reg643))}));
  assign wire705 = (((~&reg652[(3'h5):(2'h2)]) | reg622) << reg622);
  assign wire706 = (((~&reg696) ? reg638[(3'h4):(1'h1)] : (8'ha4)) ?
                       wire705[(1'h1):(1'h0)] : reg668);
  assign wire707 = ($unsigned((!$unsigned($unsigned(reg650)))) ?
                       (8'hac) : ($unsigned(($signed(reg691) ?
                               ((8'ha7) > wire616) : (^(8'hab)))) ?
                           (reg648[(3'h7):(3'h5)] < (reg689[(2'h3):(2'h2)] ?
                               (reg630 ?
                                   wire706 : reg655) : reg672)) : $signed($unsigned($unsigned(reg646)))));
  assign wire708 = (((^wire616) <= $signed($unsigned($unsigned((8'hb0))))) & reg699[(4'hd):(4'ha)]);
  always
    @(posedge clk) begin
      for (forvar709 = (1'h0); (forvar709 < (1'h0)); forvar709 = (forvar709 + (1'h1)))
        begin
          if ({{$unsigned($signed((~(8'hb2)))),
                  {((~&wire653) != (reg636 || reg655))}}})
            begin
              reg710 <= reg672;
              reg711 <= $signed($unsigned(reg622[(3'h6):(3'h5)]));
              reg712 <= (($signed(((reg622 ?
                          wire708 : (8'hab)) ^~ (reg678 & reg672))) ?
                      $signed(($unsigned((8'hbd)) ?
                          wire708[(3'h6):(1'h1)] : reg629[(2'h2):(2'h2)])) : $signed($unsigned($unsigned(reg697)))) ?
                  $unsigned($signed(($signed(reg619) ?
                      reg633 : {reg669,
                          reg655}))) : (((|reg663[(3'h6):(2'h3)]) ?
                      $signed($signed(reg694)) : ((|reg643) != reg636)) >> reg623[(2'h3):(2'h2)]));
              reg713 <= wire0[(3'h6):(2'h3)];
            end
          else
            begin
              reg710 <= ($unsigned((+(~^(reg656 < reg689)))) >>> reg691[(3'h5):(2'h3)]);
              reg714 = ((^reg711) <<< reg629[(2'h2):(1'h1)]);
              reg715 = (reg699[(2'h2):(2'h2)] ?
                  (-(((reg673 ? reg714 : wire653) && $signed(reg659)) ?
                      ({(8'ha5), wire356} ?
                          (wire2 ^ reg652) : $unsigned(reg670)) : reg642)) : ((reg661[(4'hc):(3'h4)] | ((reg677 ?
                          (8'hbb) : wire707) >>> (wire653 + wire707))) ?
                      {reg679[(4'h8):(1'h0)],
                          reg629[(1'h1):(1'h0)]} : (8'hb1)));
            end
          for (forvar716 = (1'h0); (forvar716 < (1'h0)); forvar716 = (forvar716 + (1'h1)))
            begin
              reg717 <= (reg659 & reg697);
              reg718 <= $signed(({$signed({reg714})} ?
                  (reg677 ?
                      $unsigned($unsigned(wire705)) : reg621[(4'h8):(3'h6)]) : $unsigned($unsigned((reg652 - reg636)))));
              reg719 = ((^((^~$signed(wire704)) >> ((-reg655) ?
                  wire704 : $unsigned(reg712)))) ~^ $unsigned($unsigned(((reg668 | reg678) | (reg714 ?
                  reg619 : reg656)))));
              reg720 = $unsigned($signed(reg646[(5'h14):(5'h14)]));
              reg721 <= (+wire17);
            end
          reg722 <= $signed($unsigned(reg719));
          for (forvar723 = (1'h0); (forvar723 < (1'h0)); forvar723 = (forvar723 + (1'h1)))
            begin
              reg724 = {$signed(wire618[(2'h3):(1'h0)])};
              reg725 <= reg717[(4'h9):(3'h7)];
              reg726 <= (&(^~reg623));
            end
        end
      for (forvar727 = (1'h0); (forvar727 < (1'h1)); forvar727 = (forvar727 + (1'h1)))
        begin
          for (forvar728 = (1'h0); (forvar728 < (1'h1)); forvar728 = (forvar728 + (1'h1)))
            begin
              reg729 <= reg697[(4'hb):(1'h1)];
              reg730 = (8'hb1);
              reg731 = $signed($signed({(^wire618)}));
              reg732 <= reg666;
            end
          for (forvar733 = (1'h0); (forvar733 < (1'h0)); forvar733 = (forvar733 + (1'h1)))
            begin
              reg734 <= (reg633[(1'h1):(1'h0)] ?
                  $signed((forvar727 ?
                      (^~reg721[(5'h15):(3'h6)]) : (reg655 <<< wire0[(2'h2):(1'h1)]))) : (($signed({reg663}) ?
                      reg663[(4'h8):(4'h8)] : (&(reg729 ?
                          reg622 : reg646))) >>> {$signed((8'hb4))}));
              reg735 = (^~$signed((~&$signed($signed(forvar733)))));
              reg736 <= reg666[(3'h4):(3'h4)];
            end
          reg737 <= (((~|reg735[(4'hc):(4'h9)]) ?
                  reg654 : (reg633 ? $signed($unsigned(reg623)) : reg724)) ?
              ((-{reg623, $signed((8'hbc))}) ~^ {$unsigned(reg703),
                  reg627[(2'h3):(2'h3)]}) : {(!(8'ha3))});
        end
      if ($signed({$unsigned((~$unsigned(reg631)))}))
        begin
          if (($unsigned(($signed($signed(wire705)) ?
              {wire707[(3'h5):(3'h4)],
                  (reg634 ?
                      forvar728 : reg701)} : ($unsigned(reg736) <= reg691[(3'h5):(1'h1)]))) & $signed(reg719)))
            begin
              reg738 <= {wire618[(1'h1):(1'h0)], reg650};
              reg739 <= (reg672 >= $unsigned((((wire17 ? reg721 : forvar727) ?
                      reg734 : (wire707 >= reg663)) ?
                  (+$signed((8'hb9))) : {(7'h43)})));
              reg740 = ($signed($unsigned($signed((8'hb1)))) ?
                  $signed((~|$unsigned($unsigned((8'ha9))))) : $unsigned($unsigned(($signed(reg650) > (-reg638)))));
              reg741 <= reg740;
              reg742 <= (($unsigned((-((8'hbe) ~^ reg629))) ^ ($unsigned((^reg696)) <<< (!(reg659 ?
                      reg673 : reg725)))) ?
                  (($unsigned(reg679) ?
                      ((reg668 ? reg739 : reg627) ?
                          reg726[(3'h4):(2'h3)] : (reg677 + reg739)) : $unsigned(((8'hb6) >> (8'hba)))) <= reg638[(3'h4):(1'h1)]) : reg652);
            end
          else
            begin
              reg740 = {$signed(wire2)};
            end
        end
      else
        begin
          if (({$unsigned({{reg721}}), $signed(reg699)} ?
              reg638 : ((8'hb9) ?
                  reg679[(2'h2):(2'h2)] : reg619[(5'h10):(4'hb)])))
            begin
              reg738 <= {reg621[(5'h10):(4'he)]};
              reg739 <= reg701;
              reg741 <= ($signed($unsigned((~&(reg673 <<< (7'h40))))) == {wire705,
                  reg694});
            end
          else
            begin
              reg740 = $signed({(~^reg697), reg719});
            end
          reg743 = $signed({($unsigned($unsigned(reg721)) << (reg714 ?
                  (reg694 ? reg718 : reg670) : reg738[(4'hc):(3'h4)])),
              reg646});
          if ({$signed(reg669)})
            begin
              reg744 <= wire707[(4'hd):(2'h3)];
              reg745 <= reg638[(3'h4):(1'h1)];
            end
          else
            begin
              reg744 <= (wire356[(1'h1):(1'h1)] ?
                  $unsigned((8'hb7)) : ((((forvar723 ?
                          reg738 : reg739) ^ (reg652 + reg668)) ?
                      reg646[(4'hf):(4'hc)] : (((8'hab) << reg638) | reg654[(3'h6):(1'h0)])) <<< $unsigned($unsigned(reg713))));
              reg746 = (+({forvar716[(1'h1):(1'h0)]} & $unsigned((~(reg712 ?
                  reg745 : (8'h9c))))));
              reg747 <= (reg703[(3'h7):(3'h5)] ?
                  $unsigned(((reg718[(3'h7):(3'h5)] ? {reg725} : (8'ha5)) ?
                      ((7'h40) ?
                          $signed(reg670) : (reg714 - (8'hbb))) : ($signed(reg720) ?
                          reg666 : (forvar723 ^~ reg677)))) : (reg629 ?
                      reg679 : $signed((~|reg703[(3'h6):(3'h6)]))));
              reg748 <= {((^(&$unsigned(reg730))) << (reg721 == $signed((reg722 * reg742))))};
            end
          if ($signed(((reg737 ?
              $unsigned((reg650 ?
                  reg719 : reg638)) : $unsigned((~^reg701))) || reg648[(3'h4):(2'h3)])))
            begin
              reg749 <= reg713[(3'h5):(3'h4)];
              reg750 <= {reg731[(2'h3):(2'h3)]};
              reg751 <= (^{($unsigned(((8'hb3) ? reg736 : forvar727)) ?
                      (~(forvar716 + reg722)) : (^$signed(reg679))),
                  reg648});
            end
          else
            begin
              reg749 <= $signed(reg746);
              reg752 = ((reg679[(1'h0):(1'h0)] ?
                  (~|(reg643[(4'ha):(4'h8)] ^ wire706[(1'h0):(1'h0)])) : {reg663[(2'h2):(1'h0)],
                      $signed((8'haa))}) >>> reg633[(2'h2):(1'h1)]);
            end
        end
      if (wire2)
        begin
          if ((~reg744[(3'h5):(2'h2)]))
            begin
              reg753 <= ($unsigned(($unsigned({reg750, reg732}) ?
                      $signed((reg621 + (8'h9c))) : (!(^reg633)))) ?
                  $signed((reg743[(3'h4):(1'h0)] ?
                      reg735 : (reg736 >>> reg715))) : reg721[(5'h15):(2'h2)]);
              reg754 <= ($unsigned({(-$unsigned(reg672))}) == {reg744[(4'h8):(1'h0)],
                  $signed(reg621[(4'hb):(1'h0)])});
            end
          else
            begin
              reg753 <= reg694;
              reg755 = reg661;
              reg756 = ({(reg712[(2'h3):(1'h0)] ?
                          $unsigned($signed(reg670)) : reg713)} ?
                  (((!reg753) <= $signed((reg642 ? reg629 : reg650))) ?
                      reg754[(5'h14):(4'h8)] : (reg742 ^ ((~&reg739) ?
                          (reg661 && reg631) : $unsigned((8'hb6))))) : ($signed((reg742[(1'h0):(1'h0)] != (~reg655))) ?
                      $unsigned(wire705[(3'h5):(3'h4)]) : (^~$unsigned({reg720}))));
              reg757 <= reg721[(5'h15):(2'h2)];
              reg758 <= $signed($unsigned($signed(reg713[(1'h0):(1'h0)])));
            end
          for (forvar759 = (1'h0); (forvar759 < (1'h0)); forvar759 = (forvar759 + (1'h1)))
            begin
              reg760 = (8'ha1);
            end
          reg761 = (($signed((((8'h9e) + (8'hb1)) > (reg627 ?
                      wire708 : forvar709))) ?
                  (forvar733 * reg638[(3'h6):(2'h3)]) : $unsigned(reg711[(2'h3):(1'h1)])) ?
              {{(8'had), reg726[(3'h5):(1'h0)]},
                  wire618} : (reg642[(4'hd):(3'h4)] ?
                  $signed($unsigned((-reg717))) : reg634));
        end
      else
        begin
          if (reg654)
            begin
              reg753 <= ((~|(wire616[(4'hb):(2'h2)] && ((8'hb3) >= $unsigned(reg735)))) & (reg751[(2'h3):(1'h1)] == (+$signed(reg679))));
              reg754 <= ($signed($unsigned($signed((reg711 - reg631)))) >>> (~^(|forvar709[(2'h2):(1'h1)])));
              reg755 = ($signed({(~$unsigned(reg752))}) ?
                  $signed({$unsigned(((7'h40) >= wire1)),
                      reg684[(3'h4):(2'h3)]}) : {reg741[(2'h2):(1'h1)],
                      ((reg747 < (&reg712)) >= {((7'h43) ? reg753 : reg731)})});
            end
          else
            begin
              reg753 <= (reg703[(4'hc):(3'h7)] && (-$unsigned($unsigned(reg753[(4'h9):(3'h7)]))));
              reg754 <= reg720[(2'h3):(2'h2)];
              reg755 = $unsigned(reg734);
              reg756 = $unsigned($unsigned(wire356[(3'h4):(3'h4)]));
            end
          reg759 = {(+$unsigned(wire356[(3'h6):(2'h3)]))};
        end
      for (forvar762 = (1'h0); (forvar762 < (1'h0)); forvar762 = (forvar762 + (1'h1)))
        begin
          reg763 <= reg711;
        end
    end
  assign wire764 = ({(~^(8'ha4))} + {{$signed(reg634[(4'h9):(3'h6)])},
                       $signed((&wire3))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module358
#(parameter param614 = (!(8'hb0)), 
parameter param615 = (((((8'hab) - (param614 ^ param614)) ? (^((8'haa) | param614)) : (~^(^~param614))) ? {(^~(param614 ? param614 : param614))} : ((8'hbf) ~^ param614)) ? (((~(param614 ? param614 : param614)) != ((8'hb3) ? {(8'hbb), (8'h9d)} : {param614, param614})) > {{(param614 ? (7'h44) : param614)}}) : (~param614)))
(y, clk, wire363, wire362, wire361, wire360, wire359);
  output wire [(32'h350):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire363;
  input wire [(4'ha):(1'h0)] wire362;
  input wire [(5'h12):(1'h0)] wire361;
  input wire signed [(4'hb):(1'h0)] wire360;
  input wire [(2'h2):(1'h0)] wire359;
  wire [(4'hf):(1'h0)] wire613;
  wire signed [(3'h5):(1'h0)] wire612;
  wire [(5'h15):(1'h0)] wire611;
  wire [(3'h6):(1'h0)] wire610;
  wire signed [(5'h10):(1'h0)] wire609;
  wire [(5'h14):(1'h0)] wire607;
  wire [(3'h7):(1'h0)] wire570;
  wire signed [(4'ha):(1'h0)] wire569;
  wire [(4'h8):(1'h0)] wire515;
  wire signed [(3'h7):(1'h0)] wire514;
  wire [(2'h2):(1'h0)] wire513;
  wire signed [(4'hb):(1'h0)] wire511;
  wire [(4'hf):(1'h0)] wire463;
  wire signed [(4'he):(1'h0)] wire461;
  reg signed [(4'hc):(1'h0)] reg568 = (1'h0);
  reg signed [(4'he):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg561 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg560 = (1'h0);
  reg [(4'hb):(1'h0)] reg559 = (1'h0);
  reg signed [(4'he):(1'h0)] reg555 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg553 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg550 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg547 = (1'h0);
  reg [(5'h11):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg544 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg543 = (1'h0);
  reg [(4'ha):(1'h0)] reg542 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg531 = (1'h0);
  reg [(3'h4):(1'h0)] reg541 = (1'h0);
  reg [(5'h14):(1'h0)] reg539 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg538 = (1'h0);
  reg [(4'he):(1'h0)] reg536 = (1'h0);
  reg [(4'hf):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg533 = (1'h0);
  reg [(3'h5):(1'h0)] reg532 = (1'h0);
  reg [(5'h15):(1'h0)] reg528 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg527 = (1'h0);
  reg [(5'h15):(1'h0)] reg524 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg523 = (1'h0);
  reg [(3'h6):(1'h0)] reg518 = (1'h0);
  reg [(4'hf):(1'h0)] reg517 = (1'h0);
  reg [(4'hd):(1'h0)] reg516 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg567 = (1'h0);
  reg [(4'h9):(1'h0)] reg566 = (1'h0);
  reg [(2'h3):(1'h0)] forvar565 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar564 = (1'h0);
  reg [(4'hc):(1'h0)] reg563 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg557 = (1'h0);
  reg [(3'h6):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar554 = (1'h0);
  reg [(5'h15):(1'h0)] reg551 = (1'h0);
  reg [(5'h14):(1'h0)] reg549 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg548 = (1'h0);
  reg [(3'h4):(1'h0)] reg545 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg540 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg537 = (1'h0);
  reg [(5'h11):(1'h0)] reg534 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar531 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg530 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg529 = (1'h0);
  reg [(3'h6):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg525 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg522 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg521 = (1'h0);
  reg [(3'h7):(1'h0)] reg520 = (1'h0);
  reg [(4'hf):(1'h0)] reg519 = (1'h0);
  assign y = {wire613,
                 wire612,
                 wire611,
                 wire610,
                 wire609,
                 wire607,
                 wire570,
                 wire569,
                 wire515,
                 wire514,
                 wire513,
                 wire511,
                 wire463,
                 wire461,
                 reg568,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg555,
                 reg553,
                 reg552,
                 reg550,
                 reg547,
                 reg546,
                 reg544,
                 reg543,
                 reg542,
                 reg531,
                 reg541,
                 reg539,
                 reg538,
                 reg536,
                 reg535,
                 reg533,
                 reg532,
                 reg528,
                 reg527,
                 reg524,
                 reg523,
                 reg518,
                 reg517,
                 reg516,
                 reg567,
                 reg566,
                 forvar565,
                 forvar564,
                 reg563,
                 reg558,
                 reg557,
                 reg556,
                 forvar554,
                 reg551,
                 reg549,
                 reg548,
                 reg545,
                 reg540,
                 reg537,
                 reg534,
                 forvar531,
                 reg530,
                 reg529,
                 reg526,
                 reg525,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 (1'h0)};
  module364 #() modinst462 (.y(wire461), .clk(clk), .wire368(wire360), .wire367(wire359), .wire366(wire363), .wire365(wire361));
  assign wire463 = $signed($signed($unsigned(((-wire363) <= (~^(8'ha2))))));
  module464 #() modinst512 (wire511, clk, wire461, wire463, wire363, wire361);
  assign wire513 = (~|(~$signed($unsigned({(8'hb9), wire363}))));
  assign wire514 = (wire513 <<< (($signed(wire359[(1'h1):(1'h0)]) > ($signed(wire461) ?
                       (wire361 ?
                           wire363 : (8'ha9)) : $unsigned(wire513))) >= (($signed(wire511) ?
                       $unsigned(wire463) : wire511) | ($unsigned(wire513) * wire461))));
  assign wire515 = wire463;
  always
    @(posedge clk) begin
      if (wire511)
        begin
          if (((7'h44) | wire360[(1'h0):(1'h0)]))
            begin
              reg516 <= wire361[(4'hc):(1'h0)];
              reg517 <= $unsigned((+$signed(wire514)));
              reg518 <= $unsigned({{(8'haf),
                      $signed(((8'haa) ? wire514 : wire514))},
                  $unsigned((^(|wire361)))});
            end
          else
            begin
              reg516 <= $unsigned($signed((reg518[(3'h4):(2'h2)] ?
                  {$signed(wire463), (wire362 > reg518)} : (&wire513))));
              reg519 = $unsigned($signed($unsigned(wire361[(5'h11):(4'h8)])));
              reg520 = {wire363, (&(~&(^wire362)))};
            end
          reg521 = $signed(wire461);
          if (($signed(($unsigned((-wire515)) ?
                  reg516[(2'h3):(1'h0)] : reg518[(1'h1):(1'h0)])) ?
              {$signed(wire363[(4'h9):(4'h8)]), wire463} : wire461))
            begin
              reg522 = reg517;
              reg523 <= (&(wire511 <<< (reg522 == wire514[(2'h3):(2'h3)])));
            end
          else
            begin
              reg523 <= ($unsigned(wire514[(3'h4):(1'h0)]) != $unsigned($signed($unsigned((&reg519)))));
              reg524 <= wire463;
              reg525 = wire361;
              reg526 = (~^$signed((reg523[(3'h6):(3'h4)] ?
                  $signed($unsigned(reg523)) : reg524[(4'ha):(1'h1)])));
              reg527 <= $signed(wire360[(3'h6):(3'h5)]);
            end
        end
      else
        begin
          if (($signed($unsigned($unsigned((reg524 - reg522)))) ?
              $signed($unsigned(($unsigned(wire461) ?
                  (wire363 ? (8'hab) : reg518) : (reg522 ?
                      (8'hb4) : wire514)))) : (^~$signed(reg525[(4'h9):(2'h2)]))))
            begin
              reg519 = $unsigned(reg521);
              reg523 <= $signed($signed(((|{wire461,
                  reg524}) <= ($unsigned(wire361) - (~reg525)))));
              reg525 = ($unsigned($signed(reg521[(4'h9):(1'h1)])) ?
                  reg527[(4'hc):(3'h7)] : (wire463[(4'hf):(4'h8)] <<< (reg523[(3'h5):(1'h1)] ?
                      {(reg527 ~^ reg520)} : $unsigned($signed((8'ha5))))));
              reg526 = $unsigned($signed($unsigned(reg521)));
            end
          else
            begin
              reg519 = wire360;
              reg523 <= $signed((~&$unsigned((reg523[(2'h3):(1'h1)] > (^~wire361)))));
              reg524 <= wire361[(5'h11):(4'hd)];
            end
          reg527 <= $unsigned(((8'ha0) ~^ wire359));
          reg528 <= $signed(($signed(reg516) ?
              reg527 : $signed(($signed(wire511) | wire513))));
          reg529 = $signed(wire513[(2'h2):(1'h0)]);
        end
      reg530 = ((+wire360[(3'h5):(1'h0)]) ?
          wire514[(1'h0):(1'h0)] : ($signed(reg526[(1'h0):(1'h0)]) != (wire361[(2'h3):(1'h0)] - wire463)));
      if ($signed(reg530))
        begin
          for (forvar531 = (1'h0); (forvar531 < (2'h3)); forvar531 = (forvar531 + (1'h1)))
            begin
              reg532 <= wire359;
              reg533 <= $unsigned($unsigned($unsigned(($unsigned(wire514) ?
                  reg529 : ((8'h9c) ? (8'hab) : (7'h41))))));
            end
          if (({({$unsigned(reg530)} && ((8'hb8) == (reg519 * reg519))),
              wire513} >= reg530))
            begin
              reg534 = $unsigned(reg533);
              reg535 <= (({$signed($unsigned(reg528)),
                      {$signed(reg528)}} & wire511) ?
                  $unsigned(reg518[(2'h3):(1'h0)]) : $signed($unsigned(({wire514,
                          (8'ha9)} ?
                      $signed(forvar531) : (wire514 >>> reg521)))));
              reg536 <= (($signed({((8'ha4) >>> (8'hb5)),
                      ((7'h42) ~^ reg519)}) | (wire363[(3'h4):(1'h1)] ?
                      $unsigned((~|reg529)) : $unsigned($unsigned(wire359)))) ?
                  (^$signed(((forvar531 <<< wire514) ?
                      (~^reg520) : (wire515 ?
                          wire461 : wire515)))) : wire515[(3'h4):(3'h4)]);
              reg537 = (!(7'h43));
            end
          else
            begin
              reg534 = reg528[(4'hd):(3'h6)];
              reg535 <= {$signed(($signed(wire360[(4'ha):(1'h1)]) ?
                      reg530 : (reg522[(1'h1):(1'h1)] ? (~^reg523) : wire515))),
                  $unsigned((-wire511))};
              reg537 = {wire511};
              reg538 <= (({$signed($unsigned(wire513)), {(^~wire362)}} ?
                  wire362 : (~|wire362)) ^ wire363);
              reg539 <= ((~^(&(reg525 ?
                  $signed(reg516) : $signed(reg538)))) && (8'h9e));
            end
          reg540 = reg516;
          reg541 <= ({(((wire461 << reg528) && reg537[(3'h5):(1'h1)]) ?
                  $signed((&reg518)) : (^~(~|reg528))),
              wire362} != reg523);
        end
      else
        begin
          if ((((^$unsigned($unsigned(reg519))) <= $signed(((forvar531 ?
              reg528 : reg521) < (~|wire514)))) <= reg536[(3'h4):(1'h1)]))
            begin
              reg531 <= {(^reg530),
                  $signed($unsigned(((reg538 << reg525) ? wire513 : (8'h9c))))};
            end
          else
            begin
              reg531 <= $signed({(^~$signed({wire359}))});
              reg534 = {((!(reg519[(4'hf):(1'h0)] ?
                      (reg534 && wire511) : reg535[(2'h3):(1'h0)])) == reg535[(2'h3):(2'h3)]),
                  (-$signed((~|$signed(reg539))))};
            end
          if ((8'h9c))
            begin
              reg535 <= ($signed($unsigned(((8'hbf) ?
                      (reg535 * (8'ha7)) : $signed(reg527)))) ?
                  (!$unsigned({wire511[(4'h8):(3'h6)],
                      (8'hb3)})) : (reg517[(4'h9):(3'h5)] + $unsigned((reg529 != $unsigned(reg534)))));
              reg537 = $unsigned($unsigned(($unsigned(reg522[(2'h2):(1'h1)]) & reg533)));
              reg538 <= (8'h9c);
              reg539 <= ((~|(((wire461 && reg530) ?
                  wire362 : $signed((8'hbf))) <= $signed($unsigned(reg528)))) <= reg525[(4'hc):(4'hc)]);
            end
          else
            begin
              reg537 = wire362[(3'h6):(1'h1)];
              reg538 <= $signed(reg519[(4'h9):(2'h2)]);
              reg539 <= (-$unsigned((+reg530[(4'he):(4'hd)])));
              reg540 = wire514;
              reg541 <= ((~|($signed(wire362[(1'h0):(1'h0)]) < reg522[(1'h1):(1'h1)])) ?
                  wire515 : reg522);
            end
          reg542 <= $unsigned(($unsigned(((!wire511) + (reg530 || (8'ha0)))) << $unsigned((^wire360[(3'h5):(2'h2)]))));
          if (((reg535 ^~ {{{wire360, (8'ha0)}}}) ?
              reg540 : (wire360[(4'h8):(2'h2)] ?
                  wire361[(1'h1):(1'h0)] : $signed(reg519[(1'h1):(1'h1)]))))
            begin
              reg543 <= reg518;
              reg544 <= (^reg521[(4'h9):(3'h6)]);
              reg545 = $signed(((!({wire461, reg517} ? (8'hb4) : reg543)) ?
                  $unsigned((reg534[(4'ha):(2'h3)] + forvar531[(4'hd):(3'h6)])) : wire513));
            end
          else
            begin
              reg543 <= (7'h40);
              reg545 = ((&((wire461[(3'h5):(3'h4)] + $signed(wire514)) ?
                      (-{reg531}) : {wire515[(3'h7):(3'h7)], (^reg536)})) ?
                  ($unsigned($unsigned($unsigned(reg517))) != $signed($unsigned($signed(reg527)))) : $signed($unsigned((~$unsigned((8'hab))))));
            end
        end
      if (reg522)
        begin
          if ((reg538[(2'h3):(1'h0)] || $unsigned(((+$signed((8'ha8))) - (~$signed(wire362))))))
            begin
              reg546 <= ((^(&$signed($signed(reg525)))) | (|$unsigned({(reg521 <= reg533),
                  (8'haa)})));
              reg547 <= (^$signed($unsigned(wire359)));
              reg548 = {reg525[(1'h0):(1'h0)]};
              reg549 = $signed((|wire359[(1'h1):(1'h0)]));
            end
          else
            begin
              reg548 = $unsigned({wire513[(1'h0):(1'h0)]});
              reg550 <= $unsigned($unsigned(($signed((reg540 <= reg516)) ?
                  ((~(7'h42)) ?
                      (-(8'hac)) : (reg548 <= reg535)) : (^$signed(reg544)))));
              reg551 = $unsigned($unsigned(((|(~|wire514)) ?
                  {reg539} : $signed($unsigned(reg520)))));
              reg552 <= (~(reg519[(4'hb):(4'hb)] ?
                  wire514 : ($unsigned($signed(reg534)) ^~ $unsigned($unsigned((8'hba))))));
              reg553 <= reg546[(2'h2):(1'h1)];
            end
          for (forvar554 = (1'h0); (forvar554 < (3'h4)); forvar554 = (forvar554 + (1'h1)))
            begin
              reg555 <= reg520;
            end
          reg556 = {{$signed(($signed(reg522) ?
                      (wire511 + (8'had)) : $signed(reg547)))}};
          if ($signed(((~^(^~$signed(reg539))) ?
              ({reg535} ?
                  reg555[(4'h8):(3'h5)] : reg535) : $unsigned((~&(reg550 ?
                  reg551 : reg528))))))
            begin
              reg557 = reg525[(5'h11):(2'h2)];
            end
          else
            begin
              reg557 = (8'ha1);
            end
          if (($unsigned({($unsigned(wire363) ?
                      (reg548 ? reg516 : reg532) : (~|reg541))}) ?
              $unsigned(((&reg519) ?
                  reg530 : ((wire511 > reg552) ^~ (reg540 ?
                      wire360 : reg549)))) : ({($signed(reg529) <= wire514[(3'h5):(3'h5)]),
                  reg534[(3'h6):(3'h5)]} >>> {$unsigned(reg543),
                  $signed((reg522 + reg549))})))
            begin
              reg558 = {$signed(reg518)};
              reg559 <= reg555;
            end
          else
            begin
              reg559 <= (&($unsigned({$signed(reg522)}) == (reg556[(2'h2):(2'h2)] ?
                  forvar554 : reg524[(5'h14):(4'hf)])));
              reg560 <= ((reg534[(1'h0):(1'h0)] ?
                  (reg549 ?
                      ((|reg543) ^ (forvar554 & (8'hb2))) : (8'ha8)) : reg553[(4'h9):(3'h4)]) || (reg556[(3'h4):(2'h3)] ?
                  (8'h9c) : reg522[(2'h2):(1'h0)]));
              reg561 <= (~&$unsigned($signed(((reg523 > reg544) ?
                  (reg531 | wire362) : {wire463, (8'h9e)}))));
              reg562 <= (^(~^$signed({$signed(reg558)})));
              reg563 = ($signed($signed(forvar554[(4'ha):(4'h8)])) > {wire359[(1'h1):(1'h0)],
                  $unsigned(((+reg560) ^~ $signed(reg523)))});
            end
        end
      else
        begin
          reg548 = (~(reg523 ?
              (((7'h43) ?
                  $unsigned(reg546) : reg517) != reg562[(3'h4):(2'h3)]) : ((8'ha3) >= $signed(reg553))));
        end
      for (forvar564 = (1'h0); (forvar564 < (3'h4)); forvar564 = (forvar564 + (1'h1)))
        begin
          for (forvar565 = (1'h0); (forvar565 < (2'h2)); forvar565 = (forvar565 + (1'h1)))
            begin
              reg566 = $signed($signed($signed(((&reg532) > reg549[(5'h13):(2'h3)]))));
              reg567 = (({($signed(reg562) ?
                          reg521 : $signed(reg558))} == (-$unsigned((|(8'ha0))))) ?
                  $unsigned($signed($signed(reg534))) : $unsigned((~&$signed(reg539[(1'h0):(1'h0)]))));
              reg568 <= $unsigned({{((7'h42) ? $signed(reg532) : reg553),
                      $unsigned($signed(forvar531))},
                  forvar565});
            end
        end
    end
  assign wire569 = (^(wire362[(1'h1):(1'h1)] ?
                       reg517[(3'h6):(3'h5)] : {($signed(wire514) | $unsigned(reg555)),
                           wire515[(1'h0):(1'h0)]}));
  assign wire570 = ({(wire361 ~^ ((wire360 < reg538) ?
                               (&(8'ha0)) : (reg536 ? reg550 : (8'hac)))),
                           reg536[(1'h1):(1'h1)]} ?
                       $unsigned((^~reg543)) : $signed((reg531[(4'ha):(3'h6)] || ($unsigned(reg552) ?
                           (8'hba) : $signed(reg539)))));
  module571 #() modinst608 (wire607, clk, reg533, reg559, reg524, reg560);
  assign wire609 = ((reg528 ? $signed(reg538[(3'h5):(1'h0)]) : reg538) ?
                       wire569[(1'h1):(1'h0)] : ($signed(reg550) <<< (+($unsigned(reg517) ?
                           (reg536 || reg559) : reg541))));
  assign wire610 = (^~reg527);
  assign wire611 = (^((($unsigned(reg555) ?
                       $signed(reg523) : (-wire515)) << (~|$unsigned(reg561))) && $unsigned($unsigned($unsigned(reg538)))));
  assign wire612 = reg536;
  assign wire613 = $unsigned(reg539[(4'h9):(2'h2)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module19  (y, clk, wire23, wire22, wire21, wire20);
  output wire [(32'h72a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire23;
  input wire [(4'h8):(1'h0)] wire22;
  input wire [(5'h11):(1'h0)] wire21;
  input wire signed [(5'h12):(1'h0)] wire20;
  wire signed [(4'he):(1'h0)] wire354;
  wire signed [(5'h11):(1'h0)] wire353;
  wire signed [(2'h2):(1'h0)] wire352;
  wire signed [(3'h7):(1'h0)] wire351;
  wire signed [(4'ha):(1'h0)] wire349;
  wire [(4'hc):(1'h0)] wire174;
  wire [(5'h11):(1'h0)] wire173;
  wire [(5'h14):(1'h0)] wire102;
  wire signed [(4'ha):(1'h0)] wire101;
  wire signed [(3'h7):(1'h0)] wire84;
  wire signed [(4'h9):(1'h0)] wire83;
  reg [(4'h8):(1'h0)] reg355 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg172 = (1'h0);
  reg [(3'h6):(1'h0)] reg171 = (1'h0);
  reg [(5'h14):(1'h0)] reg168 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg167 = (1'h0);
  reg [(4'hf):(1'h0)] reg164 = (1'h0);
  reg [(4'h9):(1'h0)] reg162 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg159 = (1'h0);
  reg [(5'h12):(1'h0)] reg153 = (1'h0);
  reg [(5'h12):(1'h0)] reg158 = (1'h0);
  reg [(4'hf):(1'h0)] reg157 = (1'h0);
  reg [(2'h3):(1'h0)] reg155 = (1'h0);
  reg signed [(4'he):(1'h0)] reg154 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg147 = (1'h0);
  reg [(2'h3):(1'h0)] reg146 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg143 = (1'h0);
  reg [(4'hb):(1'h0)] reg141 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg139 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg135 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg133 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg131 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg130 = (1'h0);
  reg [(3'h6):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg127 = (1'h0);
  reg [(3'h5):(1'h0)] reg126 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg124 = (1'h0);
  reg [(2'h3):(1'h0)] reg123 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg121 = (1'h0);
  reg signed [(4'he):(1'h0)] reg119 = (1'h0);
  reg [(3'h6):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg117 = (1'h0);
  reg [(4'hd):(1'h0)] reg113 = (1'h0);
  reg [(4'h8):(1'h0)] reg112 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg111 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg108 = (1'h0);
  reg [(4'hd):(1'h0)] reg105 = (1'h0);
  reg [(4'ha):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg100 = (1'h0);
  reg [(3'h5):(1'h0)] reg99 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg98 = (1'h0);
  reg [(4'h9):(1'h0)] reg97 = (1'h0);
  reg [(4'hf):(1'h0)] reg94 = (1'h0);
  reg signed [(4'he):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg91 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg90 = (1'h0);
  reg [(5'h11):(1'h0)] reg89 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg88 = (1'h0);
  reg [(5'h14):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg81 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg76 = (1'h0);
  reg [(5'h10):(1'h0)] reg73 = (1'h0);
  reg [(4'hd):(1'h0)] reg68 = (1'h0);
  reg [(5'h14):(1'h0)] reg65 = (1'h0);
  reg [(4'hc):(1'h0)] reg63 = (1'h0);
  reg [(5'h11):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg60 = (1'h0);
  reg [(4'he):(1'h0)] reg59 = (1'h0);
  reg [(4'hd):(1'h0)] reg58 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg56 = (1'h0);
  reg [(3'h4):(1'h0)] reg54 = (1'h0);
  reg [(4'ha):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg50 = (1'h0);
  reg [(5'h12):(1'h0)] reg49 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg47 = (1'h0);
  reg [(4'h8):(1'h0)] reg45 = (1'h0);
  reg [(5'h11):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg42 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg41 = (1'h0);
  reg [(4'hc):(1'h0)] reg39 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg38 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg29 = (1'h0);
  reg [(3'h7):(1'h0)] reg24 = (1'h0);
  reg [(4'h8):(1'h0)] reg170 = (1'h0);
  reg [(4'hf):(1'h0)] reg169 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg166 = (1'h0);
  reg [(5'h12):(1'h0)] reg165 = (1'h0);
  reg [(4'ha):(1'h0)] forvar163 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg161 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg160 = (1'h0);
  reg [(5'h12):(1'h0)] reg150 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg156 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar153 = (1'h0);
  reg [(3'h6):(1'h0)] reg152 = (1'h0);
  reg [(3'h6):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar150 = (1'h0);
  reg [(3'h6):(1'h0)] reg148 = (1'h0);
  reg [(3'h6):(1'h0)] forvar145 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg142 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg137 = (1'h0);
  reg [(3'h4):(1'h0)] reg140 = (1'h0);
  reg [(3'h7):(1'h0)] reg138 = (1'h0);
  reg [(5'h10):(1'h0)] forvar137 = (1'h0);
  reg [(3'h6):(1'h0)] forvar132 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg129 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg125 = (1'h0);
  reg signed [(4'he):(1'h0)] reg122 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg120 = (1'h0);
  reg [(4'h9):(1'h0)] reg116 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg115 = (1'h0);
  reg [(3'h7):(1'h0)] reg114 = (1'h0);
  reg [(2'h2):(1'h0)] reg110 = (1'h0);
  reg [(4'hd):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg107 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg106 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar103 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar85 = (1'h0);
  reg [(4'hb):(1'h0)] reg96 = (1'h0);
  reg [(5'h12):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar92 = (1'h0);
  reg [(3'h6):(1'h0)] reg87 = (1'h0);
  reg [(4'hd):(1'h0)] reg85 = (1'h0);
  reg [(3'h6):(1'h0)] reg82 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg79 = (1'h0);
  reg [(5'h10):(1'h0)] reg78 = (1'h0);
  reg [(4'hf):(1'h0)] reg77 = (1'h0);
  reg [(2'h2):(1'h0)] reg75 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg74 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg72 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg70 = (1'h0);
  reg [(5'h12):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg67 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg66 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg64 = (1'h0);
  reg [(5'h14):(1'h0)] reg62 = (1'h0);
  reg signed [(4'he):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar55 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg53 = (1'h0);
  reg [(3'h7):(1'h0)] reg51 = (1'h0);
  reg [(5'h14):(1'h0)] reg48 = (1'h0);
  reg [(5'h11):(1'h0)] forvar24 = (1'h0);
  reg [(4'h9):(1'h0)] reg46 = (1'h0);
  reg [(3'h5):(1'h0)] reg43 = (1'h0);
  reg [(4'hb):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar37 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg35 = (1'h0);
  reg signed [(4'he):(1'h0)] reg34 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg33 = (1'h0);
  reg [(3'h4):(1'h0)] reg31 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg30 = (1'h0);
  reg [(4'h9):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg27 = (1'h0);
  reg [(3'h6):(1'h0)] reg26 = (1'h0);
  reg [(3'h6):(1'h0)] reg25 = (1'h0);
  assign y = {wire354,
                 wire353,
                 wire352,
                 wire351,
                 wire349,
                 wire174,
                 wire173,
                 wire102,
                 wire101,
                 wire84,
                 wire83,
                 reg355,
                 reg172,
                 reg171,
                 reg168,
                 reg167,
                 reg164,
                 reg162,
                 reg159,
                 reg153,
                 reg158,
                 reg157,
                 reg155,
                 reg154,
                 reg149,
                 reg147,
                 reg146,
                 reg144,
                 reg143,
                 reg141,
                 reg139,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg131,
                 reg130,
                 reg128,
                 reg127,
                 reg126,
                 reg124,
                 reg123,
                 reg121,
                 reg119,
                 reg118,
                 reg117,
                 reg113,
                 reg112,
                 reg111,
                 reg108,
                 reg105,
                 reg104,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg94,
                 reg93,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg86,
                 reg81,
                 reg76,
                 reg73,
                 reg68,
                 reg65,
                 reg63,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg56,
                 reg54,
                 reg52,
                 reg50,
                 reg49,
                 reg47,
                 reg45,
                 reg44,
                 reg42,
                 reg41,
                 reg39,
                 reg38,
                 reg36,
                 reg32,
                 reg29,
                 reg24,
                 reg170,
                 reg169,
                 reg166,
                 reg165,
                 forvar163,
                 reg161,
                 reg160,
                 reg150,
                 reg156,
                 forvar153,
                 reg152,
                 reg151,
                 forvar150,
                 reg148,
                 forvar145,
                 reg142,
                 reg137,
                 reg140,
                 reg138,
                 forvar137,
                 forvar132,
                 reg129,
                 reg125,
                 reg122,
                 reg120,
                 reg116,
                 reg115,
                 reg114,
                 reg110,
                 reg109,
                 reg107,
                 reg106,
                 forvar103,
                 reg92,
                 forvar85,
                 reg96,
                 reg95,
                 forvar92,
                 reg87,
                 reg85,
                 reg82,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg75,
                 reg74,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg67,
                 reg66,
                 reg64,
                 reg62,
                 reg57,
                 forvar55,
                 reg53,
                 reg51,
                 reg48,
                 forvar24,
                 reg46,
                 reg43,
                 reg40,
                 forvar37,
                 reg35,
                 reg34,
                 reg33,
                 reg31,
                 reg30,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire23[(4'h9):(1'h0)])
        begin
          reg24 <= ({((~|(wire20 ? wire20 : wire22)) ?
                      {$signed(wire22)} : (wire20[(5'h12):(5'h10)] ?
                          wire22[(3'h6):(3'h4)] : wire21))} ?
              (!(-(~^wire21[(4'hf):(4'ha)]))) : ({$unsigned((~wire20)),
                  {(wire21 ? wire22 : wire21),
                      $signed((8'hb0))}} ~^ ((~|{wire23, wire20}) ?
                  wire20 : (wire20 > (!wire20)))));
          if ({(wire23[(4'ha):(2'h2)] <<< reg24[(1'h0):(1'h0)])})
            begin
              reg25 = $signed(wire21);
              reg26 = ($unsigned(((((8'hb2) | wire20) || (reg24 ?
                          wire22 : wire23)) ?
                      reg24[(3'h6):(3'h6)] : reg24[(2'h2):(1'h1)])) ?
                  wire23[(4'h9):(3'h6)] : (~|wire21));
              reg27 = ((8'h9c) ? (8'ha5) : (&reg25));
              reg28 = $unsigned(wire22[(3'h4):(2'h2)]);
            end
          else
            begin
              reg29 <= (&$signed($signed($signed(reg28[(3'h4):(3'h4)]))));
              reg30 = reg25;
              reg31 = (~|(reg26[(2'h2):(2'h2)] ?
                  wire23 : $signed($unsigned($unsigned(reg27)))));
              reg32 <= wire21;
            end
          if (($signed(reg30[(2'h3):(1'h0)]) ?
              wire22[(3'h7):(3'h4)] : reg25[(2'h3):(2'h3)]))
            begin
              reg33 = {reg24,
                  ($signed($unsigned($signed(reg29))) > reg24[(3'h5):(3'h4)])};
              reg34 = reg25;
              reg35 = $signed($signed(reg27));
            end
          else
            begin
              reg36 <= $signed(($unsigned($signed(reg35[(3'h5):(3'h4)])) << ({(reg30 ?
                          reg35 : reg35)} ?
                  reg25[(2'h3):(2'h3)] : (reg28 >>> reg35))));
            end
          for (forvar37 = (1'h0); (forvar37 < (3'h4)); forvar37 = (forvar37 + (1'h1)))
            begin
              reg38 <= (~|reg24[(2'h3):(2'h2)]);
              reg39 <= $unsigned(((+$unsigned((8'hbd))) ? wire23 : wire21));
              reg40 = (~|((($unsigned(reg29) ?
                      (reg24 ? reg34 : reg39) : reg32) ?
                  reg38 : (|(wire21 ? reg31 : reg39))) + ((8'ha9) & wire21)));
            end
          if (reg26)
            begin
              reg41 <= $unsigned(reg25);
              reg42 <= (~|reg28);
            end
          else
            begin
              reg43 = (~^($unsigned({$unsigned(reg30)}) ~^ (reg35 ?
                  (reg42[(3'h5):(3'h4)] * (~^reg31)) : $unsigned($signed(wire23)))));
              reg44 <= reg42;
              reg45 <= reg42;
              reg46 = (8'hb2);
              reg47 <= $signed($signed(reg45[(3'h5):(2'h3)]));
            end
        end
      else
        begin
          for (forvar24 = (1'h0); (forvar24 < (3'h4)); forvar24 = (forvar24 + (1'h1)))
            begin
              reg25 = $unsigned(reg29);
              reg26 = $unsigned(reg38[(3'h4):(2'h2)]);
              reg27 = reg32;
            end
          if ($signed($unsigned(reg30)))
            begin
              reg29 <= (|$signed((~|reg31[(2'h3):(1'h0)])));
              reg32 <= reg38;
              reg36 <= {(8'hb1), (8'ha4)};
            end
          else
            begin
              reg28 = {$signed($signed((((8'h9c) >= forvar24) ?
                      $signed(reg28) : (|reg31)))),
                  reg44};
              reg29 <= {wire22, $unsigned({{(wire23 ? (8'hb7) : reg45)}})};
              reg30 = (^($signed($signed((forvar24 ?
                  reg46 : reg24))) < ($unsigned(reg43) ?
                  ($signed((8'had)) - (forvar24 ?
                      reg29 : reg31)) : reg38[(2'h3):(1'h1)])));
              reg31 = $unsigned({wire22[(3'h4):(2'h2)]});
            end
        end
      if ({$unsigned((~|$signed((reg24 < reg27)))), reg28})
        begin
          if (reg27)
            begin
              reg48 = (|$unsigned($unsigned($signed($unsigned(wire22)))));
              reg49 <= $unsigned((~forvar37));
              reg50 <= (reg34 ?
                  (&({$signed(reg32)} - ((|reg29) ~^ (forvar24 ^~ (8'haf))))) : $signed(($unsigned(reg39[(4'hc):(2'h3)]) ^ wire20)));
            end
          else
            begin
              reg49 <= reg33;
            end
        end
      else
        begin
          if (reg27)
            begin
              reg49 <= ($unsigned(($unsigned({reg32, reg36}) ?
                      $unsigned($unsigned(reg35)) : (^~reg40))) ?
                  $unsigned(reg26[(3'h5):(3'h5)]) : reg50[(5'h11):(5'h10)]);
              reg51 = forvar24[(1'h1):(1'h0)];
              reg52 <= forvar37[(1'h0):(1'h0)];
              reg53 = $signed(reg36);
            end
          else
            begin
              reg48 = $signed($signed(wire20[(4'ha):(4'h9)]));
              reg51 = reg39[(4'ha):(4'ha)];
            end
        end
      reg54 <= (({forvar24, $signed($unsigned(reg38))} ?
          $signed((+reg39)) : (forvar24 ?
              $unsigned($signed(reg52)) : $unsigned((reg38 >> reg52)))) == $unsigned({reg46[(3'h7):(3'h5)]}));
      for (forvar55 = (1'h0); (forvar55 < (2'h2)); forvar55 = (forvar55 + (1'h1)))
        begin
          if (forvar24[(4'hb):(3'h5)])
            begin
              reg56 <= (reg30[(4'h8):(1'h0)] ^~ forvar37[(4'hb):(4'ha)]);
            end
          else
            begin
              reg57 = $unsigned($unsigned((~|{(-reg42)})));
              reg58 <= $unsigned($unsigned($unsigned($signed($signed((8'h9c))))));
              reg59 <= $signed({($signed(reg50) ?
                      ($unsigned(reg24) ?
                          $unsigned(reg25) : {reg44}) : reg36)});
              reg60 <= ((&$unsigned((reg36 ?
                      (wire22 && (8'ha5)) : reg29[(3'h5):(1'h1)]))) ?
                  {($signed($signed(reg47)) == ((reg48 <= reg53) ?
                          $unsigned(reg38) : (+(8'ha9))))} : reg38);
              reg61 <= (((forvar55 ?
                      {(|reg49)} : ((&reg50) ? {reg31} : $unsigned(wire21))) ?
                  ((reg30 ? $signed(reg35) : reg25[(3'h4):(1'h1)]) ?
                      reg51 : ({(8'hb7)} ?
                          reg39 : $signed(reg31))) : $signed(reg45)) && $signed(reg52));
            end
        end
      if (reg25[(2'h2):(1'h1)])
        begin
          if (reg35[(3'h6):(1'h0)])
            begin
              reg62 = ($unsigned(reg52[(3'h5):(2'h3)]) && reg57);
              reg63 <= wire20;
              reg64 = (reg57 ? reg63[(3'h4):(2'h2)] : reg36[(4'h8):(1'h1)]);
            end
          else
            begin
              reg63 <= (reg63[(4'h8):(2'h3)] * (8'hae));
              reg64 = reg61;
              reg65 <= reg49[(3'h4):(1'h1)];
              reg66 = $unsigned(((~($signed(reg41) ?
                  (~(8'ha8)) : reg46[(3'h7):(3'h4)])) != {(^~(reg39 << reg57))}));
              reg67 = $signed($signed({$unsigned((reg48 <= reg38)),
                  $signed($signed(reg50))}));
            end
          if ({($unsigned(reg30[(1'h1):(1'h1)]) == ((forvar37[(4'hc):(4'h8)] ?
                      reg43[(1'h1):(1'h0)] : (reg43 ? reg27 : reg59)) ?
                  reg66 : reg64))})
            begin
              reg68 <= ($unsigned({reg29[(4'ha):(4'h9)],
                  $signed((8'hac))}) ^~ $unsigned(((~{reg36, (8'haf)}) ?
                  (((8'hb6) ^ reg38) ?
                      (^~forvar37) : $unsigned(reg56)) : (reg61[(3'h4):(1'h0)] ?
                      $unsigned(reg35) : (reg66 ? reg40 : reg27)))));
              reg69 = $unsigned(reg49[(4'ha):(4'ha)]);
            end
          else
            begin
              reg68 <= {reg64};
              reg69 = $unsigned(reg58);
              reg70 = forvar37[(4'ha):(2'h3)];
              reg71 = $signed(reg38);
              reg72 = reg28;
            end
          if (((reg34 <<< $signed((~^(wire22 ? reg68 : reg31)))) ?
              forvar55 : (reg59 || (~^((~|reg51) == (reg35 ?
                  reg69 : (7'h42)))))))
            begin
              reg73 <= (((($unsigned((8'ha6)) ? $unsigned((8'ha1)) : reg30) ?
                      reg46[(2'h2):(1'h1)] : $unsigned($signed(reg47))) ~^ reg24[(1'h1):(1'h0)]) ?
                  (~^(reg28[(3'h5):(2'h3)] ?
                      reg32 : $unsigned(reg36[(4'h8):(3'h5)]))) : (reg46 ?
                      ((~|(reg51 >= reg40)) ?
                          wire23[(4'h9):(4'h8)] : reg26) : (^$unsigned((reg27 ?
                          reg53 : reg28)))));
            end
          else
            begin
              reg74 = reg65;
            end
          reg75 = $signed($unsigned(reg45));
        end
      else
        begin
          if ((~($signed((~^((8'h9e) >>> reg53))) ~^ (reg63 - reg31[(2'h3):(2'h2)]))))
            begin
              reg63 <= (reg36 >> reg60);
              reg65 <= reg26[(2'h2):(1'h1)];
              reg68 <= reg42[(3'h5):(1'h1)];
            end
          else
            begin
              reg63 <= forvar37;
              reg65 <= (&(&$unsigned({reg51[(2'h2):(2'h2)], (8'hbc)})));
              reg66 = {reg63, $signed(reg27[(3'h6):(3'h4)])};
              reg67 = (((~&(-(~^reg47))) ?
                  (reg33[(4'he):(4'he)] ?
                      $signed((~|reg29)) : (8'hb3)) : $signed((~&{reg71,
                      (8'haa)}))) <= (~|(~&$unsigned((reg35 - reg71)))));
              reg68 <= {{(~^$signed({reg42, reg41}))},
                  $signed($signed($unsigned($unsigned((8'haa)))))};
            end
          reg73 <= (reg32[(3'h6):(1'h0)] ?
              reg40[(3'h5):(1'h0)] : reg48[(4'hb):(3'h4)]);
          reg76 <= $unsigned(($signed((reg45 ?
              {forvar24,
                  reg34} : reg67[(3'h5):(3'h4)])) >>> $unsigned($signed($unsigned((8'h9c))))));
          if ($unsigned($signed($signed((|reg68[(4'h8):(3'h6)])))))
            begin
              reg77 = ($unsigned((!(reg73 ^~ (8'h9d)))) || (+reg56[(1'h1):(1'h0)]));
              reg78 = $unsigned({reg76, $signed($signed($signed(reg49)))});
              reg79 = (reg43 <<< (reg25[(2'h2):(2'h2)] ~^ reg60));
              reg80 = ((8'ha2) >= $unsigned((8'ha2)));
            end
          else
            begin
              reg81 <= $signed((~&reg34));
              reg82 = (^~reg62[(3'h5):(2'h2)]);
            end
        end
    end
  assign wire83 = (~&(reg24[(3'h6):(1'h1)] && $unsigned($signed({reg47}))));
  assign wire84 = $unsigned((wire20 ^ $signed((~|$unsigned(reg81)))));
  always
    @(posedge clk) begin
      if (((~(reg58[(4'ha):(1'h1)] ?
              reg50[(4'h8):(1'h1)] : (~$unsigned(reg68)))) ?
          {$signed(((|reg41) & (reg32 ?
                  reg81 : reg45)))} : $unsigned(($signed((8'hb5)) ?
              (!$unsigned(wire23)) : (~(wire20 ? wire21 : wire23))))))
        begin
          if ((~|((reg50 || ((reg65 ? reg52 : reg44) ?
                  reg49[(5'h10):(4'hd)] : (|reg59))) ?
              (((~^reg24) ?
                  $unsigned(reg76) : $signed(reg73)) - $signed($unsigned(reg68))) : reg59)))
            begin
              reg85 = (reg49 <<< (({$unsigned(wire22), wire83[(3'h6):(1'h0)]} ?
                  {reg73[(4'hb):(2'h3)],
                      $unsigned((8'ha0))} : (8'hae)) <= reg73[(4'he):(2'h2)]));
              reg86 <= (^reg44);
              reg87 = reg52[(3'h5):(2'h2)];
            end
          else
            begin
              reg86 <= (^~$unsigned((^~$unsigned((~|wire84)))));
              reg88 <= $unsigned((+$signed(reg45[(3'h6):(3'h4)])));
              reg89 <= ($signed($signed($signed(((8'hbc) && reg50)))) ?
                  {$signed($signed((~&reg59)))} : {reg39});
              reg90 <= $unsigned($signed(reg49));
              reg91 <= $unsigned({$signed((&(reg52 ? reg73 : reg38))),
                  (($signed((8'hb6)) < {reg41, reg86}) ^ (7'h40))});
            end
          for (forvar92 = (1'h0); (forvar92 < (3'h4)); forvar92 = (forvar92 + (1'h1)))
            begin
              reg93 <= (reg88[(2'h3):(1'h0)] >= $unsigned({((reg61 ^ wire23) != (~reg68)),
                  reg81}));
            end
          if ((7'h44))
            begin
              reg94 <= $unsigned($signed((reg87[(3'h5):(3'h5)] <<< reg36)));
            end
          else
            begin
              reg95 = ((!reg89[(3'h4):(2'h3)]) >>> {wire20});
              reg96 = $signed((-$signed((((8'hbf) ?
                  reg88 : reg87) >>> (reg85 >= (8'hab))))));
              reg97 <= (!((({(8'h9e), (8'hac)} > wire83) ?
                  (^~(reg59 * reg86)) : $signed((reg38 <<< reg29))) - reg88[(3'h5):(2'h3)]));
              reg98 <= (~&(reg63 ?
                  ((~(-reg42)) ? (8'hae) : (&wire84)) : (reg73 ?
                      {{reg94}, wire21[(4'hf):(1'h1)]} : ((~^reg58) ?
                          (~&(8'hbe)) : (reg68 ? reg44 : wire21)))));
              reg99 <= $unsigned((reg39[(4'h9):(4'h8)] ?
                  (reg39 ^~ reg81[(1'h0):(1'h0)]) : (-reg42[(1'h1):(1'h1)])));
            end
          reg100 <= reg38;
        end
      else
        begin
          for (forvar85 = (1'h0); (forvar85 < (1'h0)); forvar85 = (forvar85 + (1'h1)))
            begin
              reg86 <= (7'h44);
              reg87 = wire84;
              reg92 = (-$unsigned(reg88));
              reg93 <= (-(^~reg61[(3'h4):(2'h2)]));
              reg94 <= (reg91 ?
                  ($signed((reg85[(3'h4):(1'h0)] == reg87)) < ((~((8'h9d) ^ reg38)) | (&$signed(wire84)))) : ((-((8'hb3) ?
                          (8'hbe) : reg24[(3'h7):(3'h7)])) ?
                      (~^reg59) : $signed(({reg29} <= reg68[(3'h4):(2'h3)]))));
            end
        end
    end
  assign wire101 = $unsigned(reg32);
  assign wire102 = reg99[(3'h4):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar103 = (1'h0); (forvar103 < (2'h2)); forvar103 = (forvar103 + (1'h1)))
        begin
          if ($unsigned($unsigned((reg73[(4'he):(3'h5)] ?
              reg94[(4'h8):(3'h7)] : $signed((reg47 >> (8'hb9)))))))
            begin
              reg104 <= reg58[(4'ha):(4'h8)];
              reg105 <= {(|$signed(((reg47 ?
                      reg54 : wire101) & (reg86 ^ wire22))))};
            end
          else
            begin
              reg106 = $unsigned(reg58[(1'h0):(1'h0)]);
              reg107 = $signed(reg42);
              reg108 <= ($unsigned((^~(((8'ha8) <<< wire83) ?
                      (&reg65) : reg105[(4'hd):(3'h7)]))) ?
                  reg89[(5'h10):(3'h5)] : reg50[(5'h12):(1'h0)]);
            end
          reg109 = $signed(({(7'h44),
              reg107[(3'h4):(1'h1)]} >>> reg93[(4'hb):(4'h8)]));
          reg110 = $signed($signed(((((8'ha2) ? reg107 : reg60) ?
                  reg56[(1'h1):(1'h1)] : reg54) ?
              (wire83[(1'h1):(1'h1)] ?
                  (wire22 & reg39) : $signed((8'hb3))) : (-(reg81 ?
                  reg47 : (8'ha4))))));
          reg111 <= (|$signed($signed({((7'h43) < reg44),
              (reg110 <<< (8'hb3))})));
          if ($unsigned({(reg90[(2'h2):(2'h2)] ?
                  $signed((reg68 ?
                      (8'haf) : reg45)) : $unsigned($signed(reg104)))}))
            begin
              reg112 <= reg56;
              reg113 <= $signed(reg88[(2'h2):(1'h0)]);
            end
          else
            begin
              reg114 = (reg106 >= $unsigned((8'h9f)));
              reg115 = ($signed({($signed(reg91) >> (+(8'haa))),
                  reg38[(2'h3):(1'h1)]}) ^~ $signed($unsigned((~&((8'h9e) ?
                  reg112 : reg47)))));
              reg116 = (reg114[(2'h2):(1'h0)] << (~|reg38[(2'h2):(1'h0)]));
            end
        end
      reg117 <= reg91[(3'h7):(1'h1)];
      if (reg45)
        begin
          reg118 <= $signed({reg108, $signed(reg114)});
          if ($unsigned(wire22[(2'h3):(2'h2)]))
            begin
              reg119 <= reg105[(4'h9):(2'h3)];
              reg120 = ((~|((-{reg89,
                  reg58}) < $unsigned($unsigned((8'hbf))))) ~^ $signed(($unsigned((~&reg89)) < reg98[(4'hd):(3'h7)])));
              reg121 <= (((((wire84 == reg38) ? reg112 : reg104) & reg97) ?
                  (~^reg91[(1'h0):(1'h0)]) : {(reg89[(5'h11):(3'h6)] || (reg107 - reg108))}) > (~&$signed({wire20,
                  $unsigned(reg39)})));
              reg122 = {($signed({$unsigned(reg88)}) >= $unsigned(((wire84 ?
                          reg113 : (8'hbe)) ?
                      {reg81} : (~wire102)))),
                  (|$unsigned(wire83[(3'h5):(2'h3)]))};
            end
          else
            begin
              reg120 = $unsigned(wire21);
              reg122 = $signed(reg91);
              reg123 <= {($unsigned(reg76[(1'h0):(1'h0)]) ?
                      {$unsigned(reg29[(2'h3):(2'h2)])} : (!{(reg105 > reg116),
                          (wire102 ? reg108 : wire102)})),
                  (8'hb2)};
              reg124 <= wire22[(1'h0):(1'h0)];
              reg125 = ({wire22[(1'h0):(1'h0)], reg54} ?
                  (8'hbf) : reg111[(4'hc):(1'h0)]);
            end
        end
      else
        begin
          if (reg117[(3'h5):(1'h1)])
            begin
              reg118 <= (($signed(reg118) ^~ reg65) ?
                  $unsigned({$unsigned($unsigned((7'h43)))}) : reg91[(1'h1):(1'h0)]);
              reg119 <= $unsigned($signed((reg73 >>> reg54)));
            end
          else
            begin
              reg120 = reg118[(2'h2):(1'h1)];
              reg122 = reg120;
            end
          if ($unsigned(reg41))
            begin
              reg123 <= reg41[(2'h3):(2'h3)];
              reg124 <= $signed(reg125[(1'h0):(1'h0)]);
              reg125 = $unsigned(({($unsigned(reg88) ?
                          $unsigned(reg44) : ((8'hbc) <= reg107)),
                      $unsigned((~reg98))} ?
                  ((-((7'h40) ?
                      reg104 : reg58)) && reg68[(4'h9):(4'h8)]) : $unsigned((reg110 << reg24))));
            end
          else
            begin
              reg125 = (|(({$unsigned((8'h9f)), (reg91 + reg119)} ?
                      (~&$unsigned(forvar103)) : $signed((reg36 <= reg111))) ?
                  $unsigned(reg97) : $unsigned({reg45[(3'h7):(2'h3)]})));
              reg126 <= $unsigned(reg54);
            end
          if ($signed((~reg68[(3'h7):(2'h3)])))
            begin
              reg127 <= {reg56[(2'h3):(2'h3)]};
              reg128 <= {reg38,
                  {($unsigned({reg81, wire20}) ?
                          reg91 : {(reg63 ? (7'h40) : (8'h9f))})}};
            end
          else
            begin
              reg129 = (wire23 >>> reg112);
              reg130 <= $signed(reg104);
              reg131 <= $signed(($signed((8'h9f)) == (reg42[(1'h0):(1'h0)] != reg81[(1'h0):(1'h0)])));
            end
          for (forvar132 = (1'h0); (forvar132 < (1'h0)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 <= {$signed((($signed((8'ha5)) ?
                          wire23[(2'h3):(2'h2)] : $signed(reg114)) ?
                      reg127 : $unsigned((wire102 + reg120)))),
                  {reg76, wire102[(2'h2):(1'h0)]}};
            end
          if ({$signed(($signed(reg122) ?
                  reg88 : $unsigned($unsigned(wire101)))),
              $unsigned($signed(reg111[(4'h8):(1'h1)]))})
            begin
              reg134 <= (({((8'hb7) + reg93)} ~^ ((~|reg36[(4'h9):(3'h5)]) ?
                  $unsigned((reg129 ?
                      reg129 : reg90)) : reg106)) && reg113[(3'h4):(1'h0)]);
            end
          else
            begin
              reg134 <= $unsigned((~^{((reg38 ^~ reg49) < wire23), reg93}));
              reg135 <= (8'hb2);
              reg136 <= $unsigned($unsigned(reg39[(1'h0):(1'h0)]));
            end
        end
      if ((((reg122[(4'hd):(1'h0)] > ((^(8'ha3)) ?
          $signed(forvar103) : reg60)) - reg116) >> (^$unsigned($unsigned(((8'hb2) | reg112))))))
        begin
          for (forvar137 = (1'h0); (forvar137 < (1'h0)); forvar137 = (forvar137 + (1'h1)))
            begin
              reg138 = ({reg81, $signed(reg73)} ?
                  wire101[(4'ha):(2'h3)] : $signed(((~&reg136[(4'hb):(2'h2)]) ?
                      ($unsigned((7'h43)) ^~ reg61) : ((reg45 << reg65) | (-reg97)))));
              reg139 <= reg118;
              reg140 = {$unsigned($signed((~reg128[(3'h6):(3'h6)])))};
              reg141 <= (+$unsigned(reg61));
            end
        end
      else
        begin
          reg137 = (~|$unsigned(reg65[(4'hf):(1'h0)]));
          if ($unsigned(wire20[(1'h0):(1'h0)]))
            begin
              reg139 <= (~&$signed((reg121[(3'h4):(2'h2)] >= (((8'hb6) ?
                  reg135 : reg54) >>> reg88[(3'h6):(2'h3)]))));
              reg140 = reg123[(1'h1):(1'h0)];
              reg142 = (+{(~($unsigned(reg32) ?
                      (reg117 ? reg88 : reg68) : (reg90 != forvar137)))});
            end
          else
            begin
              reg138 = reg39[(1'h1):(1'h0)];
              reg140 = $signed(reg52);
              reg141 <= (^reg54);
              reg143 <= $signed(((!(8'hae)) + $signed((&{reg36}))));
              reg144 <= (reg111[(3'h6):(1'h0)] ^~ {($signed((reg91 ?
                          reg121 : reg65)) ?
                      (-(reg120 ? (8'ha0) : reg65)) : reg98[(3'h4):(2'h3)])});
            end
          for (forvar145 = (1'h0); (forvar145 < (3'h4)); forvar145 = (forvar145 + (1'h1)))
            begin
              reg146 <= $unsigned(reg76);
              reg147 <= (|(^~reg108));
              reg148 = (-$signed($unsigned(wire102)));
            end
          reg149 <= (wire23[(1'h0):(1'h0)] ?
              (^(({reg124} ?
                  (reg73 ? reg120 : (8'h9e)) : ((8'hbb) ?
                      reg60 : reg141)) > $unsigned((&(8'ha3))))) : ((reg124[(4'h8):(1'h1)] ?
                      (reg109 ? reg94 : (8'ha7)) : $unsigned(((8'hb7) ?
                          reg140 : reg41))) ?
                  ((reg127 || reg119[(3'h6):(3'h4)]) ?
                      (reg125[(3'h5):(1'h1)] ?
                          reg118[(3'h4):(2'h2)] : (reg148 ?
                              reg138 : reg89)) : {$unsigned(reg115),
                          $unsigned(reg44)}) : $unsigned((reg29 ?
                      $unsigned(reg52) : (reg107 ^~ wire21)))));
        end
      if ($unsigned((reg42 ?
          reg91[(3'h4):(2'h3)] : (^(&reg136[(2'h2):(1'h0)])))))
        begin
          for (forvar150 = (1'h0); (forvar150 < (2'h2)); forvar150 = (forvar150 + (1'h1)))
            begin
              reg151 = reg124;
            end
          reg152 = reg122;
          for (forvar153 = (1'h0); (forvar153 < (3'h4)); forvar153 = (forvar153 + (1'h1)))
            begin
              reg154 <= wire101[(1'h1):(1'h0)];
            end
          if (reg126[(3'h5):(3'h5)])
            begin
              reg155 <= (^forvar153);
              reg156 = reg94;
              reg157 <= (~$unsigned(reg127));
              reg158 <= (reg110[(1'h0):(1'h0)] ?
                  $unsigned(reg154) : reg135[(5'h10):(4'hd)]);
            end
          else
            begin
              reg156 = reg117[(4'h9):(4'h8)];
            end
        end
      else
        begin
          if ($unsigned(({$signed(reg59)} ^ (&forvar132))))
            begin
              reg150 = reg105;
              reg151 = reg114;
              reg153 <= reg86;
              reg156 = $signed($unsigned({(^reg61[(4'h8):(3'h5)])}));
            end
          else
            begin
              reg150 = (~^$signed(reg124[(3'h4):(3'h4)]));
              reg153 <= (~^((reg154 ?
                      ((+reg113) >= ((8'h9d) != reg29)) : (^reg136)) ?
                  reg49[(3'h4):(2'h2)] : $unsigned({reg126[(3'h4):(3'h4)],
                      reg119[(4'hd):(1'h1)]})));
              reg154 <= reg68;
              reg156 = ((&reg116[(1'h0):(1'h0)]) <<< (~|$signed(((wire84 >= reg116) & (reg65 ^~ wire20)))));
            end
          if (reg138[(3'h5):(2'h2)])
            begin
              reg157 <= ($signed(reg91[(3'h6):(3'h5)]) && wire21[(2'h3):(2'h3)]);
              reg158 <= (8'hb8);
              reg159 <= {reg56, reg52};
              reg160 = $signed(reg116);
            end
          else
            begin
              reg160 = (reg98 ?
                  reg98[(3'h7):(3'h7)] : $unsigned($unsigned(($signed(reg41) & ((8'hbc) ?
                      (8'had) : reg93)))));
              reg161 = reg109;
            end
          reg162 <= (({{((8'hb6) >>> reg118), (reg150 | reg157)},
                  reg65} ^~ $signed($signed($unsigned(reg47)))) ?
              ({$unsigned(reg112), reg159[(3'h5):(3'h5)]} ?
                  {$signed((reg49 << reg47)),
                      (reg159[(4'ha):(1'h0)] != (reg115 ?
                          reg88 : reg68))} : reg38[(2'h2):(1'h1)]) : ($unsigned((^(~^reg89))) ?
                  (~|(~reg63)) : reg29[(3'h5):(3'h4)]));
          for (forvar163 = (1'h0); (forvar163 < (2'h3)); forvar163 = (forvar163 + (1'h1)))
            begin
              reg164 <= reg162;
            end
          if ($unsigned(((~^reg133) * reg157)))
            begin
              reg165 = reg128[(3'h4):(2'h3)];
              reg166 = $unsigned((!(!wire84)));
              reg167 <= $signed($signed((reg155 ?
                  reg137[(4'ha):(4'ha)] : reg150[(4'hf):(4'hb)])));
              reg168 <= (reg127[(4'he):(4'hc)] ?
                  $signed($unsigned(reg41[(3'h5):(2'h2)])) : (&(~&(reg138 < (8'hb4)))));
              reg169 = {reg134, (~&(^reg130[(2'h2):(1'h0)]))};
            end
          else
            begin
              reg167 <= $unsigned((~wire101[(3'h5):(3'h4)]));
              reg169 = $signed(((((reg122 < reg89) ?
                  ((7'h41) << reg38) : {reg143,
                      reg136}) < reg97[(4'h8):(1'h1)]) != reg162));
              reg170 = (reg47 != (reg91 ?
                  forvar137 : {reg60, $signed(reg148[(3'h5):(3'h5)])}));
              reg171 <= (|$signed($signed($unsigned(((8'hb2) << reg99)))));
              reg172 <= $signed($unsigned(reg93[(4'h8):(3'h5)]));
            end
        end
    end
  assign wire173 = $unsigned(($unsigned((~&{reg134, reg127})) ?
                       (~^$signed($unsigned((7'h43)))) : $unsigned(((!reg154) ^~ (!(8'hbf))))));
  assign wire174 = reg153[(5'h11):(4'hd)];
  module175 #() modinst350 (wire349, clk, wire102, reg111, reg61, wire173);
  assign wire351 = $unsigned(reg154);
  assign wire352 = (~^((8'ha5) ?
                       (reg117 > {reg159[(4'h9):(3'h7)],
                           $signed(reg105)}) : $unsigned((reg76 + $signed(reg157)))));
  assign wire353 = reg123;
  assign wire354 = $signed(reg136);
  always
    @(posedge clk) begin
      reg355 <= $signed(reg119[(4'he):(2'h2)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4  (y, clk, wire9, wire8, wire7, wire6, wire5);
  output wire [(32'h45):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire9;
  input wire [(2'h3):(1'h0)] wire8;
  input wire signed [(5'h11):(1'h0)] wire7;
  input wire signed [(3'h6):(1'h0)] wire6;
  input wire signed [(4'hc):(1'h0)] wire5;
  wire signed [(3'h4):(1'h0)] wire16;
  wire [(4'h9):(1'h0)] wire15;
  wire [(4'ha):(1'h0)] wire14;
  wire signed [(4'hd):(1'h0)] wire13;
  wire signed [(4'ha):(1'h0)] wire12;
  wire [(4'ha):(1'h0)] wire11;
  wire [(4'hc):(1'h0)] wire10;
  assign y = {wire16, wire15, wire14, wire13, wire12, wire11, wire10, (1'h0)};
  assign wire10 = $unsigned({wire8[(1'h0):(1'h0)],
                      $signed(((wire9 > wire8) >> wire6[(2'h2):(1'h1)]))});
  assign wire11 = wire6;
  assign wire12 = $signed($signed(wire8[(1'h0):(1'h0)]));
  assign wire13 = ($unsigned($unsigned({wire9[(2'h3):(1'h0)],
                      $unsigned((7'h42))})) - (wire11 ?
                      ($unsigned(wire12) * wire10) : (~^((wire10 ?
                              wire5 : wire5) ?
                          $signed(wire11) : $unsigned(wire12)))));
  assign wire14 = $signed(wire7[(4'ha):(4'ha)]);
  assign wire15 = (+wire7[(2'h3):(2'h2)]);
  assign wire16 = wire15;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module175  (y, clk, wire179, wire178, wire177, wire176);
  output wire [(32'h7b9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire179;
  input wire signed [(4'hb):(1'h0)] wire178;
  input wire [(5'h11):(1'h0)] wire177;
  input wire [(5'h11):(1'h0)] wire176;
  wire signed [(4'ha):(1'h0)] wire348;
  wire signed [(5'h10):(1'h0)] wire347;
  wire signed [(4'hf):(1'h0)] wire346;
  wire [(2'h2):(1'h0)] wire309;
  wire signed [(4'hc):(1'h0)] wire308;
  wire [(4'h9):(1'h0)] wire288;
  wire signed [(4'hc):(1'h0)] wire287;
  wire signed [(4'hd):(1'h0)] wire286;
  wire [(5'h12):(1'h0)] wire185;
  wire [(4'hb):(1'h0)] wire184;
  wire signed [(2'h2):(1'h0)] wire183;
  wire [(5'h14):(1'h0)] wire182;
  wire [(2'h2):(1'h0)] wire181;
  wire [(4'hc):(1'h0)] wire180;
  reg [(5'h14):(1'h0)] reg344 = (1'h0);
  reg [(4'ha):(1'h0)] reg342 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg340 = (1'h0);
  reg signed [(4'he):(1'h0)] reg339 = (1'h0);
  reg [(5'h11):(1'h0)] reg335 = (1'h0);
  reg [(3'h5):(1'h0)] reg333 = (1'h0);
  reg [(3'h6):(1'h0)] reg332 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg331 = (1'h0);
  reg [(5'h11):(1'h0)] reg330 = (1'h0);
  reg [(3'h5):(1'h0)] reg324 = (1'h0);
  reg [(2'h3):(1'h0)] reg323 = (1'h0);
  reg [(5'h14):(1'h0)] reg322 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg320 = (1'h0);
  reg [(5'h13):(1'h0)] reg319 = (1'h0);
  reg [(3'h7):(1'h0)] reg315 = (1'h0);
  reg [(3'h4):(1'h0)] reg314 = (1'h0);
  reg [(5'h13):(1'h0)] reg313 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg307 = (1'h0);
  reg [(4'hb):(1'h0)] reg306 = (1'h0);
  reg [(4'ha):(1'h0)] reg303 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg302 = (1'h0);
  reg [(5'h13):(1'h0)] reg300 = (1'h0);
  reg [(4'he):(1'h0)] reg299 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg298 = (1'h0);
  reg [(3'h5):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg293 = (1'h0);
  reg [(5'h15):(1'h0)] reg292 = (1'h0);
  reg [(3'h5):(1'h0)] reg274 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg285 = (1'h0);
  reg [(2'h3):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg283 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg277 = (1'h0);
  reg [(4'ha):(1'h0)] reg276 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg267 = (1'h0);
  reg [(4'hb):(1'h0)] reg272 = (1'h0);
  reg [(4'hc):(1'h0)] reg271 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg269 = (1'h0);
  reg [(4'ha):(1'h0)] reg268 = (1'h0);
  reg [(4'ha):(1'h0)] reg265 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg262 = (1'h0);
  reg [(4'hc):(1'h0)] reg261 = (1'h0);
  reg [(3'h4):(1'h0)] reg260 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg259 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg258 = (1'h0);
  reg [(5'h10):(1'h0)] reg256 = (1'h0);
  reg [(3'h7):(1'h0)] reg253 = (1'h0);
  reg [(4'h8):(1'h0)] reg250 = (1'h0);
  reg [(4'h8):(1'h0)] reg249 = (1'h0);
  reg [(3'h4):(1'h0)] reg247 = (1'h0);
  reg [(3'h6):(1'h0)] reg245 = (1'h0);
  reg [(4'hc):(1'h0)] reg244 = (1'h0);
  reg [(4'hf):(1'h0)] reg243 = (1'h0);
  reg [(4'ha):(1'h0)] reg240 = (1'h0);
  reg [(4'he):(1'h0)] reg237 = (1'h0);
  reg [(5'h15):(1'h0)] reg236 = (1'h0);
  reg [(2'h2):(1'h0)] reg235 = (1'h0);
  reg [(4'hc):(1'h0)] reg233 = (1'h0);
  reg [(3'h4):(1'h0)] reg231 = (1'h0);
  reg [(4'hd):(1'h0)] reg230 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg229 = (1'h0);
  reg [(5'h12):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg226 = (1'h0);
  reg [(5'h10):(1'h0)] reg223 = (1'h0);
  reg [(5'h11):(1'h0)] reg222 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg220 = (1'h0);
  reg [(4'he):(1'h0)] reg216 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg215 = (1'h0);
  reg [(4'ha):(1'h0)] reg213 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg211 = (1'h0);
  reg [(5'h12):(1'h0)] reg210 = (1'h0);
  reg [(4'ha):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg207 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg199 = (1'h0);
  reg [(5'h11):(1'h0)] reg193 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg191 = (1'h0);
  reg [(4'h9):(1'h0)] reg190 = (1'h0);
  reg signed [(4'he):(1'h0)] reg188 = (1'h0);
  reg [(4'hf):(1'h0)] reg186 = (1'h0);
  reg [(5'h11):(1'h0)] reg345 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg343 = (1'h0);
  reg [(4'h9):(1'h0)] forvar338 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar337 = (1'h0);
  reg [(4'h9):(1'h0)] reg336 = (1'h0);
  reg [(2'h2):(1'h0)] reg334 = (1'h0);
  reg [(4'hc):(1'h0)] reg329 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar328 = (1'h0);
  reg [(4'hd):(1'h0)] reg327 = (1'h0);
  reg [(4'hd):(1'h0)] reg326 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg325 = (1'h0);
  reg [(3'h4):(1'h0)] reg321 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg318 = (1'h0);
  reg [(4'ha):(1'h0)] reg317 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar316 = (1'h0);
  reg [(5'h13):(1'h0)] reg312 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar311 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar310 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar305 = (1'h0);
  reg [(4'hf):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg301 = (1'h0);
  reg [(5'h13):(1'h0)] reg296 = (1'h0);
  reg [(4'ha):(1'h0)] forvar295 = (1'h0);
  reg [(4'hb):(1'h0)] reg291 = (1'h0);
  reg [(4'hb):(1'h0)] forvar290 = (1'h0);
  reg [(5'h12):(1'h0)] reg289 = (1'h0);
  reg [(2'h3):(1'h0)] reg282 = (1'h0);
  reg [(4'hf):(1'h0)] reg281 = (1'h0);
  reg [(4'hc):(1'h0)] forvar280 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg279 = (1'h0);
  reg [(5'h13):(1'h0)] reg278 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg275 = (1'h0);
  reg [(5'h15):(1'h0)] forvar274 = (1'h0);
  reg [(3'h5):(1'h0)] forvar268 = (1'h0);
  reg [(3'h4):(1'h0)] reg273 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg270 = (1'h0);
  reg [(5'h13):(1'h0)] forvar267 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg264 = (1'h0);
  reg [(5'h13):(1'h0)] reg263 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg255 = (1'h0);
  reg [(3'h7):(1'h0)] reg254 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg252 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg251 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg248 = (1'h0);
  reg [(5'h12):(1'h0)] forvar246 = (1'h0);
  reg [(3'h7):(1'h0)] reg242 = (1'h0);
  reg [(2'h3):(1'h0)] reg241 = (1'h0);
  reg [(5'h10):(1'h0)] reg239 = (1'h0);
  reg [(4'hb):(1'h0)] forvar231 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg238 = (1'h0);
  reg [(4'hf):(1'h0)] reg234 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg227 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg225 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg224 = (1'h0);
  reg [(5'h13):(1'h0)] reg219 = (1'h0);
  reg [(5'h12):(1'h0)] forvar218 = (1'h0);
  reg [(5'h15):(1'h0)] reg217 = (1'h0);
  reg [(3'h4):(1'h0)] reg214 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg212 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg209 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar186 = (1'h0);
  reg [(3'h7):(1'h0)] reg206 = (1'h0);
  reg [(2'h2):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg204 = (1'h0);
  reg [(3'h5):(1'h0)] forvar202 = (1'h0);
  reg signed [(4'he):(1'h0)] reg201 = (1'h0);
  reg [(4'hc):(1'h0)] reg200 = (1'h0);
  reg [(4'hd):(1'h0)] reg198 = (1'h0);
  reg [(4'h9):(1'h0)] reg197 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg196 = (1'h0);
  reg [(4'ha):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg194 = (1'h0);
  reg [(5'h12):(1'h0)] reg192 = (1'h0);
  reg [(4'h8):(1'h0)] reg189 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg187 = (1'h0);
  assign y = {wire348,
                 wire347,
                 wire346,
                 wire309,
                 wire308,
                 wire288,
                 wire287,
                 wire286,
                 wire185,
                 wire184,
                 wire183,
                 wire182,
                 wire181,
                 wire180,
                 reg344,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg335,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg324,
                 reg323,
                 reg322,
                 reg320,
                 reg319,
                 reg315,
                 reg314,
                 reg313,
                 reg307,
                 reg306,
                 reg303,
                 reg302,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg294,
                 reg293,
                 reg292,
                 reg274,
                 reg285,
                 reg284,
                 reg283,
                 reg277,
                 reg276,
                 reg267,
                 reg272,
                 reg271,
                 reg269,
                 reg268,
                 reg265,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg256,
                 reg253,
                 reg250,
                 reg249,
                 reg247,
                 reg245,
                 reg244,
                 reg243,
                 reg240,
                 reg237,
                 reg236,
                 reg235,
                 reg233,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg226,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg216,
                 reg215,
                 reg213,
                 reg211,
                 reg210,
                 reg202,
                 reg208,
                 reg207,
                 reg203,
                 reg199,
                 reg193,
                 reg191,
                 reg190,
                 reg188,
                 reg186,
                 reg345,
                 reg343,
                 forvar338,
                 forvar337,
                 reg336,
                 reg334,
                 reg329,
                 forvar328,
                 reg327,
                 reg326,
                 reg325,
                 reg321,
                 reg318,
                 reg317,
                 forvar316,
                 reg312,
                 forvar311,
                 forvar310,
                 forvar305,
                 reg304,
                 reg301,
                 reg296,
                 forvar295,
                 reg291,
                 forvar290,
                 reg289,
                 reg282,
                 reg281,
                 forvar280,
                 reg279,
                 reg278,
                 reg275,
                 forvar274,
                 forvar268,
                 reg273,
                 reg270,
                 forvar267,
                 reg266,
                 reg264,
                 reg263,
                 reg257,
                 reg255,
                 reg254,
                 reg252,
                 reg251,
                 reg248,
                 forvar246,
                 reg242,
                 reg241,
                 reg239,
                 forvar231,
                 reg238,
                 reg234,
                 reg232,
                 reg227,
                 reg225,
                 reg224,
                 reg219,
                 forvar218,
                 reg217,
                 reg214,
                 reg212,
                 reg209,
                 forvar186,
                 reg206,
                 reg205,
                 reg204,
                 forvar202,
                 reg201,
                 reg200,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg192,
                 reg189,
                 reg187,
                 (1'h0)};
  assign wire180 = wire177[(3'h7):(3'h6)];
  assign wire181 = ($signed($signed(wire177[(3'h7):(2'h2)])) ?
                       (~|{(^~$signed(wire180))}) : (wire179[(4'ha):(2'h2)] ?
                           $signed(((&wire176) && {wire177,
                               wire180})) : wire179));
  assign wire182 = (|(wire181 ^~ {wire177, {(wire177 + wire177)}}));
  assign wire183 = wire176[(1'h0):(1'h0)];
  assign wire184 = wire182;
  assign wire185 = (~&wire180[(3'h4):(3'h4)]);
  always
    @(posedge clk) begin
      if ((^$unsigned($signed(wire182[(1'h1):(1'h1)]))))
        begin
          if (wire178)
            begin
              reg186 <= (8'ha6);
              reg187 = wire183;
              reg188 <= (^((~|$signed($unsigned(wire178))) ?
                  $unsigned(wire181[(1'h1):(1'h0)]) : reg187[(2'h3):(1'h1)]));
              reg189 = (^wire178);
            end
          else
            begin
              reg187 = $signed($unsigned(wire177[(4'hf):(1'h1)]));
              reg188 <= wire181[(1'h0):(1'h0)];
              reg190 <= $unsigned((|wire184[(4'h9):(3'h6)]));
              reg191 <= (|$signed(wire179));
              reg192 = (7'h41);
            end
          if (reg190)
            begin
              reg193 <= (|$unsigned((reg188[(4'ha):(3'h4)] ?
                  $unsigned(wire185) : {(wire182 | wire185)})));
            end
          else
            begin
              reg193 <= ((~^(reg189 ?
                  {wire176,
                      reg192} : (~^$signed(wire181)))) | reg188[(4'he):(1'h1)]);
              reg194 = (wire177 ?
                  $signed($signed(((~&wire178) ?
                      wire183[(1'h0):(1'h0)] : ((8'hbf) ?
                          wire179 : (8'hb2))))) : {((wire176 ?
                          (8'hbb) : $unsigned(reg188)) & wire177),
                      {((wire176 | reg190) ?
                              wire182[(3'h5):(1'h0)] : $signed(reg190)),
                          $unsigned((~reg192))}});
              reg195 = (((~&{(^~wire179)}) || $signed(((&wire182) ?
                  (wire180 ?
                      wire180 : wire184) : ((8'ha0) >= wire176)))) | reg188);
              reg196 = $signed((reg195[(1'h0):(1'h0)] ?
                  ((^$unsigned((8'ha4))) ?
                      ($unsigned(wire177) - (reg191 ?
                          reg190 : reg195)) : (reg195[(3'h6):(1'h0)] ?
                          reg194[(4'h9):(3'h6)] : $unsigned(wire176))) : ({{wire184,
                          reg193},
                      (wire178 ?
                          wire182 : (8'hba))} && reg189[(1'h0):(1'h0)])));
            end
          if ($unsigned(wire179))
            begin
              reg197 = (({wire176} ?
                      (+(!(8'hbc))) : $unsigned($unsigned(wire180))) ?
                  $unsigned($signed(wire181)) : (!{wire184}));
              reg198 = wire182;
              reg199 <= ($unsigned((wire185[(5'h11):(1'h1)] ?
                      wire176[(1'h1):(1'h0)] : $signed({(8'h9c)}))) ?
                  ((^{$unsigned(wire180), (reg190 ? (8'ha2) : reg190)}) ?
                      $unsigned($signed($unsigned(wire185))) : ((|reg196[(2'h3):(2'h2)]) >= {$signed(wire183)})) : $signed($unsigned((reg188[(4'hb):(1'h0)] != reg194))));
              reg200 = (wire180 ? (8'h9e) : wire181[(1'h1):(1'h0)]);
              reg201 = $unsigned($signed((($unsigned(wire183) ?
                      (reg190 ? reg189 : (8'hb3)) : $signed((8'hb0))) ?
                  $signed((reg186 || reg191)) : $unsigned(wire178[(3'h7):(2'h3)]))));
            end
          else
            begin
              reg197 = reg196[(1'h0):(1'h0)];
              reg198 = ({(|$signed(reg190)), wire185[(1'h0):(1'h0)]} ?
                  (reg199 >= $unsigned($signed((reg192 * reg192)))) : ($signed((~|(wire180 ?
                          (8'hbf) : reg201))) ?
                      {wire183[(1'h0):(1'h0)], reg191} : reg197));
              reg200 = (((~^reg188) >> (($unsigned(wire183) ?
                      (wire181 ?
                          (8'ha0) : reg192) : reg199[(3'h7):(3'h5)]) * reg191)) ?
                  wire176[(4'hf):(4'hd)] : {reg193});
            end
          for (forvar202 = (1'h0); (forvar202 < (1'h1)); forvar202 = (forvar202 + (1'h1)))
            begin
              reg203 <= wire177[(4'h8):(4'h8)];
              reg204 = (!(!$unsigned(($unsigned((7'h41)) ?
                  (~&reg197) : $signed(reg188)))));
              reg205 = $unsigned($unsigned({(~^$signed(reg193)),
                  (&(reg198 ? reg203 : wire184))}));
              reg206 = $signed($unsigned(reg188[(4'h8):(2'h2)]));
              reg207 <= $unsigned(wire183);
            end
          reg208 <= reg197;
        end
      else
        begin
          for (forvar186 = (1'h0); (forvar186 < (3'h4)); forvar186 = (forvar186 + (1'h1)))
            begin
              reg188 <= {$signed($signed((reg191[(2'h3):(1'h1)] ?
                      (~^reg206) : $signed(reg199))))};
              reg189 = $unsigned(reg207[(2'h2):(1'h1)]);
            end
          if ({$unsigned(reg203)})
            begin
              reg190 <= ($signed((!reg200[(4'hb):(4'ha)])) ?
                  $unsigned(((-{wire183}) >>> (~^$signed((8'h9f))))) : $unsigned($unsigned((+$unsigned(reg200)))));
              reg192 = $signed(wire180);
              reg194 = reg194[(3'h6):(1'h1)];
              reg199 <= (8'hb2);
              reg202 <= $unsigned(wire185);
            end
          else
            begin
              reg190 <= $signed($signed(wire183));
              reg191 <= {(8'hb8)};
              reg192 = $signed((reg201 ^ {$signed($unsigned(wire185))}));
              reg194 = wire185[(3'h6):(3'h4)];
              reg195 = $unsigned((&reg208[(1'h1):(1'h0)]));
            end
          reg203 <= (reg187[(1'h0):(1'h0)] || (wire178 ?
              (^~(~|(&reg196))) : wire184));
          if (reg198[(3'h7):(3'h6)])
            begin
              reg207 <= $signed(((~&wire176) < (~^({(8'hbc), wire183} ?
                  $unsigned((8'hac)) : wire185[(4'hb):(2'h3)]))));
              reg208 <= {(({$unsigned((8'hb0)),
                      reg191} != reg187) || wire177[(3'h7):(3'h5)])};
              reg209 = (8'hb2);
            end
          else
            begin
              reg207 <= $unsigned(reg196);
              reg208 <= ((({forvar202[(3'h5):(3'h4)],
                      (&(8'ha5))} >>> (reg204[(4'he):(4'hb)] ?
                      $signed(reg192) : $signed(reg202))) || reg208) ?
                  ((8'h9f) ?
                      reg208 : (&{$unsigned(reg191),
                          ((8'ha6) ?
                              wire182 : wire177)})) : $signed((~&($signed(reg186) != (reg199 ?
                      (8'hb0) : (8'ha7))))));
              reg209 = (&(!$unsigned($unsigned(wire179[(1'h1):(1'h1)]))));
              reg210 <= reg192[(5'h10):(5'h10)];
            end
        end
      if (reg194[(5'h12):(4'hc)])
        begin
          reg211 <= {$unsigned($signed((+(^~reg194))))};
          if ({(reg186 & {reg198, (-(|reg192))})})
            begin
              reg212 = {$unsigned($unsigned($unsigned((reg208 ?
                      (8'ha6) : reg202))))};
            end
          else
            begin
              reg212 = (reg200[(3'h7):(3'h6)] != (|$signed($unsigned($unsigned((8'hb5))))));
              reg213 <= $signed(reg187);
              reg214 = reg201;
              reg215 <= (~(&$signed(((~(8'ha9)) - {reg194}))));
              reg216 <= reg195[(3'h7):(2'h3)];
            end
        end
      else
        begin
          if ($signed($signed((+reg199))))
            begin
              reg211 <= $signed((reg189[(3'h6):(2'h3)] ?
                  (((^reg214) >= {wire182}) ?
                      (-reg192[(3'h4):(2'h3)]) : (|$unsigned((8'ha5)))) : $signed(wire184[(1'h0):(1'h0)])));
              reg213 <= ($signed((~((|reg201) >>> (reg214 ?
                      reg188 : (8'ha3))))) ?
                  wire183[(1'h0):(1'h0)] : (~&$unsigned((reg201[(4'h8):(3'h5)] != (^reg195)))));
              reg214 = ({$signed($signed({wire179})), (~|$signed((^reg190)))} ?
                  $unsigned($signed($unsigned(((8'hb5) ?
                      wire177 : (8'hb3))))) : {($signed(reg213) ~^ reg205),
                      reg190});
              reg215 <= (-$unsigned($unsigned({(~&reg210)})));
              reg217 = reg196[(2'h3):(2'h3)];
            end
          else
            begin
              reg212 = (((&reg200[(2'h2):(1'h0)]) ?
                  (7'h43) : (reg193[(1'h0):(1'h0)] ?
                      (reg201[(2'h2):(1'h0)] ^ (7'h40)) : reg215[(3'h4):(2'h3)])) > ($signed(reg205) >> {$signed((reg210 ?
                      wire177 : reg211))}));
              reg214 = reg211[(2'h3):(1'h0)];
              reg217 = wire182[(4'h9):(3'h6)];
            end
          for (forvar218 = (1'h0); (forvar218 < (2'h3)); forvar218 = (forvar218 + (1'h1)))
            begin
              reg219 = reg203[(1'h0):(1'h0)];
              reg220 <= reg197;
              reg221 <= $signed($signed(((reg204[(4'ha):(1'h0)] ?
                      reg194 : $unsigned(reg212)) ?
                  (+((8'hbf) ? reg196 : wire185)) : {(~|reg219)})));
              reg222 <= {($unsigned(reg212) - {(~|(wire183 ? reg207 : reg210)),
                      $unsigned((+wire180))})};
            end
          reg223 <= (~reg201);
          if (forvar202[(1'h0):(1'h0)])
            begin
              reg224 = wire183;
              reg225 = $unsigned($signed($unsigned((-$signed(reg206)))));
              reg226 <= ($signed(($unsigned((reg212 ?
                      reg203 : reg211)) ^ (^{wire179, reg194}))) ?
                  $unsigned((~&((wire179 & wire181) >= $signed(wire185)))) : wire180);
              reg227 = reg195[(4'ha):(2'h3)];
              reg228 <= (reg224 < $unsigned((!$signed((reg204 | reg198)))));
            end
          else
            begin
              reg224 = reg220;
            end
        end
      reg229 <= reg225[(1'h1):(1'h1)];
      if (reg225)
        begin
          if ((({((wire176 >>> (8'hb7)) ? reg194[(5'h11):(1'h1)] : reg224)} ?
                  wire181 : ((|reg205[(1'h1):(1'h0)]) ?
                      reg222 : $signed($unsigned(wire183)))) ?
              $signed(($signed($signed(reg186)) ~^ $unsigned($unsigned(reg200)))) : reg199[(3'h5):(1'h0)]))
            begin
              reg230 <= ($signed($signed(reg217[(4'hc):(4'hc)])) == reg202);
            end
          else
            begin
              reg230 <= {(&$signed($unsigned($signed(reg199)))),
                  $signed((wire178 ?
                      ($signed(reg194) ?
                          $signed(reg191) : (reg199 - reg213)) : (^$unsigned(reg199))))};
              reg231 <= (^reg204[(5'h11):(4'h8)]);
              reg232 = (($signed($signed((reg217 ?
                  reg187 : reg217))) >= ($unsigned((reg219 ? reg199 : reg222)) ?
                  $signed((wire180 || reg224)) : forvar218)) | {$signed({(reg214 ?
                          reg228 : reg212),
                      (reg214 > reg204)}),
                  ((~|reg202) ? $unsigned((reg187 >>> reg221)) : reg194)});
            end
          if ($unsigned(((({reg200,
              (8'hac)} && reg224) ^~ reg198) <<< (8'hb6))))
            begin
              reg233 <= {$signed($unsigned($signed({reg223}))),
                  (~|$signed((wire179 * (+wire185))))};
            end
          else
            begin
              reg234 = ($unsigned(reg194[(5'h11):(1'h1)]) ?
                  $unsigned(($signed((reg233 ? reg200 : wire182)) ?
                      $signed((~^wire176)) : reg228)) : {wire177});
              reg235 <= $signed((reg221 <<< {((~reg208) ?
                      (&(8'h9e)) : (reg225 ? reg229 : (8'hb0)))}));
            end
          if ($unsigned({reg234, {reg203}}))
            begin
              reg236 <= $unsigned(reg232[(3'h5):(2'h2)]);
              reg237 <= {reg196};
              reg238 = reg208[(2'h2):(2'h2)];
            end
          else
            begin
              reg238 = reg217[(3'h5):(3'h4)];
            end
        end
      else
        begin
          reg230 <= $signed({(({reg222, (8'hb1)} ?
                      forvar202 : (reg200 >> reg232)) ?
                  $unsigned((reg203 ?
                      reg217 : reg213)) : reg217[(4'hc):(4'hc)])});
          for (forvar231 = (1'h0); (forvar231 < (2'h2)); forvar231 = (forvar231 + (1'h1)))
            begin
              reg232 = reg211;
              reg233 <= (({((reg234 ?
                          wire176 : reg189) >>> (~|(8'ha5)))} != ($signed((forvar231 ?
                          (7'h41) : reg229)) ?
                      wire178[(4'hb):(3'h5)] : wire181)) ?
                  $signed(wire182) : reg190);
              reg235 <= (~^(+(((reg238 >>> (8'hbb)) >= $unsigned(reg215)) ^~ $signed((^~(8'hbf))))));
              reg238 = reg233;
              reg239 = reg186[(4'ha):(2'h2)];
            end
          reg240 <= (~$unsigned(reg208));
          if (reg186)
            begin
              reg241 = reg238[(3'h5):(2'h2)];
              reg242 = ((+($unsigned(((8'haa) ? wire180 : reg197)) ?
                  reg208 : $unsigned(reg189[(3'h6):(3'h5)]))) ^ reg194);
              reg243 <= {reg205, reg194[(1'h0):(1'h0)]};
              reg244 <= reg223[(4'h8):(3'h4)];
              reg245 <= (-(!reg196[(1'h1):(1'h1)]));
            end
          else
            begin
              reg241 = (reg211 ?
                  $unsigned($signed($signed($signed(wire181)))) : (8'haa));
              reg243 <= (|($signed(reg220) & (reg195 != {$signed(reg201)})));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar246 = (1'h0); (forvar246 < (1'h1)); forvar246 = (forvar246 + (1'h1)))
        begin
          reg247 <= $unsigned(wire185);
          if ($signed((8'haf)))
            begin
              reg248 = ($unsigned((|((reg229 ? (8'hb0) : wire183) ?
                  reg211[(1'h0):(1'h0)] : ((8'ha9) ?
                      wire183 : reg228)))) >>> reg226);
              reg249 <= (reg247[(3'h4):(3'h4)] >> $signed(($unsigned(reg244[(2'h2):(1'h1)]) ?
                  reg210 : ($signed(reg208) >> {reg244}))));
              reg250 <= ((!reg211[(2'h2):(2'h2)]) ?
                  $signed({(^~(!reg208))}) : (reg193[(5'h11):(4'ha)] & (reg207[(2'h2):(2'h2)] ?
                      ($signed(reg243) & $unsigned(reg203)) : ((reg223 < wire183) > $unsigned((8'hb7))))));
            end
          else
            begin
              reg248 = (^$signed($signed($unsigned((wire177 ^ reg228)))));
            end
          if ((wire177 ?
              reg190 : (^~($unsigned($unsigned(wire179)) != $signed(reg210[(2'h3):(2'h3)])))))
            begin
              reg251 = $unsigned(wire179);
              reg252 = $signed((($signed(reg250[(1'h1):(1'h0)]) ?
                  ((wire178 ?
                      wire180 : (8'hbf)) ^~ reg248[(2'h2):(2'h2)]) : (8'ha6)) >> $unsigned($signed((reg243 ?
                  (7'h43) : wire182)))));
              reg253 <= reg237;
            end
          else
            begin
              reg253 <= reg223;
              reg254 = $unsigned({(8'haf)});
              reg255 = reg210[(1'h1):(1'h1)];
              reg256 <= (reg245 <<< reg254);
            end
          if ((~|{(({(8'hb0)} << (wire177 ?
                  reg222 : (8'haf))) >= $unsigned($unsigned(wire179))),
              $signed(wire182[(3'h7):(3'h5)])}))
            begin
              reg257 = (!reg186[(4'hc):(4'h9)]);
              reg258 <= $unsigned(((reg251 != {$unsigned(reg211), reg231}) ?
                  $unsigned($unsigned($signed(reg215))) : reg233[(4'h9):(3'h6)]));
              reg259 <= {{(~|$signed(reg223[(3'h5):(1'h0)])),
                      (reg245 && reg253[(3'h6):(3'h6)])},
                  (+(($unsigned((7'h44)) ^~ $unsigned(reg211)) != (-((8'hbd) ?
                      reg230 : (8'hb5)))))};
              reg260 <= {(^~$unsigned($signed($unsigned(reg203))))};
              reg261 <= (~|{reg257});
            end
          else
            begin
              reg257 = (reg231 ?
                  $unsigned($signed((!(reg188 ^ wire176)))) : (~|(reg210[(4'hc):(3'h5)] ^ {reg233,
                      reg190})));
              reg258 <= (((($unsigned(reg210) ?
                      (reg221 ?
                          reg213 : (8'hb0)) : reg210) != (!$signed((8'h9c)))) - ($unsigned(reg248[(5'h12):(5'h12)]) >>> (reg257 <<< {reg186}))) ?
                  {reg253[(2'h2):(1'h1)], reg215} : wire178[(1'h1):(1'h1)]);
            end
        end
      if (($unsigned(($signed(reg250) ?
          ({reg245,
              reg202} + reg260) : {(-reg259)})) < $unsigned({((reg207 + reg233) ?
              (reg222 >>> reg215) : reg260),
          (^((7'h40) ? reg249 : (8'ha9)))})))
        begin
          if (reg245[(3'h6):(3'h6)])
            begin
              reg262 <= (reg249 ?
                  wire184[(3'h4):(3'h4)] : (&(reg255[(1'h0):(1'h0)] & $signed($signed(reg245)))));
              reg263 = $unsigned($unsigned(reg236[(3'h5):(3'h4)]));
              reg264 = (7'h43);
            end
          else
            begin
              reg262 <= ((reg213[(3'h4):(2'h3)] + $unsigned(((reg249 > reg244) ?
                  $signed(reg203) : ((8'haf) || reg188)))) | $signed((reg250 ?
                  $signed((-reg257)) : {$unsigned((8'h9f))})));
              reg263 = reg226;
              reg265 <= ($signed(reg250[(2'h2):(1'h0)]) ?
                  ((~|$unsigned((reg259 ? reg260 : reg202))) ?
                      (&(reg245 + {reg203,
                          reg249})) : ($signed($unsigned(reg250)) && ((8'hb6) ?
                          $signed(reg262) : reg208[(3'h4):(3'h4)]))) : $unsigned((^($unsigned(forvar246) >> reg264[(5'h13):(5'h13)]))));
              reg266 = wire178[(2'h3):(1'h1)];
            end
          for (forvar267 = (1'h0); (forvar267 < (1'h0)); forvar267 = (forvar267 + (1'h1)))
            begin
              reg268 <= $signed((~&$signed({(reg211 <<< (7'h40))})));
              reg269 <= {{reg202}, reg233[(3'h6):(1'h0)]};
              reg270 = ((^~reg236[(4'hf):(3'h5)]) << reg255[(1'h1):(1'h1)]);
              reg271 <= reg186[(1'h0):(1'h0)];
            end
          reg272 <= (wire184[(2'h2):(1'h1)] <<< reg237);
          reg273 = (^(~$unsigned({{(8'hbc)}, (~reg271)})));
        end
      else
        begin
          if (wire179)
            begin
              reg263 = reg213[(3'h5):(2'h2)];
              reg265 <= (|reg190[(4'h9):(3'h5)]);
            end
          else
            begin
              reg262 <= (8'h9e);
              reg265 <= $signed(reg243);
              reg267 <= (~(reg258[(1'h0):(1'h0)] ?
                  ((reg251 ?
                      (~^reg264) : (reg220 ?
                          reg235 : wire184)) > ($unsigned(reg268) > (reg240 ?
                      wire183 : reg259))) : $signed(reg220)));
            end
          for (forvar268 = (1'h0); (forvar268 < (2'h2)); forvar268 = (forvar268 + (1'h1)))
            begin
              reg269 <= reg269[(4'hc):(1'h1)];
              reg271 <= $signed(reg220[(5'h11):(4'ha)]);
              reg272 <= $unsigned(wire183[(1'h0):(1'h0)]);
            end
        end
      if ((+(((wire181[(1'h1):(1'h1)] >= (reg255 ?
              reg257 : wire176)) > wire176) ?
          ((~(reg211 ?
              (7'h40) : (8'hb1))) >> reg188[(4'hb):(3'h5)]) : $signed((+{wire176})))))
        begin
          for (forvar274 = (1'h0); (forvar274 < (1'h1)); forvar274 = (forvar274 + (1'h1)))
            begin
              reg275 = reg261[(3'h4):(1'h0)];
              reg276 <= reg199[(5'h12):(2'h3)];
            end
          if (reg253)
            begin
              reg277 <= (-(^~$signed((!(reg215 ? reg260 : reg257)))));
            end
          else
            begin
              reg277 <= (8'hbd);
            end
          reg278 = (+(forvar274 ?
              {(~|reg261),
                  (reg277 ?
                      {reg229,
                          reg237} : $unsigned(reg252))} : reg210[(5'h12):(5'h11)]));
          reg279 = $unsigned((~^(&(8'h9f))));
          for (forvar280 = (1'h0); (forvar280 < (2'h2)); forvar280 = (forvar280 + (1'h1)))
            begin
              reg281 = ({(reg275 != reg237)} >>> (&$unsigned(($signed(reg270) ?
                  $unsigned(wire183) : reg216[(4'hc):(2'h2)]))));
              reg282 = reg245;
              reg283 <= (($signed($signed(reg251[(4'h9):(3'h4)])) + reg235) ?
                  reg276 : ($unsigned($signed((reg221 ?
                      reg257 : reg230))) <= (reg267[(2'h3):(1'h1)] && (~$signed(reg247)))));
              reg284 <= {$signed(reg245[(2'h2):(1'h1)]),
                  ($unsigned($unsigned((reg269 + reg276))) - ($unsigned(reg199[(3'h6):(3'h5)]) & (wire180 ?
                      (reg236 + reg236) : (+reg231))))};
              reg285 <= $signed((reg245 && {{{reg255, reg228},
                      $unsigned(reg226)},
                  $unsigned((wire184 & reg211))}));
            end
        end
      else
        begin
          if ((($unsigned((-reg245[(2'h3):(2'h3)])) ?
                  reg226 : reg248[(4'h8):(2'h2)]) ?
              (-(~|{{(8'hbb),
                      reg285}})) : ((~$signed($signed(reg213))) - ($unsigned({reg190}) ?
                  reg258 : (reg247[(2'h3):(2'h2)] ^~ reg255)))))
            begin
              reg274 <= ($signed((reg244 > ((reg203 ? reg269 : (8'hbb)) ?
                      (&reg245) : {reg202, forvar268}))) ?
                  reg275[(4'h8):(1'h1)] : wire179);
            end
          else
            begin
              reg274 <= (reg251[(2'h3):(1'h0)] ?
                  $signed(reg256) : reg236[(2'h2):(2'h2)]);
              reg276 <= $signed((^~((~&(reg279 ^~ reg235)) ?
                  reg258 : (~|reg208))));
              reg277 <= $unsigned((-$unsigned($unsigned(reg265))));
            end
        end
    end
  assign wire286 = ((|wire180) + reg256[(1'h1):(1'h1)]);
  assign wire287 = $signed($signed(reg259));
  assign wire288 = ($signed($unsigned(wire179[(5'h14):(3'h5)])) ?
                       (~^($signed(reg271) ^~ (~|reg213[(2'h3):(2'h3)]))) : $signed(reg268));
  always
    @(posedge clk) begin
      reg289 = reg231[(2'h3):(1'h0)];
      for (forvar290 = (1'h0); (forvar290 < (1'h0)); forvar290 = (forvar290 + (1'h1)))
        begin
          reg291 = (reg191 ?
              $signed((($unsigned(reg228) ?
                  (reg271 != reg213) : $signed(reg193)) - ((8'hb5) ?
                  $unsigned(wire181) : $signed(wire176)))) : reg236);
          if (reg211)
            begin
              reg292 <= $unsigned(reg253[(2'h3):(2'h2)]);
            end
          else
            begin
              reg292 <= $signed((~$unsigned($unsigned(((8'haa) < reg243)))));
              reg293 <= (reg256 ~^ (~&$unsigned($signed($signed(reg210)))));
              reg294 <= ((&reg276) ? $signed((8'hb1)) : reg272[(3'h7):(3'h5)]);
            end
        end
      for (forvar295 = (1'h0); (forvar295 < (2'h3)); forvar295 = (forvar295 + (1'h1)))
        begin
          if ((~{{(-$unsigned(reg271)),
                  ($signed(reg190) == $unsigned(wire286))}}))
            begin
              reg296 = wire288[(3'h5):(1'h1)];
            end
          else
            begin
              reg297 <= (~^$unsigned(((^wire288[(3'h4):(1'h1)]) << $unsigned((!reg265)))));
              reg298 <= (~&$signed(wire183));
            end
          if ($signed((reg208[(1'h1):(1'h1)] ?
              $unsigned($unsigned($unsigned(wire178))) : (|$unsigned($unsigned(reg228))))))
            begin
              reg299 <= (reg276 ?
                  (&$unsigned(({reg250} - $signed(reg236)))) : $unsigned($unsigned((~&reg222[(2'h2):(1'h0)]))));
              reg300 <= {reg292[(3'h7):(3'h4)]};
            end
          else
            begin
              reg301 = reg269[(1'h0):(1'h0)];
              reg302 <= reg284[(1'h0):(1'h0)];
              reg303 <= reg213;
              reg304 = $signed($signed($signed(((reg222 - reg223) | $signed(reg276)))));
            end
          for (forvar305 = (1'h0); (forvar305 < (1'h0)); forvar305 = (forvar305 + (1'h1)))
            begin
              reg306 <= $unsigned($unsigned((reg188 && ((~|reg256) < reg230[(3'h6):(2'h3)]))));
            end
        end
      reg307 <= wire182;
    end
  assign wire308 = $unsigned(reg292[(4'he):(4'he)]);
  assign wire309 = $unsigned(reg193[(3'h6):(3'h4)]);
  always
    @(posedge clk) begin
      for (forvar310 = (1'h0); (forvar310 < (1'h1)); forvar310 = (forvar310 + (1'h1)))
        begin
          for (forvar311 = (1'h0); (forvar311 < (2'h3)); forvar311 = (forvar311 + (1'h1)))
            begin
              reg312 = ({$unsigned(($signed(reg220) >= $signed(reg215)))} ?
                  forvar311[(1'h1):(1'h0)] : ((~|(8'ha4)) ~^ (reg271 < wire309)));
              reg313 <= $signed($unsigned((wire308[(4'h8):(4'h8)] ?
                  reg231[(3'h4):(2'h2)] : (^~{reg256, reg221}))));
              reg314 <= $unsigned({wire288[(1'h1):(1'h0)],
                  $unsigned(reg243[(4'hd):(2'h2)])});
              reg315 <= {$signed(reg243[(2'h3):(1'h1)])};
            end
          for (forvar316 = (1'h0); (forvar316 < (2'h3)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg317 = reg202;
              reg318 = reg230;
            end
          if (reg315)
            begin
              reg319 <= $unsigned($signed(reg243[(2'h3):(1'h1)]));
              reg320 <= $unsigned(((~&$unsigned({reg267, reg298})) ?
                  $unsigned($unsigned((&reg244))) : $unsigned(((wire286 ?
                          (8'ha3) : (8'h9e)) ?
                      $unsigned(reg230) : (reg223 - reg314)))));
              reg321 = wire185[(1'h0):(1'h0)];
            end
          else
            begin
              reg319 <= reg299;
            end
          if (wire185)
            begin
              reg322 <= ($signed((reg285[(2'h3):(1'h0)] ?
                      reg256 : $signed((reg208 < reg223)))) ?
                  wire286[(4'hd):(4'h8)] : ($signed(reg293) ?
                      reg240[(3'h7):(2'h3)] : {reg321,
                          ($unsigned(reg319) * {reg247})}));
              reg323 <= $signed({$signed($unsigned((reg253 ? reg313 : reg253))),
                  ((reg186[(1'h0):(1'h0)] ? (-wire286) : (8'hbe)) ?
                      (!reg322[(3'h4):(1'h1)]) : reg191)});
              reg324 <= $signed(wire179[(4'hd):(4'h9)]);
            end
          else
            begin
              reg325 = {(~$signed((^(|(8'haf)))))};
              reg326 = $unsigned((reg292 ?
                  $signed(($unsigned(wire288) ?
                      $signed(reg299) : $unsigned(wire180))) : $signed($unsigned($signed(forvar316)))));
              reg327 = $unsigned($unsigned(reg314[(2'h3):(2'h3)]));
            end
          for (forvar328 = (1'h0); (forvar328 < (2'h3)); forvar328 = (forvar328 + (1'h1)))
            begin
              reg329 = ((~|($unsigned(reg233) > $signed(wire178))) ?
                  (~|(~^reg267[(3'h6):(3'h5)])) : $signed($unsigned($unsigned((~(8'hbf))))));
              reg330 <= $unsigned({$signed(reg283)});
              reg331 <= wire308;
              reg332 <= ($unsigned(((~|reg294) * $signed($signed(reg229)))) >>> $signed((~&(~|$unsigned((8'ha4))))));
              reg333 <= reg203[(1'h1):(1'h0)];
            end
        end
      if ((reg313 <= (!$signed(reg319[(4'hb):(2'h3)]))))
        begin
          reg334 = wire308[(3'h7):(3'h5)];
          reg335 <= reg302[(2'h3):(1'h1)];
        end
      else
        begin
          reg335 <= (($signed((^~(8'h9f))) | (((forvar328 ?
                      forvar316 : reg274) <= (wire180 != (8'hbf))) ?
                  {reg235} : (&reg210[(4'hc):(1'h0)]))) ?
              forvar310 : {$signed(((^~reg202) * $unsigned(wire181))),
                  $signed({$unsigned((7'h42)), (8'hae)})});
          reg336 = reg222;
        end
      for (forvar337 = (1'h0); (forvar337 < (2'h3)); forvar337 = (forvar337 + (1'h1)))
        begin
          for (forvar338 = (1'h0); (forvar338 < (3'h4)); forvar338 = (forvar338 + (1'h1)))
            begin
              reg339 <= reg188;
              reg340 <= (wire182 ?
                  {$signed((!(wire176 ? (8'hb4) : reg327)))} : (reg303 ?
                      $unsigned($signed($signed(forvar328))) : (reg221[(2'h3):(1'h1)] << $unsigned(reg258))));
              reg341 <= $unsigned($unsigned((^$signed((^reg203)))));
              reg342 <= reg203;
            end
          reg343 = $unsigned(reg276[(4'h8):(3'h5)]);
          if ((^~(reg283[(4'h9):(4'h8)] | $unsigned(((wire288 ?
                  reg298 : reg324) ?
              (reg268 || reg317) : reg260)))))
            begin
              reg344 <= reg221[(1'h0):(1'h0)];
            end
          else
            begin
              reg344 <= (~^$signed($unsigned({(!forvar338),
                  reg262[(3'h4):(2'h3)]})));
              reg345 = (reg208[(1'h0):(1'h0)] * reg315);
            end
        end
    end
  assign wire346 = reg340;
  assign wire347 = (reg276[(4'ha):(2'h2)] ?
                       $signed($signed(wire287[(4'hb):(3'h4)])) : (&$unsigned(reg216[(1'h0):(1'h0)])));
  assign wire348 = reg274;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module571  (y, clk, wire575, wire574, wire573, wire572);
  output wire [(32'h188):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire575;
  input wire signed [(4'hb):(1'h0)] wire574;
  input wire [(5'h12):(1'h0)] wire573;
  input wire [(5'h11):(1'h0)] wire572;
  wire signed [(5'h13):(1'h0)] wire606;
  wire signed [(4'hf):(1'h0)] wire605;
  wire signed [(5'h10):(1'h0)] wire604;
  wire signed [(5'h13):(1'h0)] wire603;
  wire signed [(3'h5):(1'h0)] wire602;
  wire signed [(5'h11):(1'h0)] wire601;
  wire signed [(4'h9):(1'h0)] wire600;
  wire [(4'hc):(1'h0)] wire599;
  wire signed [(5'h15):(1'h0)] wire598;
  wire signed [(4'h9):(1'h0)] wire597;
  wire signed [(4'he):(1'h0)] wire596;
  wire [(4'hd):(1'h0)] wire580;
  wire [(3'h5):(1'h0)] wire579;
  wire [(4'hb):(1'h0)] wire578;
  wire [(5'h12):(1'h0)] wire577;
  wire [(4'hb):(1'h0)] wire576;
  reg [(4'hb):(1'h0)] reg595 = (1'h0);
  reg [(5'h14):(1'h0)] reg592 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg591 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg590 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg588 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg586 = (1'h0);
  reg [(4'hb):(1'h0)] reg585 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg584 = (1'h0);
  reg [(4'hf):(1'h0)] reg582 = (1'h0);
  reg [(2'h3):(1'h0)] reg594 = (1'h0);
  reg [(4'ha):(1'h0)] forvar593 = (1'h0);
  reg [(3'h7):(1'h0)] reg589 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg587 = (1'h0);
  reg [(4'hd):(1'h0)] forvar583 = (1'h0);
  reg [(4'he):(1'h0)] reg581 = (1'h0);
  assign y = {wire606,
                 wire605,
                 wire604,
                 wire603,
                 wire602,
                 wire601,
                 wire600,
                 wire599,
                 wire598,
                 wire597,
                 wire596,
                 wire580,
                 wire579,
                 wire578,
                 wire577,
                 wire576,
                 reg595,
                 reg592,
                 reg591,
                 reg590,
                 reg588,
                 reg586,
                 reg585,
                 reg584,
                 reg582,
                 reg594,
                 forvar593,
                 reg589,
                 reg587,
                 forvar583,
                 reg581,
                 (1'h0)};
  assign wire576 = wire572[(4'h9):(3'h4)];
  assign wire577 = (|wire573[(4'h8):(3'h6)]);
  assign wire578 = (wire574 ? wire576 : (^~(-$unsigned($unsigned(wire572)))));
  assign wire579 = (-$unsigned((&$signed((wire572 ? wire573 : wire573)))));
  assign wire580 = (^{($signed((+(8'haa))) ?
                           ($signed((7'h40)) ?
                               (wire578 <<< (8'hb9)) : wire576[(2'h2):(1'h0)]) : {(~&wire573)}),
                       (($signed((8'hbc)) ?
                           $unsigned(wire577) : ((8'hbe) <= wire577)) && {(wire578 || wire575)})});
  always
    @(posedge clk) begin
      reg581 = $signed(wire573[(3'h4):(2'h2)]);
      reg582 <= wire572[(5'h10):(4'hb)];
      for (forvar583 = (1'h0); (forvar583 < (1'h1)); forvar583 = (forvar583 + (1'h1)))
        begin
          reg584 <= (-(&$signed(reg581[(4'hc):(1'h1)])));
          reg585 <= {(~|{$unsigned($unsigned(wire573))})};
          if ((~(&$unsigned($unsigned(wire573[(4'h9):(3'h4)])))))
            begin
              reg586 <= (^wire575[(4'ha):(3'h7)]);
              reg587 = (reg581[(3'h7):(3'h4)] ?
                  (|($unsigned((reg581 ?
                      reg586 : reg585)) ~^ reg586)) : wire572[(4'ha):(3'h4)]);
              reg588 <= (wire579 ?
                  ((($signed((8'hbf)) ?
                      (~^(8'ha7)) : (wire576 < reg587)) + (+$unsigned(reg581))) <<< ((wire579[(1'h1):(1'h1)] && $unsigned(reg585)) ?
                      $signed(wire574) : (~$signed(wire573)))) : (wire576[(4'hb):(2'h2)] ?
                      (8'hac) : wire577));
              reg589 = ($unsigned(((&(~^wire580)) > (((8'ha7) >>> wire579) * (+(8'hb3))))) ?
                  reg582[(4'hc):(1'h1)] : $signed($unsigned(wire575)));
            end
          else
            begin
              reg587 = (8'hbc);
              reg588 <= $signed(reg589);
              reg590 <= ($unsigned((-((wire578 < wire578) ?
                      (wire572 ~^ wire577) : $unsigned((8'hb1))))) ?
                  reg584[(4'h8):(3'h7)] : $unsigned((wire573[(3'h4):(1'h0)] >>> (wire574[(2'h2):(1'h1)] ?
                      (~&forvar583) : {reg582}))));
              reg591 <= {wire576[(1'h0):(1'h0)]};
              reg592 <= (($unsigned(reg589) ^~ $signed($signed({(8'ha4),
                      wire576}))) ?
                  ($signed((~^forvar583[(3'h6):(1'h1)])) & $unsigned((^~(reg591 ?
                      reg591 : reg591)))) : reg582[(3'h4):(3'h4)]);
            end
        end
      for (forvar593 = (1'h0); (forvar593 < (1'h0)); forvar593 = (forvar593 + (1'h1)))
        begin
          if (wire573)
            begin
              reg594 = ((wire577[(4'he):(4'hb)] ?
                      (reg592 < {{reg585,
                              reg585}}) : ((~|reg584[(2'h3):(2'h3)]) ?
                          $unsigned({reg591}) : (wire579[(3'h4):(1'h0)] ?
                              $signed(reg586) : (wire579 ?
                                  wire575 : wire576)))) ?
                  (^(&((wire580 ? reg585 : reg590) == reg588))) : forvar593);
            end
          else
            begin
              reg595 <= (($unsigned((wire580 ^~ reg590)) >>> $unsigned((&((8'ha3) ?
                  reg581 : wire573)))) ~^ reg592[(2'h2):(2'h2)]);
            end
        end
    end
  assign wire596 = {((wire579[(1'h1):(1'h1)] ^ ((|(8'hb7)) ?
                               $unsigned(wire573) : (wire580 ?
                                   reg586 : reg582))) ?
                           {wire575[(1'h1):(1'h1)], reg592} : (wire580 ?
                               (!$unsigned(reg595)) : {(wire579 ?
                                       reg585 : reg585)}))};
  assign wire597 = reg585[(2'h2):(2'h2)];
  assign wire598 = $signed(((($unsigned(wire576) + reg585[(1'h1):(1'h0)]) >>> wire578) + $signed($unsigned($unsigned(wire573)))));
  assign wire599 = (|(~|(!{(~^(8'h9e)), (reg582 < wire598)})));
  assign wire600 = wire575[(4'he):(3'h5)];
  assign wire601 = (-$unsigned(wire598));
  assign wire602 = wire574[(3'h4):(1'h1)];
  assign wire603 = wire573[(3'h5):(1'h0)];
  assign wire604 = (~|reg588);
  assign wire605 = reg590[(3'h5):(2'h2)];
  assign wire606 = wire605;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module464  (y, clk, wire468, wire467, wire466, wire465);
  output wire [(32'h1f8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire468;
  input wire [(3'h6):(1'h0)] wire467;
  input wire [(3'h6):(1'h0)] wire466;
  input wire [(2'h2):(1'h0)] wire465;
  wire [(4'ha):(1'h0)] wire510;
  wire [(5'h12):(1'h0)] wire472;
  wire signed [(3'h7):(1'h0)] wire471;
  wire [(5'h10):(1'h0)] wire470;
  wire signed [(5'h14):(1'h0)] wire469;
  reg [(2'h3):(1'h0)] reg508 = (1'h0);
  reg [(3'h7):(1'h0)] reg507 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg503 = (1'h0);
  reg [(5'h10):(1'h0)] reg501 = (1'h0);
  reg [(4'he):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg497 = (1'h0);
  reg signed [(4'he):(1'h0)] reg496 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg490 = (1'h0);
  reg [(4'he):(1'h0)] reg486 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg485 = (1'h0);
  reg [(4'hb):(1'h0)] reg484 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg482 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg478 = (1'h0);
  reg [(4'ha):(1'h0)] reg477 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg474 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg473 = (1'h0);
  reg [(4'hf):(1'h0)] reg509 = (1'h0);
  reg [(3'h5):(1'h0)] reg506 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg502 = (1'h0);
  reg [(4'he):(1'h0)] forvar500 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg498 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg495 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg494 = (1'h0);
  reg [(5'h10):(1'h0)] forvar493 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg491 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg489 = (1'h0);
  reg [(4'hb):(1'h0)] forvar488 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg487 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg483 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg481 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg479 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar476 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg475 = (1'h0);
  assign y = {wire510,
                 wire472,
                 wire471,
                 wire470,
                 wire469,
                 reg508,
                 reg507,
                 reg505,
                 reg504,
                 reg503,
                 reg501,
                 reg499,
                 reg497,
                 reg496,
                 reg492,
                 reg490,
                 reg486,
                 reg485,
                 reg484,
                 reg482,
                 reg480,
                 reg478,
                 reg477,
                 reg474,
                 reg473,
                 reg509,
                 reg506,
                 reg502,
                 forvar500,
                 reg498,
                 reg495,
                 reg494,
                 forvar493,
                 reg491,
                 reg489,
                 forvar488,
                 reg487,
                 reg483,
                 reg481,
                 reg479,
                 forvar476,
                 reg475,
                 (1'h0)};
  assign wire469 = (((!$signed($unsigned(wire467))) ?
                           wire465[(1'h0):(1'h0)] : wire465) ?
                       (-wire465) : ({$signed((&wire468)),
                               $unsigned({wire466, wire466})} ?
                           $signed((+wire465)) : $unsigned(wire467[(3'h4):(2'h3)])));
  assign wire470 = $signed((~{wire468}));
  assign wire471 = (wire465[(1'h1):(1'h0)] >> {$unsigned($signed((wire467 ?
                           wire466 : wire466)))});
  assign wire472 = wire468;
  always
    @(posedge clk) begin
      if (wire466)
        begin
          if (wire470[(3'h4):(2'h2)])
            begin
              reg473 <= wire467;
            end
          else
            begin
              reg473 <= wire472;
              reg474 <= ($signed(((~&(wire471 ~^ wire465)) ?
                  wire470[(4'hf):(4'hc)] : ((wire471 ? wire465 : wire469) ?
                      wire469 : (&wire467)))) || wire465);
              reg475 = $signed({(wire472 ?
                      (~^$unsigned(wire469)) : ({(8'ha9)} >= $signed(wire468))),
                  $unsigned($unsigned((&(8'ha5))))});
            end
          for (forvar476 = (1'h0); (forvar476 < (1'h1)); forvar476 = (forvar476 + (1'h1)))
            begin
              reg477 <= (+$unsigned((wire467 ?
                  $unsigned($signed(wire469)) : (-$signed((8'hbb))))));
              reg478 <= wire471;
              reg479 = (wire469[(3'h6):(3'h4)] ?
                  reg477[(4'h8):(4'h8)] : $signed(wire468[(2'h3):(1'h0)]));
              reg480 <= ($unsigned(($signed($unsigned(reg479)) ?
                      wire465 : ((-reg479) ?
                          ((8'h9e) || wire467) : $signed(wire471)))) ?
                  reg474 : wire472[(4'hf):(3'h6)]);
              reg481 = $unsigned(wire466);
            end
          reg482 <= wire465[(1'h0):(1'h0)];
        end
      else
        begin
          reg475 = (7'h43);
          for (forvar476 = (1'h0); (forvar476 < (1'h1)); forvar476 = (forvar476 + (1'h1)))
            begin
              reg479 = $signed((-$signed((&$unsigned(wire472)))));
              reg480 <= ((8'ha7) ?
                  (($unsigned($unsigned(reg477)) * ($signed(wire467) | (8'ha5))) - (reg475 ?
                      reg482[(3'h7):(2'h2)] : reg473[(5'h10):(1'h0)])) : $signed(((~$unsigned(wire467)) ?
                      $signed((^reg474)) : reg475[(4'hd):(2'h2)])));
              reg482 <= (^$signed($signed(reg482)));
              reg483 = ({($signed((reg478 != reg481)) ?
                      ((wire470 ? wire469 : wire469) ?
                          (8'ha0) : wire472[(3'h4):(2'h3)]) : reg474[(2'h2):(1'h1)]),
                  $signed(wire468)} ^ (~^forvar476));
              reg484 <= $signed((^(~^forvar476[(3'h4):(2'h2)])));
            end
        end
      reg485 <= $signed((7'h44));
      reg486 <= reg473[(2'h2):(1'h1)];
      if ((8'ha7))
        begin
          reg487 = wire468[(1'h0):(1'h0)];
        end
      else
        begin
          reg487 = wire466[(1'h0):(1'h0)];
          for (forvar488 = (1'h0); (forvar488 < (2'h2)); forvar488 = (forvar488 + (1'h1)))
            begin
              reg489 = ((wire467[(2'h3):(2'h2)] ?
                  wire467 : (!(reg481 ?
                      ((8'h9f) ?
                          wire469 : wire471) : (~wire469)))) << $unsigned((reg481 << $unsigned((forvar488 ^ reg485)))));
              reg490 <= reg474[(3'h5):(3'h4)];
              reg491 = $signed(wire468);
              reg492 <= (^~reg490[(4'he):(4'h9)]);
            end
          for (forvar493 = (1'h0); (forvar493 < (2'h2)); forvar493 = (forvar493 + (1'h1)))
            begin
              reg494 = (~^$unsigned((~|forvar493)));
              reg495 = reg492;
              reg496 <= (forvar488[(1'h0):(1'h0)] ?
                  (~^(!$signed($unsigned(wire467)))) : (^~(wire471[(2'h2):(1'h0)] ?
                      (reg486[(3'h7):(3'h6)] && forvar493) : {{wire469,
                              (8'haf)}})));
            end
          reg497 <= ((8'hb3) || ($signed(wire468[(3'h5):(1'h1)]) >= (reg494[(2'h2):(1'h1)] ?
              {(&wire467)} : ($signed(reg481) >> (forvar493 ?
                  reg483 : wire466)))));
          if (wire471[(3'h4):(2'h3)])
            begin
              reg498 = (^(!$signed(reg485)));
            end
          else
            begin
              reg499 <= (({$unsigned(reg482)} ?
                      reg478[(3'h7):(1'h1)] : ((~&$signed(reg484)) << $signed(((8'ha7) >= wire472)))) ?
                  reg485 : (~^(&($unsigned((8'ha0)) ~^ reg484))));
            end
        end
      for (forvar500 = (1'h0); (forvar500 < (2'h3)); forvar500 = (forvar500 + (1'h1)))
        begin
          if ((&((8'hbe) * (reg475 ?
              {$signed(forvar488),
                  $unsigned(reg474)} : reg497[(4'h9):(3'h6)]))))
            begin
              reg501 <= $signed($signed($unsigned($unsigned((!(8'ha2))))));
            end
          else
            begin
              reg502 = reg498[(2'h2):(2'h2)];
              reg503 <= $signed((wire471[(1'h0):(1'h0)] ?
                  (-(wire472[(5'h11):(4'hd)] ?
                      ((8'haf) ?
                          forvar500 : wire468) : (wire471 & reg481))) : {reg474[(2'h3):(1'h0)],
                      $unsigned((reg496 + reg478))}));
            end
          if ({$unsigned((+$unsigned((reg486 && reg497))))})
            begin
              reg504 <= (&forvar488[(4'h9):(3'h7)]);
              reg505 <= ((~|{$signed($unsigned(reg497))}) < (^(!reg501)));
            end
          else
            begin
              reg504 <= $signed(reg485);
              reg506 = reg494[(1'h1):(1'h1)];
              reg507 <= $unsigned($unsigned($unsigned($signed({reg497,
                  wire469}))));
              reg508 <= ((8'ha6) < (8'hbd));
              reg509 = (^wire472);
            end
        end
    end
  assign wire510 = (|(+(&((^reg474) ? (8'hbd) : (^reg478)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module364  (y, clk, wire368, wire367, wire366, wire365);
  output wire [(32'h417):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire368;
  input wire [(2'h2):(1'h0)] wire367;
  input wire [(3'h6):(1'h0)] wire366;
  input wire signed [(4'h8):(1'h0)] wire365;
  wire signed [(5'h13):(1'h0)] wire460;
  wire signed [(2'h3):(1'h0)] wire459;
  wire signed [(5'h13):(1'h0)] wire425;
  wire signed [(4'h9):(1'h0)] wire424;
  wire signed [(5'h14):(1'h0)] wire395;
  wire [(3'h5):(1'h0)] wire394;
  wire [(5'h13):(1'h0)] wire393;
  wire signed [(4'hd):(1'h0)] wire392;
  wire [(3'h6):(1'h0)] wire391;
  wire [(3'h7):(1'h0)] wire372;
  wire signed [(2'h2):(1'h0)] wire371;
  wire signed [(4'h9):(1'h0)] wire370;
  wire signed [(5'h13):(1'h0)] wire369;
  reg signed [(4'ha):(1'h0)] reg457 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg456 = (1'h0);
  reg [(4'hd):(1'h0)] reg455 = (1'h0);
  reg signed [(4'he):(1'h0)] reg453 = (1'h0);
  reg [(3'h5):(1'h0)] reg450 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg448 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg447 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg441 = (1'h0);
  reg [(4'he):(1'h0)] reg439 = (1'h0);
  reg [(5'h13):(1'h0)] reg435 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg433 = (1'h0);
  reg [(2'h2):(1'h0)] reg432 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg429 = (1'h0);
  reg [(5'h15):(1'h0)] reg423 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg422 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg421 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg418 = (1'h0);
  reg [(4'h8):(1'h0)] reg417 = (1'h0);
  reg [(2'h2):(1'h0)] reg415 = (1'h0);
  reg [(5'h12):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg405 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg404 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg403 = (1'h0);
  reg [(5'h15):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg398 = (1'h0);
  reg [(4'he):(1'h0)] reg390 = (1'h0);
  reg [(2'h3):(1'h0)] reg388 = (1'h0);
  reg [(4'h8):(1'h0)] reg387 = (1'h0);
  reg [(4'h9):(1'h0)] reg386 = (1'h0);
  reg [(3'h6):(1'h0)] reg384 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg381 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg380 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg377 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg376 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg374 = (1'h0);
  reg [(5'h10):(1'h0)] reg373 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg458 = (1'h0);
  reg [(4'he):(1'h0)] reg454 = (1'h0);
  reg [(4'h9):(1'h0)] reg452 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg451 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg449 = (1'h0);
  reg [(4'hf):(1'h0)] forvar446 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar445 = (1'h0);
  reg [(3'h6):(1'h0)] reg444 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar443 = (1'h0);
  reg [(5'h10):(1'h0)] reg442 = (1'h0);
  reg [(4'hf):(1'h0)] reg440 = (1'h0);
  reg signed [(4'he):(1'h0)] reg438 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg437 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg436 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar434 = (1'h0);
  reg [(3'h4):(1'h0)] reg431 = (1'h0);
  reg [(3'h4):(1'h0)] reg430 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg428 = (1'h0);
  reg [(4'h9):(1'h0)] reg427 = (1'h0);
  reg [(2'h2):(1'h0)] forvar426 = (1'h0);
  reg signed [(4'he):(1'h0)] reg420 = (1'h0);
  reg [(5'h15):(1'h0)] reg419 = (1'h0);
  reg [(3'h5):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar414 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg413 = (1'h0);
  reg signed [(4'he):(1'h0)] reg412 = (1'h0);
  reg [(5'h13):(1'h0)] forvar411 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg410 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg408 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg407 = (1'h0);
  reg [(5'h12):(1'h0)] reg406 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg402 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar400 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg399 = (1'h0);
  reg [(3'h4):(1'h0)] forvar397 = (1'h0);
  reg [(3'h7):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg389 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg385 = (1'h0);
  reg [(3'h6):(1'h0)] reg383 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg382 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar378 = (1'h0);
  reg [(3'h7):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar373 = (1'h0);
  assign y = {wire460,
                 wire459,
                 wire425,
                 wire424,
                 wire395,
                 wire394,
                 wire393,
                 wire392,
                 wire391,
                 wire372,
                 wire371,
                 wire370,
                 wire369,
                 reg457,
                 reg456,
                 reg455,
                 reg453,
                 reg450,
                 reg448,
                 reg447,
                 reg441,
                 reg439,
                 reg435,
                 reg433,
                 reg432,
                 reg429,
                 reg423,
                 reg422,
                 reg421,
                 reg418,
                 reg417,
                 reg415,
                 reg409,
                 reg405,
                 reg404,
                 reg403,
                 reg401,
                 reg398,
                 reg390,
                 reg388,
                 reg387,
                 reg386,
                 reg384,
                 reg381,
                 reg380,
                 reg379,
                 reg377,
                 reg376,
                 reg374,
                 reg373,
                 reg458,
                 reg454,
                 reg452,
                 reg451,
                 reg449,
                 forvar446,
                 forvar445,
                 reg444,
                 forvar443,
                 reg442,
                 reg440,
                 reg438,
                 reg437,
                 reg436,
                 forvar434,
                 reg431,
                 reg430,
                 reg428,
                 reg427,
                 forvar426,
                 reg420,
                 reg419,
                 reg416,
                 forvar414,
                 reg413,
                 reg412,
                 forvar411,
                 reg410,
                 reg408,
                 reg407,
                 reg406,
                 reg402,
                 forvar400,
                 reg399,
                 forvar397,
                 reg396,
                 reg389,
                 reg385,
                 reg383,
                 reg382,
                 forvar378,
                 reg375,
                 forvar373,
                 (1'h0)};
  assign wire369 = $unsigned(({(8'h9e)} >> $signed((&wire368))));
  assign wire370 = ({wire369[(5'h12):(4'ha)]} >>> wire368);
  assign wire371 = wire366[(3'h5):(3'h4)];
  assign wire372 = $unsigned(wire368);
  always
    @(posedge clk) begin
      if ($signed($signed(wire372)))
        begin
          if ((^~(wire367 ?
              (^(!$signed(wire368))) : $unsigned((wire368[(3'h5):(1'h0)] ?
                  (wire371 ^~ wire371) : wire366[(3'h6):(3'h5)])))))
            begin
              reg373 <= (&$unsigned({wire369, $unsigned($unsigned(wire369))}));
              reg374 <= (^$signed((~(((8'hbb) ? wire365 : (8'hbb)) * (wire365 ?
                  wire371 : wire370)))));
            end
          else
            begin
              reg373 <= (wire372 ?
                  (|wire371[(2'h2):(1'h1)]) : $unsigned($unsigned($unsigned((-wire370)))));
            end
        end
      else
        begin
          for (forvar373 = (1'h0); (forvar373 < (2'h3)); forvar373 = (forvar373 + (1'h1)))
            begin
              reg375 = wire365;
              reg376 <= forvar373;
              reg377 <= (&wire368[(4'h8):(1'h0)]);
            end
        end
      for (forvar378 = (1'h0); (forvar378 < (1'h0)); forvar378 = (forvar378 + (1'h1)))
        begin
          if ((^(~^(8'hb0))))
            begin
              reg379 <= reg375;
              reg380 <= wire367;
              reg381 <= $unsigned({$unsigned(wire369),
                  $unsigned($signed(wire366))});
            end
          else
            begin
              reg379 <= $unsigned(($unsigned(reg380) ?
                  $signed($unsigned(reg377[(3'h4):(3'h4)])) : (({reg381} ?
                          {forvar378, wire372} : wire368[(3'h4):(1'h1)]) ?
                      (forvar378[(5'h10):(5'h10)] ?
                          (|(8'ha7)) : $unsigned((8'hab))) : (+(8'hbb)))));
              reg382 = forvar373[(2'h2):(2'h2)];
              reg383 = $signed({(~&$unsigned((wire370 >= forvar373))), reg379});
              reg384 <= forvar373;
            end
          if ((~&$signed((&((reg381 ? reg380 : reg375) ?
              (+reg377) : $signed(wire370))))))
            begin
              reg385 = $unsigned($unsigned($signed(((!wire368) ?
                  (reg377 + reg380) : forvar373))));
            end
          else
            begin
              reg386 <= $signed($signed($unsigned({((8'haa) ?
                      reg381 : (8'h9d))})));
              reg387 <= (^((forvar373[(2'h2):(1'h1)] ?
                  (^~(reg377 ? wire365 : wire368)) : (-reg376)) ~^ reg384));
              reg388 <= {$signed((~^$unsigned((reg382 <= reg382))))};
              reg389 = $signed(({(^((8'ha1) ? reg382 : reg380))} ?
                  (+reg380) : (reg384 >> {wire371, $signed(reg387)})));
            end
          reg390 <= $unsigned($unsigned($signed(reg387)));
        end
    end
  assign wire391 = ($unsigned($signed($unsigned(reg390))) ?
                       wire372 : (((+wire365[(4'h8):(1'h0)]) ?
                               ((reg387 >= reg390) < $signed(wire368)) : reg377) ?
                           (reg384 == ({(8'hb0), reg379} ?
                               reg373 : reg379[(4'h9):(3'h5)])) : {$signed($signed(reg390)),
                               $unsigned(wire371[(1'h0):(1'h0)])}));
  assign wire392 = {(8'ha6)};
  assign wire393 = ($unsigned($signed(wire392[(3'h5):(1'h1)])) | reg381[(2'h3):(1'h0)]);
  assign wire394 = (~^($signed({(reg381 ? wire370 : reg374),
                           (wire371 ? reg387 : (8'hb6))}) ?
                       {($signed(reg387) ?
                               reg377 : $unsigned(reg386))} : wire367[(1'h1):(1'h0)]));
  assign wire395 = wire367[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg396 = wire394;
      for (forvar397 = (1'h0); (forvar397 < (1'h0)); forvar397 = (forvar397 + (1'h1)))
        begin
          if (({(^(reg374[(3'h5):(2'h3)] && ((8'hae) ? (8'hb9) : wire394))),
                  (($unsigned((8'ha9)) <<< $signed(reg390)) ~^ wire392[(3'h5):(1'h0)])} ?
              (($signed($signed(wire392)) ?
                      (~|reg376) : ((reg396 && wire371) ^~ wire392[(2'h2):(2'h2)])) ?
                  $signed((((8'hbc) <<< reg384) ~^ (wire365 != reg390))) : (!$signed((8'haf)))) : $signed(reg373[(3'h4):(3'h4)])))
            begin
              reg398 <= forvar397[(2'h3):(1'h0)];
              reg399 = $unsigned(((^((~|wire368) ?
                      reg386 : (wire394 < reg387))) ?
                  ((~^wire370[(2'h2):(1'h0)]) ?
                      $signed($unsigned((8'hb3))) : wire395) : {{(&reg388)},
                      (reg398[(2'h2):(1'h0)] ?
                          wire392 : reg387[(3'h6):(2'h2)])}));
            end
          else
            begin
              reg398 <= wire371[(1'h0):(1'h0)];
            end
          for (forvar400 = (1'h0); (forvar400 < (2'h3)); forvar400 = (forvar400 + (1'h1)))
            begin
              reg401 <= $unsigned((((((8'had) >> wire394) < $unsigned(reg374)) ?
                  $unsigned((|reg374)) : $signed($signed(reg386))) ^~ $unsigned($signed((wire368 < wire371)))));
              reg402 = $signed($signed(wire369));
              reg403 <= $signed((^~(forvar397 & (reg386[(2'h2):(1'h1)] && reg388[(1'h1):(1'h0)]))));
              reg404 <= reg381;
            end
          if ($unsigned((wire370 ?
              $signed({wire365}) : (($unsigned(reg377) && ((8'hbf) ?
                      reg377 : wire368)) ?
                  (reg387[(2'h3):(2'h3)] ?
                      $unsigned(wire370) : $unsigned(wire369)) : $unsigned($unsigned(reg398))))))
            begin
              reg405 <= ($unsigned(reg396) >= (^reg404[(1'h0):(1'h0)]));
              reg406 = reg380[(1'h0):(1'h0)];
              reg407 = wire370;
              reg408 = {(((~$signed(wire366)) ?
                          {(reg402 > wire394),
                              reg406} : ({wire367} || (-(8'hb3)))) ?
                      $unsigned(($unsigned(reg379) & $signed(reg384))) : (wire371[(1'h0):(1'h0)] <= $unsigned(reg377)))};
            end
          else
            begin
              reg406 = reg376[(1'h0):(1'h0)];
              reg407 = reg373;
            end
          if ((8'hb7))
            begin
              reg409 <= (wire368[(3'h5):(3'h4)] >= ($signed($unsigned($signed((8'hb8)))) ?
                  $unsigned(wire370[(3'h7):(2'h2)]) : (^~wire365[(2'h3):(2'h3)])));
              reg410 = ($signed((~&reg398[(4'he):(4'hb)])) ?
                  reg374 : $unsigned($signed(($signed((7'h43)) ?
                      {wire367, reg408} : forvar397[(2'h2):(1'h1)]))));
            end
          else
            begin
              reg410 = (reg374 > (forvar400 ~^ $unsigned($unsigned($signed(reg402)))));
            end
        end
      for (forvar411 = (1'h0); (forvar411 < (2'h3)); forvar411 = (forvar411 + (1'h1)))
        begin
          reg412 = $signed(reg402);
          reg413 = wire369[(4'ha):(4'ha)];
          for (forvar414 = (1'h0); (forvar414 < (3'h4)); forvar414 = (forvar414 + (1'h1)))
            begin
              reg415 <= reg401;
              reg416 = $signed($unsigned(wire394[(3'h4):(3'h4)]));
            end
          reg417 <= $signed(reg413);
          if ((^((~|((!wire367) * {reg374})) - $signed(($unsigned(reg373) ?
              {reg386, (8'hb3)} : (wire366 ^~ forvar400))))))
            begin
              reg418 <= ($signed(($signed(wire372) | $signed((reg387 ^ forvar414)))) ?
                  (wire394 ?
                      $signed(($signed(wire395) != (reg401 + forvar411))) : (^((&(8'hb2)) ?
                          $unsigned(reg399) : wire393[(3'h4):(2'h3)]))) : reg417);
              reg419 = (&$signed($unsigned({((8'hbc) && reg416)})));
              reg420 = $signed((~&$signed((8'ha1))));
              reg421 <= $unsigned((+reg413[(2'h3):(1'h1)]));
              reg422 <= forvar414[(4'hf):(2'h2)];
            end
          else
            begin
              reg419 = ((($unsigned((reg377 <<< reg417)) ?
                      {(forvar400 * reg379)} : (~^(reg384 <= wire372))) << $unsigned(($unsigned(forvar414) ?
                      (~reg415) : (8'hb7)))) ?
                  (reg420 ^~ (~^$signed({(8'hb6)}))) : ($unsigned((8'haf)) ?
                      $unsigned(((wire391 ?
                          reg401 : reg407) && reg390)) : reg381[(1'h1):(1'h1)]));
              reg421 <= reg421;
              reg422 <= reg413;
              reg423 <= ((^(~($signed(forvar414) == reg398))) <<< ($signed((^(reg421 ?
                  reg399 : wire368))) ^ {$unsigned(wire394[(3'h4):(3'h4)])}));
            end
        end
    end
  assign wire424 = {$unsigned($unsigned((reg374 << (~reg417)))),
                       (reg388[(2'h2):(2'h2)] | $unsigned(wire371[(2'h2):(2'h2)]))};
  assign wire425 = reg417;
  always
    @(posedge clk) begin
      for (forvar426 = (1'h0); (forvar426 < (1'h1)); forvar426 = (forvar426 + (1'h1)))
        begin
          reg427 = (-(reg390 ? wire392 : reg401));
          if (reg417)
            begin
              reg428 = $signed(reg384[(2'h3):(1'h1)]);
            end
          else
            begin
              reg429 <= (^$signed((~|reg376[(3'h4):(2'h2)])));
              reg430 = wire366;
              reg431 = (8'h9f);
              reg432 <= wire367[(1'h1):(1'h0)];
              reg433 <= wire370;
            end
        end
      for (forvar434 = (1'h0); (forvar434 < (2'h2)); forvar434 = (forvar434 + (1'h1)))
        begin
          if (wire369)
            begin
              reg435 <= (((reg418[(2'h2):(1'h0)] ?
                          wire372 : reg427[(3'h7):(3'h6)]) ?
                      wire424 : reg409) ?
                  $unsigned((|$unsigned($unsigned(reg428)))) : reg430[(3'h4):(2'h2)]);
              reg436 = $unsigned($signed(reg432));
              reg437 = reg379;
              reg438 = $unsigned(wire367);
            end
          else
            begin
              reg436 = reg421[(3'h4):(2'h3)];
              reg439 <= {wire393,
                  $signed(((~$unsigned(reg435)) ?
                      ($unsigned(reg433) ?
                          (8'ha4) : (-reg415)) : (|(reg427 != reg380))))};
              reg440 = ({(({reg432, reg418} ?
                              $signed(reg423) : $unsigned(reg415)) ?
                          reg376 : {$signed(wire366)}),
                      reg381} ?
                  (&(^$unsigned((reg403 <<< reg417)))) : $unsigned(forvar434[(3'h7):(3'h4)]));
              reg441 <= $unsigned($unsigned($signed($unsigned((+reg428)))));
              reg442 = $unsigned($unsigned({(!reg437)}));
            end
        end
      for (forvar443 = (1'h0); (forvar443 < (2'h2)); forvar443 = (forvar443 + (1'h1)))
        begin
          reg444 = $signed(reg404[(2'h2):(1'h0)]);
        end
      for (forvar445 = (1'h0); (forvar445 < (3'h4)); forvar445 = (forvar445 + (1'h1)))
        begin
          for (forvar446 = (1'h0); (forvar446 < (2'h3)); forvar446 = (forvar446 + (1'h1)))
            begin
              reg447 <= $signed((|(reg438[(4'h8):(3'h5)] ?
                  $unsigned($unsigned(reg435)) : $signed((wire424 & wire370)))));
            end
          if ((^(({(reg405 ? reg441 : reg433)} ?
              (&$signed(reg415)) : wire425[(4'h8):(1'h1)]) * reg388[(1'h0):(1'h0)])))
            begin
              reg448 <= (($unsigned(reg405[(4'h9):(3'h6)]) >= reg428) >>> ({wire391[(3'h6):(2'h2)]} ^~ forvar426));
              reg449 = (+$unsigned($unsigned({reg405[(3'h7):(3'h7)]})));
              reg450 <= $signed($unsigned(reg380));
            end
          else
            begin
              reg448 <= $unsigned((~^((+$unsigned(wire367)) ?
                  reg437[(4'h8):(3'h4)] : reg379)));
              reg449 = (~&$unsigned($unsigned(reg449)));
              reg450 <= reg415;
              reg451 = ($signed((~$unsigned(wire394))) ?
                  reg405 : {wire372[(2'h2):(1'h1)], (8'ha7)});
              reg452 = ($unsigned(wire393) ?
                  $signed(reg401[(5'h13):(2'h3)]) : {$signed(({wire368} ?
                          ((8'hbb) && reg438) : reg377[(4'hc):(4'hc)]))});
            end
          if ($unsigned($signed($signed($unsigned((^reg432))))))
            begin
              reg453 <= (8'hb2);
              reg454 = $unsigned(reg427[(1'h1):(1'h1)]);
              reg455 <= reg454;
              reg456 <= {{$unsigned((|reg390[(2'h3):(1'h0)])),
                      (((~|reg422) <<< (^forvar443)) ?
                          (^~{wire393, forvar426}) : ((reg373 ?
                              reg415 : reg374) + (forvar434 ?
                              wire424 : reg404)))},
                  (~reg387)};
              reg457 <= $unsigned(wire371[(2'h2):(1'h1)]);
            end
          else
            begin
              reg453 <= ((~&(($unsigned(reg386) * (reg455 >= reg438)) <= ((reg442 | reg432) > (reg415 == reg448)))) + $unsigned(((~(reg433 ?
                      reg422 : (8'h9e))) ?
                  (reg437 * reg428) : $signed(((8'ha5) ? reg377 : (8'h9d))))));
              reg454 = $signed(({$signed((wire366 ? wire367 : wire370)),
                      ($unsigned(forvar445) == (~|reg437))} ?
                  reg415 : ($unsigned((&wire366)) << (^reg401))));
              reg455 <= (reg453[(1'h0):(1'h0)] != $signed({($signed((8'ha4)) ?
                      $unsigned(reg388) : (wire370 ? wire424 : reg409))}));
              reg458 = $unsigned($signed((($signed(reg440) ?
                  (wire391 ?
                      wire394 : (8'ha7)) : wire370[(3'h6):(2'h3)]) ^~ (!{reg441,
                  wire366}))));
            end
        end
    end
  assign wire459 = (((~wire367[(2'h2):(1'h1)]) * (wire365 ?
                           wire366[(3'h5):(3'h4)] : (reg390[(4'hb):(3'h7)] ?
                               $signed(wire393) : reg409[(4'he):(1'h1)]))) ?
                       wire365 : (8'hbd));
  assign wire460 = reg381;
endmodule