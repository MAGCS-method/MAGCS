(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'hb2a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire3;
  input wire [(5'h1c):(1'h0)] wire2;
  input wire signed [(5'h15):(1'h0)] wire1;
  input wire [(5'h17):(1'h0)] wire0;
  wire signed [(3'h7):(1'h0)] wire222;
  wire signed [(4'hc):(1'h0)] wire90;
  wire [(4'hd):(1'h0)] wire89;
  wire signed [(5'h10):(1'h0)] wire4;
  wire signed [(5'h19):(1'h0)] wire2119;
  wire [(5'h14):(1'h0)] wire2196;
  wire signed [(3'h4):(1'h0)] wire2197;
  reg signed [(3'h7):(1'h0)] reg7 = (1'h0);
  reg [(5'h19):(1'h0)] reg8 = (1'h0);
  reg [(4'hb):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg10 = (1'h0);
  reg [(4'hd):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg13 = (1'h0);
  reg [(5'h13):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg19 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg25 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg34 = (1'h0);
  reg [(4'hb):(1'h0)] reg35 = (1'h0);
  reg [(5'h12):(1'h0)] reg37 = (1'h0);
  reg [(4'hc):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg40 = (1'h0);
  reg [(5'h17):(1'h0)] reg42 = (1'h0);
  reg [(5'h19):(1'h0)] reg44 = (1'h0);
  reg [(5'h1c):(1'h0)] reg45 = (1'h0);
  reg [(4'hd):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg49 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg54 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg56 = (1'h0);
  reg [(3'h7):(1'h0)] reg58 = (1'h0);
  reg [(5'h18):(1'h0)] reg64 = (1'h0);
  reg [(5'h1d):(1'h0)] reg65 = (1'h0);
  reg [(4'he):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg68 = (1'h0);
  reg [(4'ha):(1'h0)] reg73 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg77 = (1'h0);
  reg [(5'h18):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg75 = (1'h0);
  reg [(3'h7):(1'h0)] reg85 = (1'h0);
  reg [(5'h15):(1'h0)] reg2121 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2123 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2124 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2128 = (1'h0);
  reg [(4'hd):(1'h0)] reg2129 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2131 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2133 = (1'h0);
  reg [(5'h19):(1'h0)] reg2134 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2137 = (1'h0);
  reg [(3'h4):(1'h0)] reg2138 = (1'h0);
  reg [(4'hb):(1'h0)] reg2140 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2144 = (1'h0);
  reg [(2'h2):(1'h0)] reg2145 = (1'h0);
  reg [(3'h5):(1'h0)] reg2149 = (1'h0);
  reg [(4'hf):(1'h0)] reg2151 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2152 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2153 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2158 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2159 = (1'h0);
  reg [(3'h5):(1'h0)] reg2160 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2162 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2167 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2170 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2175 = (1'h0);
  reg [(4'hd):(1'h0)] reg2177 = (1'h0);
  reg [(4'h9):(1'h0)] reg2179 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2180 = (1'h0);
  reg [(4'h8):(1'h0)] reg2181 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2182 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2183 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2184 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2186 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2187 = (1'h0);
  reg [(5'h10):(1'h0)] reg2190 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2191 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2193 = (1'h0);
  reg [(5'h17):(1'h0)] reg2195 = (1'h0);
  reg [(5'h14):(1'h0)] reg2194 = (1'h0);
  reg [(5'h10):(1'h0)] reg2192 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2189 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2188 = (1'h0);
  reg [(4'he):(1'h0)] reg2185 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2178 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2176 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2174 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2173 = (1'h0);
  reg [(5'h15):(1'h0)] reg2172 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2171 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2169 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2168 = (1'h0);
  reg [(2'h2):(1'h0)] reg2166 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2165 = (1'h0);
  reg [(3'h5):(1'h0)] reg2164 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2163 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar2161 = (1'h0);
  reg [(5'h17):(1'h0)] reg2150 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2157 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2156 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2155 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2154 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2150 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2148 = (1'h0);
  reg [(5'h18):(1'h0)] reg2147 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2146 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2143 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2142 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2141 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2139 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2136 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2135 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2132 = (1'h0);
  reg [(3'h7):(1'h0)] reg2130 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2127 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2126 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2125 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2122 = (1'h0);
  reg [(3'h7):(1'h0)] reg88 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg87 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg84 = (1'h0);
  reg [(5'h14):(1'h0)] reg83 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg82 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg80 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg79 = (1'h0);
  reg [(5'h1b):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg76 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar75 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg72 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg71 = (1'h0);
  reg [(4'hd):(1'h0)] reg70 = (1'h0);
  reg signed [(4'he):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg66 = (1'h0);
  reg [(5'h1c):(1'h0)] reg63 = (1'h0);
  reg [(3'h6):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg61 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg60 = (1'h0);
  reg [(5'h18):(1'h0)] reg59 = (1'h0);
  reg [(5'h1c):(1'h0)] reg57 = (1'h0);
  reg [(5'h17):(1'h0)] reg55 = (1'h0);
  reg [(4'ha):(1'h0)] reg53 = (1'h0);
  reg [(4'h8):(1'h0)] forvar48 = (1'h0);
  reg [(5'h1f):(1'h0)] reg51 = (1'h0);
  reg [(5'h16):(1'h0)] reg50 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg43 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg41 = (1'h0);
  reg [(5'h1d):(1'h0)] reg38 = (1'h0);
  reg signed [(4'he):(1'h0)] reg36 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg33 = (1'h0);
  reg [(5'h17):(1'h0)] forvar32 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5 = (1'h0);
  reg [(3'h6):(1'h0)] reg31 = (1'h0);
  reg [(5'h1a):(1'h0)] reg30 = (1'h0);
  reg [(5'h1b):(1'h0)] reg29 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg28 = (1'h0);
  reg [(5'h10):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg23 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg20 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg16 = (1'h0);
  reg signed [(4'he):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg12 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6 = (1'h0);
  reg [(4'hd):(1'h0)] reg5 = (1'h0);
  assign y = {wire222,
                 wire90,
                 wire89,
                 wire4,
                 wire2119,
                 wire2196,
                 wire2197,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg13,
                 reg14,
                 reg18,
                 reg19,
                 reg21,
                 reg24,
                 reg25,
                 reg26,
                 reg34,
                 reg35,
                 reg37,
                 reg39,
                 reg40,
                 reg42,
                 reg44,
                 reg45,
                 reg48,
                 reg49,
                 reg52,
                 reg54,
                 reg56,
                 reg58,
                 reg64,
                 reg65,
                 reg67,
                 reg68,
                 reg73,
                 reg74,
                 reg77,
                 reg81,
                 reg75,
                 reg85,
                 reg2121,
                 reg2123,
                 reg2124,
                 reg2128,
                 reg2129,
                 reg2131,
                 reg2133,
                 reg2134,
                 reg2137,
                 reg2138,
                 reg2140,
                 reg2144,
                 reg2145,
                 reg2149,
                 reg2151,
                 reg2152,
                 reg2153,
                 reg2158,
                 reg2159,
                 reg2160,
                 reg2162,
                 reg2167,
                 reg2170,
                 reg2175,
                 reg2177,
                 reg2179,
                 reg2180,
                 reg2181,
                 reg2182,
                 reg2183,
                 reg2184,
                 reg2186,
                 reg2187,
                 reg2190,
                 reg2191,
                 reg2193,
                 reg2195,
                 reg2194,
                 reg2192,
                 forvar2189,
                 forvar2188,
                 reg2185,
                 reg2178,
                 reg2176,
                 reg2174,
                 reg2173,
                 reg2172,
                 reg2171,
                 forvar2169,
                 reg2168,
                 reg2166,
                 reg2165,
                 reg2164,
                 reg2163,
                 forvar2161,
                 reg2150,
                 reg2157,
                 reg2156,
                 forvar2155,
                 reg2154,
                 forvar2150,
                 forvar2148,
                 reg2147,
                 forvar2146,
                 reg2143,
                 reg2142,
                 reg2141,
                 reg2139,
                 reg2136,
                 reg2135,
                 reg2132,
                 reg2130,
                 reg2127,
                 reg2126,
                 reg2125,
                 reg2122,
                 reg88,
                 reg87,
                 reg86,
                 reg84,
                 reg83,
                 reg82,
                 reg80,
                 reg79,
                 reg78,
                 reg76,
                 forvar75,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg66,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg57,
                 reg55,
                 reg53,
                 forvar48,
                 reg51,
                 reg50,
                 reg47,
                 reg46,
                 reg43,
                 reg41,
                 reg38,
                 reg36,
                 reg33,
                 forvar32,
                 forvar5,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg23,
                 reg22,
                 reg20,
                 reg17,
                 reg16,
                 reg15,
                 reg12,
                 reg6,
                 reg5,
                 (1'h0)};
  assign wire4 = $unsigned((!wire2[(5'h10):(2'h3)]));
  always
    @(posedge clk) begin
      if (wire0)
        begin
          if ((wire4 > wire3))
            begin
              reg5 = (~$unsigned(((wire1[(5'h12):(2'h2)] ?
                      (wire3 * wire3) : (^~wire2)) ?
                  wire4[(3'h5):(1'h1)] : $unsigned((wire1 * wire4)))));
              reg6 = $unsigned((({((8'haa) <<< wire3), (reg5 > wire4)} ?
                  $unsigned($unsigned(reg5)) : ((wire4 ? wire1 : wire1) ?
                      reg5[(4'h8):(2'h2)] : $signed(wire3))) * (^~wire3)));
            end
          else
            begin
              reg7 <= {(~^(^(~$unsigned(reg6)))),
                  (~^wire0[(1'h1):(1'h1)]),
                  $unsigned(wire4)};
              reg8 <= (($unsigned((~(8'ha4))) ?
                  (!$unsigned($unsigned(reg7))) : $signed(($signed(reg7) ^ wire4[(4'he):(4'hd)]))) < (wire1 ?
                  (^~((wire2 >>> (8'ha0)) ?
                      $unsigned(wire1) : $signed(wire2))) : wire4[(4'ha):(4'ha)]));
              reg9 <= $signed({$signed(($signed(reg7) ?
                      wire0[(5'h14):(5'h11)] : $unsigned(wire4))),
                  $signed(($unsigned((8'hbb)) && wire4)),
                  {(wire2[(4'hf):(1'h0)] ? $signed(reg6) : ((8'hb1) <= reg8)),
                      (wire1 ? reg5[(4'hb):(2'h2)] : (reg7 ? reg5 : (8'hb8))),
                      wire0}});
              reg10 <= ((~wire0[(2'h2):(2'h2)]) ?
                  $unsigned($unsigned($unsigned((wire1 >> wire0)))) : ($unsigned((~wire1[(4'hb):(3'h5)])) >>> reg9));
              reg11 <= ($signed(((^$unsigned((8'hbb))) > $signed(wire1[(1'h0):(1'h0)]))) ?
                  ({reg8[(2'h3):(1'h0)], (7'h55), $signed(reg10)} ?
                      $unsigned(($signed(wire1) | reg8)) : wire4[(4'he):(1'h0)]) : reg7[(1'h1):(1'h0)]);
              reg12 = reg9;
              reg13 <= (~(wire3 ?
                  ($signed(reg7) || (reg9[(4'h9):(3'h6)] ?
                      (reg8 & wire2) : {wire3, wire2, wire4})) : (-(reg10 ?
                      $signed(reg6) : $unsigned(reg12)))));
            end
          reg14 <= ($unsigned($signed($unsigned(wire4))) << wire2[(5'h13):(5'h13)]);
          if (wire0[(4'h8):(3'h4)])
            begin
              reg15 = {$signed(reg8),
                  ((((~^reg14) ? (wire3 * reg13) : $unsigned(wire2)) ?
                          (7'h51) : $signed((|reg8))) ?
                      $unsigned((reg12 >> (reg14 >= reg11))) : (!reg10[(2'h3):(1'h1)])),
                  $unsigned(({(+reg9), {wire4}} ?
                      ($signed(wire4) ? reg6 : {(8'h9e), (7'h4c)}) : reg12))};
              reg16 = (~|($unsigned($unsigned(reg5)) <<< $unsigned((~^(wire2 * reg15)))));
              reg17 = $unsigned(wire0[(4'ha):(4'h8)]);
            end
          else
            begin
              reg18 <= (wire3[(3'h4):(1'h0)] ^ $unsigned(((reg7 <= $unsigned((8'ha7))) < (~&wire3))));
              reg19 <= ({$signed((reg12 | (reg11 ? reg13 : reg15))),
                  $unsigned($unsigned((8'ha9)))} && $unsigned((((8'ha5) >>> $signed((8'hb1))) >> $unsigned((reg9 ?
                  (7'h53) : reg8)))));
              reg20 = reg17[(1'h1):(1'h0)];
              reg21 <= ($unsigned({$unsigned((wire1 ? reg7 : reg9)),
                  ((~reg10) & (reg20 ? (8'hbc) : reg5)),
                  (wire4[(4'h8):(3'h7)] >= (reg6 || reg17))}) >= {reg12,
                  ($signed((wire0 && (8'hbc))) ?
                      ($signed(reg20) ? wire4 : (~&reg17)) : reg20),
                  (8'hab)});
              reg22 = {((8'h9f) << reg15)};
            end
          reg23 = $unsigned($signed({(reg6[(4'h9):(1'h0)] ?
                  ((7'h41) ? reg15 : reg12) : ((8'hb4) ? wire3 : reg7)),
              ((~|reg10) ? (|reg19) : ((8'ha7) ? reg5 : reg19)),
              wire0[(3'h4):(1'h0)]}));
          if ($unsigned((((~&reg16[(2'h2):(2'h2)]) <= wire1) ?
              $unsigned(reg16[(1'h1):(1'h1)]) : (~&(&((8'h9d) < reg14))))))
            begin
              reg24 <= (7'h4c);
            end
          else
            begin
              reg24 <= (8'hbc);
              reg25 <= (7'h44);
              reg26 <= (7'h42);
              reg27 = ((((^$unsigned(reg8)) ?
                          ($unsigned(reg14) < (reg11 - reg13)) : reg6) ?
                      (8'ha4) : $signed((~|$signed(wire3)))) ?
                  $unsigned(reg6[(4'hc):(3'h6)]) : (&(~^reg7)));
              reg28 = (8'hbb);
              reg29 = (reg6 | reg20[(5'h10):(2'h3)]);
            end
          reg30 = ((+(~&($signed(reg11) >>> reg10))) || reg23[(3'h4):(3'h4)]);
          reg31 = (8'h9d);
        end
      else
        begin
          for (forvar5 = (1'h0); (forvar5 < (3'h4)); forvar5 = (forvar5 + (1'h1)))
            begin
              reg7 <= (reg31[(1'h0):(1'h0)] ?
                  (($signed($signed(reg13)) ?
                      (7'h4a) : $signed({reg6})) << ({$signed(wire3),
                      (reg17 | wire1),
                      (7'h44)} >= $signed(reg19[(5'h17):(2'h3)]))) : (^((reg11[(4'h8):(2'h3)] >> {reg10,
                          (8'hb6)}) ?
                      reg7 : (+(-wire3)))));
            end
        end
      for (forvar32 = (1'h0); (forvar32 < (3'h6)); forvar32 = (forvar32 + (1'h1)))
        begin
          reg33 = ($unsigned(reg15[(4'ha):(4'ha)]) > $unsigned({{(reg9 == wire3),
                  reg13[(1'h1):(1'h0)],
                  (&reg16)},
              $signed(reg12),
              ((reg26 ? reg7 : reg12) + (reg17 ? reg8 : (7'h56)))}));
          reg34 <= (^wire3[(1'h0):(1'h0)]);
          if ((($signed(reg31) ?
                  (|($signed(reg5) ?
                      forvar32[(4'hc):(3'h4)] : {reg33})) : $signed(({reg21,
                          reg8,
                          reg21} ?
                      $unsigned(forvar32) : $signed(reg34)))) ?
              ($signed($unsigned((wire3 ~^ reg16))) ?
                  $unsigned((7'h51)) : $unsigned(($signed(reg8) && $signed(reg10)))) : $unsigned(($unsigned(((8'ha8) ?
                  reg13 : (7'h41))) <= ({reg17, forvar5} > $unsigned(reg20))))))
            begin
              reg35 <= {reg25[(4'he):(3'h5)],
                  $unsigned(forvar5[(3'h6):(3'h4)])};
              reg36 = $unsigned((($unsigned((~^reg33)) <<< $unsigned($signed(reg33))) ?
                  (~(^(reg27 >= reg29))) : $signed(reg28)));
              reg37 <= ((reg9[(1'h0):(1'h0)] >>> (forvar5[(3'h4):(3'h4)] ?
                  (~(reg11 == (7'h4f))) : (reg30 - (~&(7'h45))))) & $signed($unsigned(({reg23,
                      reg20,
                      wire2} ?
                  reg30[(4'hb):(4'h8)] : (reg33 ? reg15 : reg29)))));
              reg38 = ((~{($signed(reg35) ? {reg29, wire3} : $signed((7'h56))),
                  (~&(7'h51)),
                  $unsigned((reg19 ? (8'ha3) : reg9))}) >> (+$unsigned({reg27,
                  (reg36 ^ reg34),
                  $unsigned(reg33)})));
              reg39 <= (8'haa);
              reg40 <= $signed($signed(reg8));
              reg41 = ({{((~|reg24) ? (~|wire3) : ((7'h49) ? wire4 : reg6))},
                  (^(reg17 ? $signed((8'ha2)) : (reg8 || wire4))),
                  {reg12,
                      {(wire3 | reg9), (&reg26), $signed(reg25)},
                      {(reg18 ?
                              reg36 : (8'had))}}} >>> (reg11[(1'h1):(1'h1)] >= {$unsigned((reg7 ?
                      forvar5 : wire4)),
                  (|$unsigned(reg33))}));
            end
          else
            begin
              reg35 <= {reg37, reg21, {$unsigned(reg33[(1'h1):(1'h1)])}};
              reg36 = $signed((reg28 << ((~^$signed(reg11)) * {$unsigned(forvar5),
                  $signed(wire0)})));
              reg38 = reg24[(5'h16):(5'h14)];
            end
        end
      reg42 <= ((reg39[(4'hb):(4'ha)] ?
              (!reg5) : (({reg15} - $unsigned(reg35)) < (!reg30))) ?
          (|$signed($signed($unsigned(reg22)))) : $signed((reg35[(2'h2):(1'h0)] ?
              $unsigned(reg11[(4'ha):(1'h1)]) : ((~&reg35) > reg37[(3'h4):(1'h1)]))));
      if ($unsigned($signed({$unsigned($unsigned((8'hb7))),
          (^reg18[(3'h7):(1'h1)]),
          (8'hba)})))
        begin
          if ((~^{(((reg9 ? reg33 : reg34) || (~&reg9)) ?
                  $unsigned($unsigned(reg35)) : ((8'hbf) <<< reg38)),
              ($unsigned((reg14 ? reg38 : reg33)) || ($unsigned(reg20) ?
                  reg5 : $unsigned(reg14))),
              forvar32}))
            begin
              reg43 = (~(reg16 >= (~^$signed(reg19[(3'h5):(3'h4)]))));
              reg44 <= $unsigned(((reg30 ?
                      $unsigned((reg7 ?
                          reg36 : reg39)) : (~&$unsigned(wire1))) ?
                  reg29[(4'he):(1'h1)] : $unsigned({(~^reg42)})));
              reg45 <= reg35[(3'h7):(3'h4)];
              reg46 = (~|(reg33[(2'h2):(2'h2)] ? $unsigned(reg25) : (8'hb8)));
              reg47 = (((reg26[(1'h1):(1'h0)] ?
                      ((reg25 ? reg10 : reg28) ?
                          (wire1 < reg28) : (reg19 ? reg30 : reg25)) : {reg39,
                          (reg35 ? wire2 : reg15)}) - wire3) ?
                  {reg28, wire3[(3'h6):(2'h2)]} : $unsigned($signed((&reg36))));
              reg48 <= reg37;
              reg49 <= (!(8'hb1));
            end
          else
            begin
              reg44 <= (~$unsigned(reg21[(4'hc):(4'hc)]));
              reg46 = ({reg13,
                      reg8[(1'h1):(1'h1)],
                      (^$unsigned(((8'hbe) <<< reg14)))} ?
                  forvar5[(2'h3):(1'h0)] : (({(~&(7'h53)), (!reg17)} ?
                      (reg19[(4'he):(3'h6)] != (reg41 * reg27)) : reg8[(4'hf):(3'h4)]) >>> $signed(((reg38 << reg21) ?
                      $signed(forvar5) : (reg40 < reg9)))));
              reg47 = $signed(forvar32);
              reg50 = {({{$unsigned(reg29),
                          $signed(reg46),
                          reg16[(3'h5):(2'h3)]}} & (~|{$signed(wire0)})),
                  (((~|{reg16, reg46}) ?
                      wire4[(3'h4):(2'h3)] : ((reg46 <<< reg22) || (reg25 ^~ (7'h40)))) || (&({reg23,
                      reg24} <<< reg27[(3'h5):(2'h3)])))};
              reg51 = (!$unsigned((({reg7, forvar32} ?
                      {reg11} : reg49[(3'h6):(2'h2)]) ?
                  $signed((reg30 >>> reg17)) : (reg45 ?
                      (~(8'hb3)) : (^~reg14)))));
            end
          reg52 <= ({reg33[(1'h1):(1'h0)]} ?
              (7'h41) : {(reg15 ?
                      {reg28[(2'h3):(2'h3)],
                          (+wire3)} : ((reg38 << reg38) || wire0)),
                  (~|$unsigned({wire0, reg25, reg16})),
                  (^~((8'hb2) ? {reg35, reg40} : $signed(reg17)))});
        end
      else
        begin
          reg44 <= (~^(wire1 ? (-reg50) : $signed($signed($unsigned(reg40)))));
          reg46 = (({reg28[(1'h1):(1'h1)],
                  (reg6[(3'h4):(1'h1)] ? $signed(reg21) : ((8'ha9) > reg30)),
                  reg14} ?
              $signed((~|reg27[(4'he):(2'h3)])) : ($unsigned((reg31 ?
                      forvar32 : reg9)) ?
                  reg20[(5'h1a):(3'h4)] : reg42)) <= reg31[(1'h0):(1'h0)]);
          reg47 = (|((~(8'ha5)) != (8'hb3)));
          for (forvar48 = (1'h0); (forvar48 < (3'h4)); forvar48 = (forvar48 + (1'h1)))
            begin
              reg49 <= reg7;
              reg52 <= $signed((&(($signed((8'had)) > forvar48) ?
                  reg48 : (7'h49))));
              reg53 = reg8[(4'h9):(3'h5)];
              reg54 <= ({{$unsigned((reg11 << reg30)),
                      forvar32[(5'h10):(4'hc)],
                      ($unsigned(reg53) * (reg38 ? reg27 : forvar48))},
                  wire1,
                  (&reg26[(1'h1):(1'h0)])} | $signed($signed(({reg43,
                  reg7,
                  reg20} << (~|reg21)))));
              reg55 = ($signed($signed($unsigned(reg36))) ?
                  ($signed($signed($unsigned(wire0))) - {$unsigned((~reg28)),
                      (~^$unsigned(reg18)),
                      reg27[(3'h4):(3'h4)]}) : reg41);
              reg56 <= wire4[(4'ha):(4'h9)];
            end
          reg57 = (({($signed(forvar48) ? (|reg55) : reg50),
                  (reg53 ? (~|reg38) : wire0[(4'hb):(2'h2)]),
                  ($signed(reg21) ?
                      {reg8} : $signed(reg26))} - {reg13[(3'h7):(2'h3)],
                  ((reg56 ? reg53 : (8'hb0)) ?
                      (reg55 - forvar48) : reg36[(1'h1):(1'h0)])}) ?
              $unsigned($signed((~|$unsigned(reg18)))) : (reg26[(2'h2):(1'h1)] ?
                  $unsigned($signed(((8'h9d) ^~ reg34))) : reg22));
          reg58 <= reg14;
        end
      reg59 = $signed(($unsigned($unsigned((reg13 ?
          reg33 : reg26))) * reg24[(4'hd):(1'h0)]));
      reg60 = (~^$signed(($signed((reg55 ?
          reg20 : (7'h47))) ~^ reg49[(5'h14):(4'hf)])));
      reg61 = $signed((8'ha6));
    end
  always
    @(posedge clk) begin
      reg62 = (reg40[(4'hb):(4'h8)] ?
          (~reg34) : ({$unsigned($unsigned((8'h9f)))} <= (($unsigned(reg26) ?
              reg54[(4'hc):(4'hb)] : (^reg45)) | reg39[(4'ha):(4'ha)])));
      reg63 = {(|(((reg39 ? reg49 : reg42) ^~ (reg45 ? reg39 : reg21)) ?
              reg40 : $unsigned((8'haf)))),
          $signed(reg49[(4'hc):(1'h0)])};
      if (reg49[(4'hb):(4'h9)])
        begin
          reg64 <= $signed(reg45[(4'hd):(3'h5)]);
          reg65 <= reg62;
          if ($unsigned($unsigned(((reg18[(1'h1):(1'h1)] == (reg10 ?
                  reg44 : reg11)) ?
              reg21[(2'h3):(1'h0)] : $signed((wire4 ? (7'h42) : (8'hbe)))))))
            begin
              reg66 = (((+wire1) ?
                      reg21[(1'h0):(1'h0)] : reg19[(3'h4):(1'h1)]) ?
                  $unsigned(reg42[(4'h9):(2'h3)]) : $signed(reg37));
              reg67 <= ($signed((!$unsigned({wire2, reg49}))) ?
                  $unsigned($signed(reg45[(4'hc):(3'h7)])) : (reg34 ?
                      wire1 : (&{(reg44 * reg21), $signed(wire2)})));
              reg68 <= {$unsigned((7'h42))};
            end
          else
            begin
              reg66 = reg40[(4'h8):(2'h3)];
              reg67 <= reg67;
              reg69 = $signed(reg39);
              reg70 = ({(reg25 ~^ $signed((reg14 <= (8'ha4))))} ?
                  ((^~reg35[(4'h8):(3'h7)]) ?
                      reg67 : (reg62[(2'h2):(1'h0)] >= (7'h55))) : $signed((reg66[(3'h6):(2'h3)] ?
                      ({wire1, (7'h57)} ?
                          reg65 : wire0) : (reg62[(2'h3):(1'h0)] ?
                          reg64 : reg62[(3'h4):(2'h3)]))));
              reg71 = wire3[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg64 <= reg9[(1'h1):(1'h1)];
          reg65 <= wire4[(4'h9):(3'h4)];
          reg66 = $unsigned(reg14[(4'h8):(4'h8)]);
        end
      if ($unsigned(wire2[(4'hf):(4'hb)]))
        begin
          reg72 = {$signed(reg11[(2'h2):(1'h0)])};
          reg73 <= ((7'h40) << reg8);
          reg74 <= ((wire4 ?
                  reg70[(3'h4):(3'h4)] : $unsigned(({reg34, reg8} ?
                      ((7'h49) ? reg45 : reg34) : (-reg11)))) ?
              (reg39[(3'h6):(1'h1)] ?
                  ((((7'h45) ? reg58 : reg49) ? $signed(reg49) : (&reg44)) ?
                      {(reg42 ? wire3 : reg14),
                          $signed(reg68),
                          (reg68 > reg73)} : ($unsigned((8'hbd)) ?
                          $signed(reg13) : reg56)) : $signed((+reg56[(3'h7):(3'h5)]))) : (($unsigned($unsigned(reg14)) ?
                  reg21 : $unsigned(reg25)) * reg68[(1'h0):(1'h0)]));
          for (forvar75 = (1'h0); (forvar75 < (1'h0)); forvar75 = (forvar75 + (1'h1)))
            begin
              reg76 = ($unsigned($unsigned(reg63)) != $unsigned({$unsigned(reg73[(4'h9):(3'h7)]),
                  ($signed(reg64) >> (8'hba)),
                  $signed($signed(reg9))}));
              reg77 <= ($unsigned((($signed(reg26) ? wire0 : $unsigned(reg11)) ?
                  wire4[(3'h6):(2'h2)] : (reg9[(2'h3):(1'h1)] & (8'ha0)))) ~^ reg8[(4'h9):(2'h3)]);
            end
          if (reg54)
            begin
              reg78 = $signed($signed((|((reg40 ?
                  (8'hb8) : forvar75) ^ {reg58}))));
              reg79 = wire1[(4'hb):(3'h7)];
              reg80 = $signed(reg67[(4'h9):(2'h3)]);
              reg81 <= (reg45 ?
                  ($unsigned(wire4) ?
                      (reg73 ?
                          (^$unsigned(reg65)) : ((~reg63) ?
                              (^reg14) : (forvar75 ?
                                  reg21 : reg67))) : {((reg18 ?
                                  (7'h44) : reg7) ?
                              $signed(reg67) : (reg69 <= wire0)),
                          (7'h4a),
                          ($unsigned((8'ha5)) ?
                              (8'ha9) : (~^reg34))}) : (^$unsigned((~^(8'had)))));
              reg82 = reg74;
            end
          else
            begin
              reg78 = reg10[(4'hc):(4'h8)];
              reg79 = (~&$signed(wire1));
              reg81 <= $unsigned(((reg49 ?
                      ($signed(reg35) && $unsigned(reg80)) : $signed((reg14 ?
                          wire4 : reg63))) ?
                  reg25 : (~$unsigned((reg71 ^ (8'haf))))));
              reg82 = reg8[(1'h1):(1'h1)];
              reg83 = reg39[(3'h5):(2'h2)];
            end
        end
      else
        begin
          reg73 <= {reg10};
          reg74 <= wire0;
          if ((~|$signed($signed((~(|reg82))))))
            begin
              reg75 <= $signed(reg70[(1'h0):(1'h0)]);
              reg76 = $signed(($unsigned((8'hbe)) ? (~|reg24) : reg79));
              reg78 = (~{$signed({(&reg80), reg19[(5'h16):(1'h1)]})});
              reg81 <= (+($unsigned(reg79) < (~&((reg82 ?
                  reg34 : reg69) + $signed(wire4)))));
              reg82 = $unsigned($unsigned(($unsigned($unsigned(reg37)) ?
                  (^~reg70[(2'h2):(2'h2)]) : (^reg34))));
              reg83 = $unsigned($unsigned(reg44[(5'h14):(4'h8)]));
              reg84 = wire1[(4'ha):(1'h0)];
            end
          else
            begin
              reg76 = ($unsigned((reg48[(4'h9):(4'h9)] >= reg19)) ?
                  (^~(reg13[(3'h7):(1'h1)] ?
                      reg84[(5'h11):(4'hf)] : (~|reg13[(1'h0):(1'h0)]))) : $unsigned((!(+(~&(8'hae))))));
              reg78 = reg68[(3'h4):(3'h4)];
              reg81 <= {{$signed((7'h4e)),
                      {((reg14 && reg79) ?
                              reg48[(3'h6):(3'h5)] : (reg56 ? reg18 : reg9))}}};
              reg85 <= wire1[(2'h3):(2'h2)];
              reg86 = $unsigned((-reg56[(5'h1a):(5'h16)]));
            end
          reg87 = reg19[(5'h15):(1'h0)];
          reg88 = $unsigned((-(-({reg62} | reg69[(4'hb):(4'ha)]))));
        end
    end
  assign wire89 = (($unsigned(((reg7 ^~ reg11) ?
                              reg73[(3'h6):(3'h6)] : reg52[(4'hb):(4'hb)])) ?
                          {$unsigned(reg11[(4'hc):(4'h8)]),
                              {$unsigned(reg39), (reg75 + reg77), (|reg68)},
                              reg37[(3'h6):(1'h1)]} : (reg65[(4'hc):(2'h2)] ?
                              reg65 : ((reg67 ?
                                  reg42 : (8'h9c)) < $signed(wire2)))) ?
                      (~&$unsigned(((reg19 || reg35) ^~ (+reg21)))) : (~|$signed(((reg9 != wire0) - (reg37 ~^ reg18)))));
  assign wire90 = (($signed(reg40) ~^ (reg58[(3'h5):(3'h4)] && ((reg24 ?
                          reg35 : reg34) ?
                      (reg65 ?
                          wire3 : reg49) : $unsigned(reg25)))) * {((reg26 - (reg35 ?
                              wire4 : reg44)) ?
                          {reg42[(3'h7):(3'h4)]} : ((wire0 ? wire3 : reg45) ?
                              reg35 : $unsigned(reg58))),
                      ($unsigned((reg74 ? reg75 : wire1)) ?
                          $unsigned($unsigned(reg48)) : reg10)});
  module91 #() modinst223 (.wire94(reg11), .wire95(reg24), .y(wire222), .wire92(wire90), .wire96(reg85), .clk(clk), .wire93(reg34));
  module224 #() modinst2120 (.wire228(reg24), .y(wire2119), .wire226(reg75), .wire227(reg21), .wire225(reg81), .clk(clk));
  always
    @(posedge clk) begin
      if ($unsigned($unsigned((reg68 || ($signed(wire4) >>> (~&reg52))))))
        begin
          reg2121 <= $unsigned(reg21);
          if (((7'h56) ?
              {reg75[(4'hf):(3'h7)]} : $unsigned($unsigned(($unsigned(wire222) ?
                  reg52 : (wire222 || wire3))))))
            begin
              reg2122 = reg18[(1'h0):(1'h0)];
              reg2123 <= (((wire4 ? reg2122 : (~^reg45)) ?
                      $unsigned({{(8'ha6), (7'h58)},
                          $signed(reg73)}) : (^(~|wire4[(3'h4):(2'h2)]))) ?
                  $signed($signed($unsigned($unsigned(reg52)))) : (((reg85 > (reg65 ?
                      reg25 : reg9)) >>> ((reg39 <<< reg25) ?
                      (reg39 ?
                          wire89 : reg65) : (reg2122 >> reg34))) | (((reg8 ?
                              reg2122 : reg40) ?
                          (~|wire3) : wire2119[(5'h17):(5'h15)]) ?
                      (reg75[(5'h16):(3'h4)] ^ $unsigned((8'hb8))) : {(+reg21)})));
              reg2124 <= (((~&$signed(reg45)) ?
                      $unsigned($signed((~wire4))) : reg37) ?
                  $signed((({reg25, reg11} ?
                      (|(7'h52)) : (~wire4)) <<< $signed(reg54[(2'h2):(1'h0)]))) : wire2);
            end
          else
            begin
              reg2122 = (~|(wire90 ? reg45 : (8'hac)));
              reg2125 = reg40[(4'he):(1'h1)];
              reg2126 = (~^$signed(reg54));
            end
          if (reg2122[(3'h4):(2'h2)])
            begin
              reg2127 = (|$signed((8'hbd)));
              reg2128 <= $signed(({reg7[(3'h5):(3'h5)],
                  (^~reg65[(4'ha):(3'h6)])} & (reg19[(4'he):(4'h8)] ~^ reg18)));
              reg2129 <= ((reg14[(5'h11):(4'hc)] && ((^~reg21[(4'hd):(3'h7)]) < $unsigned((reg40 ~^ reg2122)))) != wire222);
              reg2130 = $unsigned(($signed((((8'ha7) & reg64) ?
                      reg48[(4'hc):(3'h6)] : $signed(reg11))) ?
                  ((wire0 ?
                      $signed((7'h56)) : $signed(reg18)) <<< reg67) : $signed((^~{reg42,
                      wire1,
                      (8'hb6)}))));
            end
          else
            begin
              reg2128 <= (~|reg77);
              reg2130 = reg26;
              reg2131 <= (+$signed((reg65[(3'h4):(2'h3)] ?
                  ((reg37 < reg85) ?
                      reg2125[(5'h12):(4'hf)] : (+wire4)) : (|(|wire90)))));
            end
          if ($signed(reg24[(5'h1c):(3'h6)]))
            begin
              reg2132 = (reg39[(2'h3):(2'h2)] * $unsigned(($unsigned((reg14 | reg18)) <= (~|reg7[(1'h0):(1'h0)]))));
              reg2133 <= $unsigned(($signed(((reg44 ? reg11 : reg40) ?
                  reg2124 : (reg44 >= (7'h49)))) <= ($signed(reg7[(3'h5):(3'h5)]) ?
                  $signed($signed(wire90)) : $unsigned($signed(reg14)))));
              reg2134 <= $signed(reg11[(4'hb):(3'h6)]);
              reg2135 = ({(|((^reg35) ? $unsigned(reg65) : $signed(reg42))),
                  reg68,
                  ((8'hb7) * (~&reg44))} == (|(reg2123[(5'h18):(5'h11)] > (reg2124[(3'h4):(2'h3)] - reg2122[(1'h1):(1'h1)]))));
              reg2136 = $unsigned(($signed(((reg34 ?
                      reg2135 : wire90) << reg74[(3'h6):(3'h6)])) ?
                  (~reg21[(2'h3):(1'h1)]) : (^~$signed($unsigned(reg54)))));
              reg2137 <= (^~$signed(reg2131[(3'h4):(3'h4)]));
              reg2138 <= (($unsigned($signed(wire3)) ?
                  reg49 : reg74) >>> ((|(reg48[(4'hd):(2'h2)] + (wire1 ?
                      reg40 : reg48))) ?
                  {(-(^~reg49)),
                      ((reg54 | reg40) ?
                          (reg42 ? reg73 : wire90) : {wire0,
                              reg54})} : (8'hbb)));
            end
          else
            begin
              reg2133 <= ((^(((reg2127 + reg77) ?
                          reg2129[(4'hd):(1'h0)] : (reg2132 ?
                              reg2135 : reg13)) ?
                      $unsigned({reg52, (8'hbf), reg2129}) : $unsigned({reg7,
                          wire1}))) ?
                  (wire0 ?
                      reg40 : {$unsigned((wire1 < (8'hab))),
                          $signed(reg21[(3'h4):(2'h3)])}) : $unsigned(($unsigned({reg2136,
                      (8'hbd),
                      reg37}) > $signed((reg75 - reg25)))));
              reg2135 = reg2130;
            end
          reg2139 = $unsigned(reg45);
        end
      else
        begin
          reg2121 <= (7'h58);
        end
      if (reg10[(4'hf):(4'h9)])
        begin
          reg2140 <= reg67[(4'he):(1'h1)];
        end
      else
        begin
          if (reg2138[(3'h4):(3'h4)])
            begin
              reg2140 <= (~&(reg2136 ?
                  (~^reg75) : (^$signed($unsigned(reg7)))));
            end
          else
            begin
              reg2141 = reg2138[(3'h4):(1'h0)];
              reg2142 = {reg2132};
              reg2143 = ((|$signed(reg21)) ?
                  $signed({(reg2142[(5'h14):(1'h1)] || (wire222 ?
                          reg14 : (8'hba))),
                      {$signed(reg44), $signed(reg9), {reg2134, (8'hbc)}},
                      reg11}) : (((+$signed(wire4)) ?
                      ($unsigned((8'hae)) ?
                          $signed(reg25) : (7'h4e)) : $unsigned($signed(reg24))) ^ (!($unsigned(reg2141) == $unsigned((7'h46))))));
              reg2144 <= $signed((~(reg2125 ^ {(reg2131 ? reg65 : (7'h55)),
                  reg19,
                  $signed(wire4)})));
              reg2145 <= ($signed($unsigned($unsigned((^(8'hb3))))) ?
                  (~|$unsigned(((reg2133 ? reg18 : reg81) ?
                      reg2131[(1'h0):(1'h0)] : (reg2144 <<< reg2139)))) : $signed($unsigned(($signed(reg21) ?
                      (7'h51) : reg67))));
            end
          for (forvar2146 = (1'h0); (forvar2146 < (2'h2)); forvar2146 = (forvar2146 + (1'h1)))
            begin
              reg2147 = ((|($unsigned((|reg2142)) ?
                      reg2126[(4'hd):(2'h2)] : reg34[(4'he):(2'h3)])) ?
                  reg8 : reg2127);
            end
        end
      for (forvar2148 = (1'h0); (forvar2148 < (3'h4)); forvar2148 = (forvar2148 + (1'h1)))
        begin
          reg2149 <= $signed(((~|$unsigned((+reg2127))) ?
              (&$signed((wire2119 ?
                  reg85 : reg11))) : $signed((+reg44[(4'h8):(2'h2)]))));
        end
      if (((+$signed(reg2123)) ?
          (($unsigned(reg52) * (&(!reg2145))) ?
              (7'h45) : {{$signed(reg2131),
                      $unsigned(wire90),
                      $unsigned(wire222)},
                  (+$signed(reg2143))}) : ($signed((~^reg45[(2'h3):(2'h3)])) ?
              $unsigned({(reg68 < reg7)}) : ({reg2140} ?
                  $unsigned($signed(reg11)) : reg2137))))
        begin
          for (forvar2150 = (1'h0); (forvar2150 < (3'h5)); forvar2150 = (forvar2150 + (1'h1)))
            begin
              reg2151 <= (reg2131 ? $signed(reg48) : (8'h9e));
              reg2152 <= (reg85 - $unsigned(wire222[(3'h7):(3'h5)]));
              reg2153 <= (reg52 ?
                  (($signed((~^reg2136)) ~^ $unsigned(((8'ha8) << (7'h48)))) ?
                      $unsigned(reg49) : (^wire4[(1'h0):(1'h0)])) : (7'h58));
              reg2154 = reg19;
            end
          for (forvar2155 = (1'h0); (forvar2155 < (3'h4)); forvar2155 = (forvar2155 + (1'h1)))
            begin
              reg2156 = reg2136;
              reg2157 = (($unsigned(($signed(reg2125) ?
                      $signed((7'h50)) : (reg48 ? reg2129 : reg25))) ?
                  ((reg45 ?
                      reg2141 : (reg81 == reg45)) >>> $signed((8'ha7))) : (reg21[(1'h1):(1'h0)] ?
                      (~|(^~reg26)) : $signed((reg74 ?
                          forvar2150 : reg21)))) == $unsigned(forvar2150[(4'he):(3'h6)]));
              reg2158 <= reg73;
              reg2159 <= wire89;
            end
        end
      else
        begin
          reg2150 = $signed($unsigned($signed($unsigned((~^reg77)))));
        end
    end
  always
    @(posedge clk) begin
      reg2160 <= (~^$signed(reg48));
      for (forvar2161 = (1'h0); (forvar2161 < (1'h0)); forvar2161 = (forvar2161 + (1'h1)))
        begin
          if (reg2138[(2'h2):(2'h2)])
            begin
              reg2162 <= $unsigned(reg18);
              reg2163 = $signed((reg48 > reg2160[(2'h3):(1'h1)]));
              reg2164 = (reg18[(1'h1):(1'h1)] || reg54);
              reg2165 = {$unsigned(reg85[(2'h3):(1'h0)]),
                  ((((reg65 ?
                      (7'h53) : (8'hbe)) <<< $unsigned((8'hb9))) ^ {(!wire90),
                      reg68}) && reg2134)};
              reg2166 = (~^((!reg2158) ^ ((^~(reg2123 - reg35)) - ($unsigned(reg85) ?
                  ((8'hbe) ? reg2123 : reg39) : {(7'h40)}))));
            end
          else
            begin
              reg2162 <= $unsigned(reg26[(1'h1):(1'h1)]);
              reg2167 <= reg2124;
              reg2168 = (^($unsigned((8'ha1)) == (+(((8'hac) ?
                  wire89 : (8'hb5)) >> {reg2144, reg85, wire2}))));
            end
        end
      for (forvar2169 = (1'h0); (forvar2169 < (1'h1)); forvar2169 = (forvar2169 + (1'h1)))
        begin
          if (reg81[(5'h15):(3'h7)])
            begin
              reg2170 <= reg39[(2'h2):(2'h2)];
            end
          else
            begin
              reg2171 = $signed(($signed({wire1, reg2138, reg2152}) ?
                  ($signed($signed(reg73)) ?
                      (~$unsigned(reg45)) : (((7'h50) ?
                          reg42 : (8'hab)) * (reg44 ?
                          wire3 : (7'h4a)))) : $signed(reg26[(1'h1):(1'h0)])));
            end
          reg2172 = reg37;
        end
      if ({wire2})
        begin
          reg2173 = $unsigned($signed((!reg68[(1'h1):(1'h1)])));
          reg2174 = ($signed(((reg8[(4'ha):(3'h7)] ?
                      {reg2128, reg2128} : reg21[(3'h4):(1'h0)]) ?
                  reg2145[(1'h1):(1'h1)] : (&reg19[(3'h5):(2'h2)]))) ?
              (wire2119 >= (~^(8'ha2))) : $signed($unsigned({{wire2119,
                      reg64,
                      reg45},
                  $signed(reg2163),
                  reg68})));
          reg2175 <= (reg2149 >= ({$signed(reg45),
                  ($signed(wire3) == (8'ha4))} ?
              reg21 : $unsigned($signed(reg2162[(5'h17):(2'h3)]))));
        end
      else
        begin
          reg2173 = {$unsigned((^~$signed({wire3})))};
          if (((($unsigned(reg49) ?
                      ((reg2129 || reg18) | ((8'hb5) + wire0)) : {reg2144[(2'h3):(1'h0)],
                          reg2166}) ?
                  {reg2158} : (!forvar2161[(2'h3):(2'h2)])) ?
              $signed(reg21[(3'h7):(3'h6)]) : (($unsigned(((8'h9d) || reg2128)) ?
                  reg68 : (reg2137[(1'h1):(1'h0)] ?
                      (reg10 | reg49) : reg35)) & reg34[(1'h1):(1'h0)])))
            begin
              reg2175 <= $unsigned((reg39[(1'h1):(1'h1)] ?
                  ((~|$signed((8'hb5))) * {(reg49 > (8'had)),
                      reg2171[(4'h8):(4'h8)]}) : $unsigned($unsigned($unsigned(reg75)))));
              reg2176 = reg73[(4'h8):(3'h7)];
              reg2177 <= (8'ha8);
            end
          else
            begin
              reg2175 <= $signed($unsigned($signed(($signed((7'h4f)) && reg2134[(5'h14):(1'h0)]))));
              reg2176 = $signed($unsigned((|reg81)));
              reg2178 = $unsigned($unsigned($signed(({(8'ha3), reg19} ?
                  (reg18 ? (8'hb1) : reg49) : wire2119))));
              reg2179 <= $signed(wire89[(3'h5):(1'h1)]);
            end
          if ($unsigned((reg75 && $unsigned($unsigned((|reg2158))))))
            begin
              reg2180 <= $signed(({$signed((~^reg2129))} | ((-(reg64 && reg2145)) & ($unsigned(reg52) ?
                  (wire4 * (7'h48)) : $unsigned((8'ha0))))));
              reg2181 <= reg2170[(4'hf):(2'h2)];
              reg2182 <= $signed(($signed($unsigned(((8'h9d) ?
                      (8'ha6) : reg37))) ?
                  {$unsigned({reg24,
                          reg58,
                          (7'h4e)})} : {reg2173[(3'h4):(1'h1)],
                      reg74[(1'h1):(1'h1)]}));
              reg2183 <= (^{(&$unsigned((reg65 - reg35)))});
              reg2184 <= $unsigned(((^reg2168[(2'h2):(1'h1)]) ?
                  reg2176[(4'hf):(2'h3)] : reg11[(3'h6):(3'h4)]));
            end
          else
            begin
              reg2185 = reg2170;
              reg2186 <= $signed(($signed(reg74) ?
                  reg2152[(5'h1b):(1'h0)] : $unsigned($unsigned((reg56 ~^ wire1)))));
            end
        end
      reg2187 <= $signed(($unsigned(reg2160) >>> (|(~&(|reg44)))));
      for (forvar2188 = (1'h0); (forvar2188 < (3'h6)); forvar2188 = (forvar2188 + (1'h1)))
        begin
          for (forvar2189 = (1'h0); (forvar2189 < (2'h2)); forvar2189 = (forvar2189 + (1'h1)))
            begin
              reg2190 <= ((8'ha7) ?
                  {{(^(reg2123 ? reg2179 : reg14))},
                      $unsigned($unsigned((reg2186 ?
                          (8'hac) : forvar2189)))} : ((!reg2149[(1'h0):(1'h0)]) + (((^reg2171) ?
                          {reg2165, reg68, reg2165} : reg2137) ?
                      (reg2124[(2'h2):(1'h0)] ?
                          {reg2124, (7'h50)} : {reg49,
                              wire222,
                              reg25}) : $signed($unsigned(reg2181)))));
              reg2191 <= reg42[(3'h6):(2'h3)];
              reg2192 = ((~&{reg2158[(3'h6):(1'h1)],
                  $unsigned($signed(reg2160)),
                  $unsigned((|reg77))}) ~^ reg2179);
              reg2193 <= ($signed({(~&(reg18 <= reg2129))}) ?
                  (($unsigned($unsigned(reg68)) ? reg2173 : (8'hb5)) ?
                      (~reg25) : (((~&reg2158) ? (7'h4e) : $signed(reg2158)) ?
                          (reg2191 | $signed((8'hbc))) : {(reg2176 >>> reg19)})) : ((~&reg2184[(3'h7):(3'h6)]) <<< $unsigned(reg40[(5'h10):(3'h5)])));
              reg2194 = $signed($signed(reg58[(1'h1):(1'h1)]));
            end
        end
      reg2195 = {(reg45 >= ($signed({reg2194, (7'h52), reg2191}) ?
              reg74 : reg18[(4'h9):(4'h9)])),
          $unsigned((|$signed($unsigned(reg2182)))),
          (^$unsigned((|$signed((8'hbe)))))};
    end
  assign wire2196 = reg2134;
  module100 #() modinst2198 (.wire103(reg8), .clk(clk), .wire104(reg2144), .wire101(reg2181), .y(wire2197), .wire102(wire1), .wire106(reg2133), .wire105(reg21));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module224
#(parameter param2118 = (&({(((7'h4b) != (7'h4a)) >> ((8'ha8) ? (7'h45) : (7'h49)))} ? (({(7'h42), (7'h4c), (7'h49)} && ((7'h4a) >= (8'h9e))) ? ((7'h4e) ? ((7'h57) ? (8'hb6) : (8'hb4)) : ((7'h48) ? (7'h55) : (7'h54))) : ({(7'h56), (8'hba)} ? ((8'ha4) < (8'hb8)) : ((8'hba) ? (8'h9f) : (7'h53)))) : ((8'h9e) != {(~&(7'h4c)), (-(8'haf))}))))
(y, clk, wire228, wire227, wire226, wire225);
  output wire [(32'h163c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire228;
  input wire [(4'hd):(1'h0)] wire227;
  input wire signed [(5'h17):(1'h0)] wire226;
  input wire [(5'h10):(1'h0)] wire225;
  wire [(4'he):(1'h0)] wire2098;
  wire signed [(5'h1e):(1'h0)] wire2000;
  wire signed [(3'h6):(1'h0)] wire1999;
  wire [(4'hf):(1'h0)] wire1997;
  wire signed [(5'h10):(1'h0)] wire319;
  wire [(2'h2):(1'h0)] wire293;
  wire signed [(3'h7):(1'h0)] wire292;
  wire signed [(2'h3):(1'h0)] wire291;
  wire signed [(5'h1d):(1'h0)] wire229;
  reg signed [(5'h1a):(1'h0)] reg2100 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2116 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2115 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2114 = (1'h0);
  reg [(2'h3):(1'h0)] reg2112 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2111 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2108 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2107 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2106 = (1'h0);
  reg [(4'hb):(1'h0)] reg2104 = (1'h0);
  reg [(3'h6):(1'h0)] reg2102 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2101 = (1'h0);
  reg [(5'h16):(1'h0)] reg2096 = (1'h0);
  reg [(3'h4):(1'h0)] reg2093 = (1'h0);
  reg [(3'h5):(1'h0)] reg2089 = (1'h0);
  reg [(4'he):(1'h0)] reg2085 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2084 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2083 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2065 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2082 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2080 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2079 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2078 = (1'h0);
  reg [(4'hc):(1'h0)] reg2076 = (1'h0);
  reg [(5'h11):(1'h0)] reg2074 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2072 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2071 = (1'h0);
  reg [(4'hc):(1'h0)] reg2067 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2066 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2064 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2063 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2062 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2060 = (1'h0);
  reg [(4'he):(1'h0)] reg2058 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2056 = (1'h0);
  reg [(5'h18):(1'h0)] reg2054 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2049 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2046 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2045 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2044 = (1'h0);
  reg [(4'hd):(1'h0)] reg2042 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2041 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2039 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2036 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2035 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2031 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2029 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2024 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2022 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2020 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2017 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2015 = (1'h0);
  reg [(3'h7):(1'h0)] reg2014 = (1'h0);
  reg [(5'h11):(1'h0)] reg2012 = (1'h0);
  reg [(4'hf):(1'h0)] reg2011 = (1'h0);
  reg [(4'h8):(1'h0)] reg2009 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2008 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2006 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2005 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2003 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2002 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2001 = (1'h0);
  reg [(3'h7):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg232 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg238 = (1'h0);
  reg [(4'he):(1'h0)] reg239 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg240 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg246 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg248 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg250 = (1'h0);
  reg [(5'h1e):(1'h0)] reg252 = (1'h0);
  reg [(5'h12):(1'h0)] reg253 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg257 = (1'h0);
  reg [(5'h1e):(1'h0)] reg262 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg273 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg274 = (1'h0);
  reg [(4'hb):(1'h0)] reg277 = (1'h0);
  reg [(4'hf):(1'h0)] reg279 = (1'h0);
  reg [(5'h10):(1'h0)] reg280 = (1'h0);
  reg [(5'h1e):(1'h0)] reg281 = (1'h0);
  reg [(4'he):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg284 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg295 = (1'h0);
  reg [(4'he):(1'h0)] reg296 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg299 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg301 = (1'h0);
  reg [(3'h7):(1'h0)] reg302 = (1'h0);
  reg [(5'h1b):(1'h0)] reg303 = (1'h0);
  reg [(2'h2):(1'h0)] reg304 = (1'h0);
  reg [(3'h4):(1'h0)] reg307 = (1'h0);
  reg [(4'ha):(1'h0)] reg311 = (1'h0);
  reg [(4'h8):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg314 = (1'h0);
  reg [(5'h1c):(1'h0)] reg316 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg320 = (1'h0);
  reg [(4'hc):(1'h0)] reg325 = (1'h0);
  reg [(5'h17):(1'h0)] reg327 = (1'h0);
  reg [(5'h13):(1'h0)] reg328 = (1'h0);
  reg [(5'h1a):(1'h0)] reg329 = (1'h0);
  reg [(5'h1f):(1'h0)] reg330 = (1'h0);
  reg [(5'h13):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg332 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg334 = (1'h0);
  reg [(4'h9):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg342 = (1'h0);
  reg [(5'h1a):(1'h0)] reg343 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg345 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg348 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg351 = (1'h0);
  reg [(3'h5):(1'h0)] reg353 = (1'h0);
  reg [(5'h10):(1'h0)] reg355 = (1'h0);
  reg [(4'ha):(1'h0)] reg358 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg371 = (1'h0);
  reg [(2'h2):(1'h0)] reg378 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg379 = (1'h0);
  reg [(5'h15):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg384 = (1'h0);
  reg [(4'ha):(1'h0)] reg385 = (1'h0);
  reg [(5'h1b):(1'h0)] reg388 = (1'h0);
  reg [(4'he):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg391 = (1'h0);
  reg [(5'h18):(1'h0)] reg392 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg394 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg397 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg400 = (1'h0);
  reg signed [(4'he):(1'h0)] reg401 = (1'h0);
  reg [(5'h1b):(1'h0)] reg403 = (1'h0);
  reg [(5'h11):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg405 = (1'h0);
  reg [(5'h1f):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg409 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg410 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg412 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg413 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg415 = (1'h0);
  reg [(4'hd):(1'h0)] reg417 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg420 = (1'h0);
  reg [(5'h1f):(1'h0)] reg421 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg423 = (1'h0);
  reg [(4'h8):(1'h0)] reg426 = (1'h0);
  reg [(3'h4):(1'h0)] reg430 = (1'h0);
  reg [(3'h6):(1'h0)] reg431 = (1'h0);
  reg signed [(4'he):(1'h0)] reg432 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2117 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2106 = (1'h0);
  reg [(4'hf):(1'h0)] reg2113 = (1'h0);
  reg [(3'h4):(1'h0)] reg2110 = (1'h0);
  reg [(5'h14):(1'h0)] reg2109 = (1'h0);
  reg [(4'ha):(1'h0)] reg2105 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2103 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar2100 = (1'h0);
  reg [(4'hc):(1'h0)] reg2099 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2097 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2095 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2094 = (1'h0);
  reg [(4'ha):(1'h0)] reg2092 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2091 = (1'h0);
  reg [(4'he):(1'h0)] reg2090 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2088 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2087 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2086 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2081 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar2076 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2073 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2064 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2081 = (1'h0);
  reg [(4'h8):(1'h0)] reg2077 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2075 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2073 = (1'h0);
  reg [(2'h2):(1'h0)] reg2070 = (1'h0);
  reg [(4'ha):(1'h0)] reg2069 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2068 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2065 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2061 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2059 = (1'h0);
  reg [(3'h6):(1'h0)] reg2057 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2055 = (1'h0);
  reg [(4'he):(1'h0)] reg2053 = (1'h0);
  reg [(5'h17):(1'h0)] reg2052 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2051 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2050 = (1'h0);
  reg [(5'h19):(1'h0)] reg2048 = (1'h0);
  reg [(5'h14):(1'h0)] reg2047 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2043 = (1'h0);
  reg [(3'h6):(1'h0)] reg2040 = (1'h0);
  reg [(2'h3):(1'h0)] reg2038 = (1'h0);
  reg [(5'h12):(1'h0)] reg2037 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2034 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2033 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2032 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar2030 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2028 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2027 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2026 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2025 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2023 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2021 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2019 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2018 = (1'h0);
  reg [(4'hb):(1'h0)] reg2016 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2013 = (1'h0);
  reg [(5'h16):(1'h0)] reg2010 = (1'h0);
  reg [(2'h3):(1'h0)] reg2007 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2004 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg425 = (1'h0);
  reg [(5'h10):(1'h0)] reg433 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar429 = (1'h0);
  reg [(3'h7):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg427 = (1'h0);
  reg [(4'hc):(1'h0)] forvar425 = (1'h0);
  reg [(3'h5):(1'h0)] reg424 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg422 = (1'h0);
  reg [(5'h12):(1'h0)] reg419 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar402 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg414 = (1'h0);
  reg [(4'hd):(1'h0)] reg411 = (1'h0);
  reg [(3'h5):(1'h0)] reg407 = (1'h0);
  reg signed [(4'he):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar398 = (1'h0);
  reg [(5'h18):(1'h0)] reg396 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg395 = (1'h0);
  reg [(2'h3):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg389 = (1'h0);
  reg [(5'h16):(1'h0)] reg387 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar386 = (1'h0);
  reg [(4'ha):(1'h0)] reg383 = (1'h0);
  reg [(5'h17):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg380 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg377 = (1'h0);
  reg [(4'hf):(1'h0)] reg376 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar375 = (1'h0);
  reg [(3'h7):(1'h0)] reg374 = (1'h0);
  reg [(4'he):(1'h0)] reg373 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg372 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg370 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg369 = (1'h0);
  reg [(3'h4):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar367 = (1'h0);
  reg [(4'hf):(1'h0)] reg366 = (1'h0);
  reg [(5'h1b):(1'h0)] reg365 = (1'h0);
  reg [(5'h11):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar361 = (1'h0);
  reg [(5'h10):(1'h0)] reg360 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg357 = (1'h0);
  reg [(5'h1b):(1'h0)] reg356 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar354 = (1'h0);
  reg [(5'h15):(1'h0)] reg352 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg350 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg349 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg347 = (1'h0);
  reg [(4'hd):(1'h0)] reg346 = (1'h0);
  reg [(3'h7):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg341 = (1'h0);
  reg [(5'h1c):(1'h0)] reg340 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg339 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg338 = (1'h0);
  reg signed [(4'he):(1'h0)] reg337 = (1'h0);
  reg [(5'h1c):(1'h0)] reg333 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg326 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar324 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar323 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar321 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg315 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg309 = (1'h0);
  reg [(4'h9):(1'h0)] reg308 = (1'h0);
  reg [(5'h1e):(1'h0)] reg306 = (1'h0);
  reg [(5'h16):(1'h0)] reg305 = (1'h0);
  reg [(5'h10):(1'h0)] reg298 = (1'h0);
  reg [(5'h1a):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg289 = (1'h0);
  reg [(4'hb):(1'h0)] reg286 = (1'h0);
  reg [(5'h1d):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar273 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg283 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar278 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg276 = (1'h0);
  reg [(5'h10):(1'h0)] reg275 = (1'h0);
  reg [(5'h10):(1'h0)] forvar272 = (1'h0);
  reg [(5'h1d):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg270 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg269 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg267 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg266 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar265 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg261 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg260 = (1'h0);
  reg [(5'h13):(1'h0)] forvar259 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg258 = (1'h0);
  reg [(4'hb):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg255 = (1'h0);
  reg [(4'hf):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar251 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg249 = (1'h0);
  reg [(5'h1b):(1'h0)] reg245 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg241 = (1'h0);
  reg [(5'h1d):(1'h0)] reg237 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg236 = (1'h0);
  reg [(5'h1c):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg233 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar230 = (1'h0);
  assign y = {wire2098,
                 wire2000,
                 wire1999,
                 wire1997,
                 wire319,
                 wire293,
                 wire292,
                 wire291,
                 wire229,
                 reg2100,
                 reg2116,
                 reg2115,
                 reg2114,
                 reg2112,
                 reg2111,
                 reg2108,
                 reg2107,
                 reg2106,
                 reg2104,
                 reg2102,
                 reg2101,
                 reg2096,
                 reg2093,
                 reg2089,
                 reg2085,
                 reg2084,
                 reg2083,
                 reg2065,
                 reg2082,
                 reg2080,
                 reg2079,
                 reg2078,
                 reg2076,
                 reg2074,
                 reg2072,
                 reg2071,
                 reg2067,
                 reg2066,
                 reg2064,
                 reg2063,
                 reg2062,
                 reg2060,
                 reg2058,
                 reg2056,
                 reg2054,
                 reg2049,
                 reg2046,
                 reg2045,
                 reg2044,
                 reg2042,
                 reg2041,
                 reg2039,
                 reg2036,
                 reg2035,
                 reg2031,
                 reg2029,
                 reg2024,
                 reg2022,
                 reg2020,
                 reg2017,
                 reg2015,
                 reg2014,
                 reg2012,
                 reg2011,
                 reg2009,
                 reg2008,
                 reg2006,
                 reg2005,
                 reg2003,
                 reg2002,
                 reg2001,
                 reg231,
                 reg232,
                 reg238,
                 reg239,
                 reg240,
                 reg242,
                 reg243,
                 reg246,
                 reg247,
                 reg248,
                 reg250,
                 reg252,
                 reg253,
                 reg257,
                 reg262,
                 reg264,
                 reg273,
                 reg274,
                 reg277,
                 reg279,
                 reg280,
                 reg281,
                 reg282,
                 reg284,
                 reg272,
                 reg278,
                 reg287,
                 reg288,
                 reg295,
                 reg296,
                 reg299,
                 reg300,
                 reg301,
                 reg302,
                 reg303,
                 reg304,
                 reg307,
                 reg311,
                 reg312,
                 reg314,
                 reg316,
                 reg317,
                 reg320,
                 reg325,
                 reg327,
                 reg328,
                 reg329,
                 reg330,
                 reg331,
                 reg332,
                 reg334,
                 reg335,
                 reg336,
                 reg342,
                 reg343,
                 reg345,
                 reg348,
                 reg351,
                 reg353,
                 reg355,
                 reg358,
                 reg362,
                 reg371,
                 reg378,
                 reg379,
                 reg381,
                 reg384,
                 reg385,
                 reg388,
                 reg390,
                 reg391,
                 reg392,
                 reg394,
                 reg397,
                 reg400,
                 reg401,
                 reg403,
                 reg404,
                 reg405,
                 reg406,
                 reg408,
                 reg409,
                 reg410,
                 reg412,
                 reg413,
                 reg415,
                 reg417,
                 reg420,
                 reg421,
                 reg423,
                 reg426,
                 reg430,
                 reg431,
                 reg432,
                 reg2117,
                 forvar2106,
                 reg2113,
                 reg2110,
                 reg2109,
                 reg2105,
                 reg2103,
                 forvar2100,
                 reg2099,
                 reg2097,
                 reg2095,
                 forvar2094,
                 reg2092,
                 reg2091,
                 reg2090,
                 reg2088,
                 reg2087,
                 forvar2086,
                 reg2081,
                 forvar2076,
                 reg2073,
                 forvar2064,
                 forvar2081,
                 reg2077,
                 reg2075,
                 forvar2073,
                 reg2070,
                 reg2069,
                 reg2068,
                 forvar2065,
                 reg2061,
                 reg2059,
                 reg2057,
                 reg2055,
                 reg2053,
                 reg2052,
                 reg2051,
                 reg2050,
                 reg2048,
                 reg2047,
                 reg2043,
                 reg2040,
                 reg2038,
                 reg2037,
                 reg2034,
                 reg2033,
                 reg2032,
                 forvar2030,
                 reg2028,
                 reg2027,
                 reg2026,
                 forvar2025,
                 reg2023,
                 reg2021,
                 reg2019,
                 reg2018,
                 reg2016,
                 reg2013,
                 reg2010,
                 reg2007,
                 reg2004,
                 reg425,
                 reg433,
                 forvar429,
                 reg428,
                 reg427,
                 forvar425,
                 reg424,
                 reg422,
                 reg419,
                 reg418,
                 forvar402,
                 reg398,
                 reg416,
                 reg414,
                 reg411,
                 reg407,
                 reg402,
                 reg399,
                 forvar398,
                 reg396,
                 reg395,
                 reg393,
                 reg389,
                 reg387,
                 forvar386,
                 reg383,
                 reg382,
                 reg380,
                 reg377,
                 reg376,
                 forvar375,
                 reg374,
                 reg373,
                 reg372,
                 reg370,
                 reg369,
                 reg368,
                 forvar367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 forvar361,
                 reg360,
                 reg359,
                 reg357,
                 reg356,
                 forvar354,
                 reg352,
                 reg350,
                 reg349,
                 reg347,
                 reg346,
                 reg344,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg333,
                 reg326,
                 forvar324,
                 forvar323,
                 reg322,
                 forvar321,
                 reg318,
                 reg315,
                 reg313,
                 reg310,
                 reg309,
                 reg308,
                 reg306,
                 reg305,
                 reg298,
                 reg297,
                 reg294,
                 reg290,
                 reg289,
                 reg286,
                 reg285,
                 forvar273,
                 reg283,
                 forvar278,
                 reg276,
                 reg275,
                 forvar272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 forvar265,
                 reg263,
                 reg261,
                 reg260,
                 forvar259,
                 reg258,
                 reg256,
                 reg255,
                 reg254,
                 forvar251,
                 reg249,
                 reg245,
                 reg244,
                 reg241,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 forvar230,
                 (1'h0)};
  assign wire229 = (^~$unsigned({(wire225 ?
                           $signed(wire228) : $unsigned(wire227))}));
  always
    @(posedge clk) begin
      for (forvar230 = (1'h0); (forvar230 < (2'h3)); forvar230 = (forvar230 + (1'h1)))
        begin
          if ((wire227[(1'h1):(1'h1)] ?
              $signed($unsigned({$unsigned(wire229),
                  $unsigned((8'ha9)),
                  $signed((8'ha5))})) : $signed(forvar230)))
            begin
              reg231 <= {(7'h51),
                  $unsigned(((|{wire228, wire228, wire226}) ?
                      (wire228 ? (^~wire228) : ((8'ha9) < wire225)) : wire225)),
                  (wire225[(3'h4):(2'h3)] != $signed($unsigned((wire225 - wire225))))};
              reg232 <= ((((!$unsigned(wire225)) ^ $unsigned(forvar230[(1'h0):(1'h0)])) & $signed(wire229)) || ((~&$unsigned((wire225 ?
                  wire227 : (8'h9d)))) >> (-($unsigned(forvar230) * (reg231 ?
                  wire226 : wire225)))));
              reg233 = $unsigned((($signed({wire226, wire226, wire227}) ?
                      wire226 : wire226) ?
                  $unsigned(wire228[(3'h7):(3'h5)]) : ($signed((wire226 + reg232)) ?
                      {$unsigned(wire227),
                          reg231[(1'h1):(1'h0)],
                          $unsigned(wire228)} : $signed($signed((8'hb4))))));
              reg234 = $signed(reg232);
              reg235 = $signed(((~&(&(~&wire228))) >>> (wire229[(1'h1):(1'h0)] ?
                  (|(wire228 ? (7'h50) : wire227)) : (|(wire229 >= wire225)))));
              reg236 = ((~&$signed(reg234)) - wire226);
              reg237 = {($unsigned((forvar230 ~^ $unsigned(wire225))) * (^~reg233)),
                  (7'h4e),
                  ($unsigned($signed((reg234 && wire229))) ?
                      (wire227[(3'h4):(1'h1)] ?
                          {((7'h52) ? wire229 : reg231)} : $signed({wire228,
                              reg235})) : wire226)};
            end
          else
            begin
              reg231 <= $signed(wire228);
              reg232 <= (($signed({{(7'h41)}, reg235, {wire228, reg234}}) ?
                      reg235[(4'hc):(3'h4)] : $signed(({(7'h44),
                          reg231,
                          reg231} - $signed(wire227)))) ?
                  ({{(~|reg237), $signed(wire228)}} ?
                      $unsigned(($unsigned(reg236) ^~ (^reg231))) : wire227) : wire229[(4'hd):(2'h2)]);
              reg233 = forvar230;
              reg234 = reg231;
              reg238 <= $unsigned(wire225);
              reg239 <= $signed(wire227);
              reg240 <= (!wire228[(3'h4):(1'h0)]);
            end
          if (reg231)
            begin
              reg241 = $signed(((($unsigned(reg239) ?
                  (reg231 * reg234) : (~wire225)) >> reg231) <= $unsigned(wire229)));
            end
          else
            begin
              reg242 <= $unsigned((({$signed(reg236),
                      (wire227 ? reg239 : (7'h4d))} >>> wire227) ?
                  reg231[(3'h4):(1'h1)] : ((wire225 <<< reg236[(4'h8):(3'h4)]) ?
                      (+$unsigned(wire228)) : $unsigned(reg241))));
              reg243 <= {({(wire225 ~^ (&reg232)),
                          (7'h43),
                          ($unsigned((8'hab)) >>> ((8'hac) ?
                              wire228 : reg238))} ?
                      (($signed(reg241) ? (reg237 * reg239) : (8'ha7)) ?
                          (+(wire229 ?
                              reg233 : reg232)) : $unsigned(wire229[(5'h15):(4'h9)])) : reg231),
                  (reg234[(4'h9):(4'h8)] ?
                      $unsigned((~|reg232)) : (reg232 ~^ (+(~^wire229)))),
                  (+$signed((+(reg233 << (8'ha6)))))};
              reg244 = $unsigned((!$unsigned($unsigned(reg234))));
              reg245 = (($unsigned({(^reg243),
                          $signed(wire225),
                          {(7'h55), (7'h43), reg243}}) ?
                      $signed(reg240) : (8'h9d)) ?
                  {(forvar230[(1'h1):(1'h0)] ?
                          (reg237[(3'h5):(3'h4)] || $signed(reg237)) : (reg232[(1'h1):(1'h0)] ?
                              wire229[(2'h2):(1'h1)] : (wire226 < reg241))),
                      $unsigned((reg243[(3'h4):(1'h0)] ?
                          (reg239 ~^ reg243) : (wire228 ? (8'hab) : reg235))),
                      $signed((-((7'h4a) == wire228)))} : wire228[(3'h4):(2'h2)]);
            end
          if (($unsigned($signed($unsigned(wire225[(4'hc):(3'h6)]))) ?
              forvar230 : $signed($unsigned((((7'h4a) ?
                  (8'hb2) : reg244) & $unsigned(reg235))))))
            begin
              reg246 <= $signed($unsigned(reg243[(5'h13):(4'he)]));
              reg247 <= (wire227 << (!reg235));
              reg248 <= reg245;
              reg249 = ((-$unsigned(reg233)) == (+wire228));
            end
          else
            begin
              reg246 <= forvar230;
              reg247 <= $signed(((^(^(-wire226))) ?
                  (&(^(reg246 != reg242))) : reg246[(4'hb):(4'hb)]));
              reg249 = wire227;
              reg250 <= $signed($signed((8'h9d)));
            end
          for (forvar251 = (1'h0); (forvar251 < (3'h6)); forvar251 = (forvar251 + (1'h1)))
            begin
              reg252 <= $signed((($unsigned($signed((7'h4a))) ?
                  (~&(|reg249)) : (7'h4a)) <= (|((reg236 == reg244) == reg243))));
              reg253 <= {$unsigned(($signed((~^reg237)) ?
                      (+reg240[(3'h5):(2'h3)]) : (+$unsigned(reg239)))),
                  ((+{(reg237 & reg233)}) ? reg243 : (+reg249[(1'h0):(1'h0)]))};
              reg254 = ((~^$unsigned($signed(reg244[(2'h2):(2'h2)]))) != $unsigned(reg252[(3'h5):(2'h3)]));
              reg255 = (~|(-{$unsigned((&reg236)),
                  ($signed(reg248) ? {reg252, reg246, reg248} : (~&(8'hbf))),
                  wire226}));
              reg256 = (8'ha1);
              reg257 <= ($unsigned(((8'ha9) >> ($unsigned(reg244) != $unsigned(reg252)))) - $signed($unsigned(reg241)));
              reg258 = $unsigned(reg247[(3'h5):(1'h0)]);
            end
          for (forvar259 = (1'h0); (forvar259 < (1'h0)); forvar259 = (forvar259 + (1'h1)))
            begin
              reg260 = (reg235 ? reg258 : reg240[(1'h0):(1'h0)]);
              reg261 = ((^(($unsigned(reg231) ~^ $unsigned(reg235)) < $unsigned($signed(reg244)))) >>> $unsigned(reg247[(5'h13):(3'h7)]));
            end
          reg262 <= (($signed($signed((~^forvar230))) <<< ($signed((reg246 ?
                  wire229 : reg233)) & $unsigned((reg241 << wire226)))) ?
              reg243 : $unsigned((~^($unsigned(reg260) ?
                  reg247[(5'h1e):(5'h10)] : $signed(reg237)))));
          reg263 = (|$unsigned(($signed($unsigned(reg232)) ?
              $unsigned((~&reg261)) : ($signed(reg250) > (reg260 ?
                  forvar251 : reg231)))));
        end
      reg264 <= (~^(wire228[(4'hc):(4'ha)] << $signed({wire227})));
      for (forvar265 = (1'h0); (forvar265 < (3'h5)); forvar265 = (forvar265 + (1'h1)))
        begin
          reg266 = forvar265[(4'h8):(4'h8)];
          reg267 = (!reg249);
          if (reg267)
            begin
              reg268 = (+$unsigned((~|((reg237 ^~ reg234) ?
                  (forvar251 ? wire226 : reg242) : ((7'h4d) >= reg250)))));
              reg269 = reg261;
              reg270 = reg261[(3'h4):(2'h3)];
            end
          else
            begin
              reg268 = reg254[(4'h8):(1'h0)];
            end
        end
      reg271 = $signed($signed(reg241));
      if ({(reg235 | $unsigned((|reg235[(5'h15):(3'h7)]))),
          $signed($signed(((~|(7'h41)) ? {reg268} : (reg268 && (8'hb3)))))})
        begin
          for (forvar272 = (1'h0); (forvar272 < (3'h4)); forvar272 = (forvar272 + (1'h1)))
            begin
              reg273 <= wire226[(4'hf):(3'h5)];
              reg274 <= $signed(forvar272[(1'h0):(1'h0)]);
              reg275 = $signed($unsigned({wire228}));
              reg276 = (((((reg237 ? reg249 : wire229) ?
                  {reg261,
                      reg241,
                      reg240} : $signed(reg256)) <= $unsigned((~reg231))) >> (!($unsigned((7'h4f)) - (reg260 && reg252)))) >> $signed((($unsigned(reg231) > (wire226 ?
                      wire225 : forvar251)) ?
                  $signed(reg254[(3'h6):(1'h0)]) : $signed(reg271))));
              reg277 <= reg271;
            end
          for (forvar278 = (1'h0); (forvar278 < (3'h6)); forvar278 = (forvar278 + (1'h1)))
            begin
              reg279 <= ({reg257[(4'hb):(4'ha)]} == (~&{reg277,
                  reg257[(4'ha):(3'h5)],
                  reg269[(3'h6):(2'h2)]}));
              reg280 <= $signed(wire228);
              reg281 <= wire226[(4'h9):(4'h8)];
              reg282 <= ((~|forvar230[(4'h8):(3'h5)]) ?
                  reg239 : {(reg236 ?
                          {reg239, reg281[(5'h1e):(5'h1b)]} : $signed(reg276)),
                      forvar259[(3'h4):(1'h0)]});
              reg283 = ($unsigned(((((7'h55) ~^ reg282) ?
                          reg238 : $signed(reg241)) ?
                      ($signed(reg240) < wire228[(3'h7):(2'h2)]) : ((reg255 ?
                          reg277 : reg279) ^~ (+reg240)))) ?
                  reg253 : (~^(+($unsigned(reg233) ?
                      (~&reg234) : $signed(reg240)))));
              reg284 <= $signed($unsigned($signed($signed({reg276}))));
            end
        end
      else
        begin
          reg272 <= (reg242[(2'h2):(1'h0)] ?
              (reg249[(4'he):(4'h8)] >> reg279) : $signed(reg245[(5'h18):(5'h12)]));
          for (forvar273 = (1'h0); (forvar273 < (1'h1)); forvar273 = (forvar273 + (1'h1)))
            begin
              reg274 <= ((~($signed((reg232 ? reg246 : wire227)) ^ (7'h4e))) ?
                  (8'hbb) : ((((reg249 ? reg271 : reg254) ?
                      (~&reg240) : $signed(reg254)) <<< (!reg236)) ^~ $unsigned(forvar278)));
              reg277 <= {reg241[(3'h5):(3'h5)]};
              reg278 <= ((+forvar278[(3'h5):(1'h0)]) << (($unsigned($unsigned(reg242)) ?
                  $signed($signed(reg248)) : ((reg257 ? reg255 : reg240) ?
                      (wire227 + reg236) : reg242)) || $signed((reg256[(3'h5):(3'h5)] <<< reg252))));
              reg283 = {$signed(reg237[(5'h1c):(2'h3)]), reg255[(3'h4):(2'h3)]};
              reg285 = (reg233 ?
                  $unsigned((&(~&(~^reg257)))) : ($signed(reg271) >> reg257[(3'h6):(2'h3)]));
              reg286 = $unsigned(($signed({$unsigned(reg231),
                      reg252,
                      (~&reg278)}) ?
                  ($signed((|reg278)) ?
                      $unsigned((7'h56)) : $unsigned((wire227 ?
                          reg237 : forvar259))) : (($signed(reg271) == $unsigned(reg281)) ?
                      reg247 : ((reg233 ?
                          (7'h40) : (7'h56)) >>> $signed((8'hac))))));
            end
          reg287 <= $signed($signed(reg254));
          reg288 <= reg246;
          reg289 = $signed($unsigned(((!(reg278 == wire227)) >> ($signed(reg278) | (reg278 ^~ reg254)))));
        end
      reg290 = reg278[(5'h13):(4'he)];
    end
  assign wire291 = reg238;
  assign wire292 = $unsigned($signed(reg279));
  assign wire293 = (wire227[(1'h0):(1'h0)] ?
                       (reg242[(3'h4):(1'h0)] ?
                           {(+(reg274 <<< reg272)),
                               (~^(^~reg284)),
                               reg277} : $unsigned({$unsigned(reg278),
                               reg240[(2'h3):(2'h3)]})) : ((|reg280[(4'hb):(2'h2)]) >> $signed((~$signed(reg257)))));
  always
    @(posedge clk) begin
      if (((((|reg252) ? reg242 : (reg248 ? (~wire293) : $signed((7'h4d)))) ?
              $unsigned((reg273[(2'h2):(1'h0)] ?
                  (~|reg239) : reg250[(3'h4):(3'h4)])) : ((((7'h41) >= (7'h44)) >= (reg232 != reg282)) * reg246[(1'h1):(1'h1)])) ?
          (wire292 ?
              (reg247[(4'he):(3'h7)] - ($unsigned(reg262) && (+reg231))) : {(|(reg288 <= reg273))}) : {(^(-((7'h51) ?
                  reg262 : wire229)))}))
        begin
          reg294 = (wire229 >> $unsigned(wire229[(3'h6):(1'h0)]));
          reg295 <= $signed((&$signed(($unsigned(reg279) || $unsigned((8'haa))))));
          reg296 <= $signed($signed({((wire225 <= reg239) | (reg242 ?
                  (7'h53) : (7'h55))),
              reg250}));
          reg297 = $signed(({(~$signed(wire229)),
                  (reg284 ^ wire228),
                  {(!(8'hbf)), (~|reg277)}} ?
              (($unsigned(wire227) ^~ $unsigned(wire229)) ^ (reg281 == (reg231 >> reg231))) : (reg252 ?
                  reg240 : (((7'h49) & reg231) ~^ (&reg295)))));
          if ($signed((|(~^$signed(reg257[(4'ha):(1'h0)])))))
            begin
              reg298 = $unsigned((~|(((reg240 > wire292) ^~ $unsigned(reg274)) ?
                  $signed((!reg274)) : {(~&reg297),
                      ((8'hbd) ? reg278 : reg262)})));
              reg299 <= ({(8'hb4)} ?
                  (-($unsigned((reg250 ?
                      reg253 : wire225)) & ($signed(wire227) - reg294[(4'hb):(4'h9)]))) : reg242[(1'h0):(1'h0)]);
              reg300 <= {reg232, reg282, reg247};
              reg301 <= ({$unsigned((reg299[(1'h1):(1'h0)] && $signed(reg247))),
                      reg274[(4'h9):(4'h8)],
                      (reg231 ?
                          $signed($signed(wire226)) : reg277[(4'h9):(4'h9)])} ?
                  (~|(reg294[(5'h19):(5'h16)] ^~ {$unsigned(reg298)})) : {$unsigned(($unsigned(reg297) ?
                          $signed(reg277) : (wire293 ? (8'hb0) : reg299))),
                      ((!$unsigned(reg284)) >> {{wire225}}),
                      $unsigned(reg246[(2'h3):(1'h1)])});
              reg302 <= (reg264 ~^ $unsigned((($signed(reg282) ?
                      reg242 : $unsigned(reg299)) ?
                  {$unsigned(reg264),
                      (wire225 ~^ reg247),
                      (reg301 >= reg284)} : ({reg257, wire292, reg273} ?
                      (reg264 != reg294) : $signed(reg252)))));
              reg303 <= $signed($signed($signed(((reg273 >> reg278) ?
                  reg282[(3'h6):(3'h6)] : $unsigned(reg242)))));
              reg304 <= $signed({reg246[(5'h13):(1'h0)],
                  wire225,
                  reg239[(3'h7):(3'h6)]});
            end
          else
            begin
              reg299 <= reg301[(4'hf):(3'h5)];
              reg305 = reg240;
              reg306 = (~^reg296[(1'h0):(1'h0)]);
              reg307 <= {$unsigned(($unsigned((wire291 ? reg250 : reg300)) ?
                      wire292 : reg240)),
                  $unsigned((~^$unsigned((7'h52)))),
                  reg281[(5'h1c):(3'h6)]};
              reg308 = (((^~(|(reg240 ? wire293 : (8'ha9)))) >>> (((8'had) ?
                      reg294 : $unsigned(reg306)) ?
                  $signed((wire293 != reg301)) : $unsigned({(8'hab)}))) > $signed(wire225));
              reg309 = (-(~&reg302[(3'h6):(3'h6)]));
              reg310 = $unsigned($signed((~|reg248[(4'hf):(4'hc)])));
            end
          reg311 <= wire226[(5'h15):(4'ha)];
        end
      else
        begin
          if ($signed(reg247[(5'h13):(5'h12)]))
            begin
              reg295 <= wire292;
              reg297 = $unsigned($unsigned(reg274[(1'h1):(1'h0)]));
              reg299 <= (wire225 * ((~(~&(reg301 ? wire292 : reg232))) ?
                  $signed($unsigned($unsigned(reg243))) : $signed($signed((8'hb7)))));
            end
          else
            begin
              reg295 <= reg277;
              reg296 <= (($signed((((8'h9e) || reg301) ?
                      reg257[(1'h0):(1'h0)] : reg250)) ?
                  {(((7'h4c) ~^ reg288) ^ reg305)} : (({reg248} || ((7'h51) ?
                      reg243 : (8'h9c))) && $unsigned((reg311 ?
                      (8'ha9) : reg280)))) && {wire228[(2'h2):(2'h2)], reg279});
              reg297 = {{{{$signed(reg272)}}, reg274},
                  $unsigned(reg242[(2'h3):(1'h1)]),
                  reg302[(3'h7):(2'h2)]};
              reg299 <= $signed(reg309[(2'h2):(1'h0)]);
              reg300 <= $signed(wire229);
              reg301 <= reg288[(4'hf):(3'h7)];
              reg302 <= $signed(($signed(reg250[(3'h4):(1'h0)]) ?
                  reg287 : (reg294 || $signed((wire292 - reg299)))));
            end
          reg303 <= ((&reg248) ?
              ($signed($signed((~&wire228))) ?
                  (+(~|(reg281 >>> reg294))) : reg300[(2'h2):(2'h2)]) : reg264);
          reg305 = ($unsigned($unsigned(((reg311 ? reg303 : reg296) ?
                  (reg295 || reg232) : reg281))) ?
              {$signed(reg298),
                  ((^reg287) >>> reg311[(2'h3):(2'h3)])} : (~^((reg298[(4'he):(3'h4)] != $unsigned(reg274)) ?
                  reg253[(4'h9):(1'h1)] : ($unsigned(wire226) ^ reg287))));
          reg307 <= ((reg274 > (7'h43)) ?
              (-(reg299[(1'h0):(1'h0)] - $signed(reg302))) : reg296);
          if ({(reg239 ^~ reg303[(5'h17):(3'h7)])})
            begin
              reg311 <= (|($unsigned(({reg299} ?
                      reg299[(2'h2):(1'h1)] : ((8'ha4) ? wire293 : reg246))) ?
                  $unsigned((~(reg273 > wire229))) : (&((reg239 & reg277) ?
                      ((7'h4a) ? (7'h41) : reg300) : (wire228 ?
                          reg310 : reg253)))));
              reg312 <= $unsigned(reg239[(3'h7):(3'h5)]);
              reg313 = ((~|((reg278 ? reg250 : (^~(8'ha5))) ?
                  $unsigned((reg277 ?
                      reg287 : reg277)) : reg296[(3'h4):(3'h4)])) < reg264);
              reg314 <= ((~^$signed((~reg308[(3'h4):(1'h0)]))) + (reg247 & $signed(reg295)));
              reg315 = $unsigned((~&reg280[(2'h3):(2'h3)]));
              reg316 <= ((^((^$unsigned(reg288)) ?
                  ((&(8'ha3)) ?
                      {reg238,
                          wire293} : reg253) : ((reg303 ^ (8'hb1)) == $unsigned((8'ha8))))) ^ ($unsigned(((reg277 || reg307) * {reg247})) ?
                  $signed(((&reg297) >= reg312[(3'h7):(3'h5)])) : ($unsigned((+reg253)) ?
                      $unsigned(((7'h42) > reg284)) : ((reg312 ?
                          reg257 : reg309) == (~|(8'ha8))))));
              reg317 <= $unsigned(($unsigned(((~|reg248) < reg302)) ?
                  reg303[(2'h3):(2'h2)] : reg281));
            end
          else
            begin
              reg311 <= ((~^(8'haa)) ^~ $signed(({$signed(reg242)} ?
                  reg302 : $signed((^reg281)))));
              reg312 <= $signed(($signed(($unsigned(reg287) + (reg232 ?
                      reg274 : (8'ha6)))) ?
                  ((+((7'h43) >= reg240)) < ($unsigned(reg274) ?
                      reg305 : $unsigned(reg310))) : wire229));
            end
          reg318 = (&$signed({((wire293 != reg294) ^~ reg312[(3'h5):(2'h3)])}));
        end
    end
  assign wire319 = ($unsigned(($unsigned((reg304 ? (8'hb6) : reg231)) ?
                           $signed((reg301 ^ reg231)) : ({reg238, reg250} ?
                               $unsigned(reg279) : $signed(wire291)))) ?
                       $signed($signed(reg300)) : wire225);
  always
    @(posedge clk) begin
      reg320 <= reg279[(1'h0):(1'h0)];
      for (forvar321 = (1'h0); (forvar321 < (3'h6)); forvar321 = (forvar321 + (1'h1)))
        begin
          reg322 = $signed(wire319);
        end
      for (forvar323 = (1'h0); (forvar323 < (1'h0)); forvar323 = (forvar323 + (1'h1)))
        begin
          for (forvar324 = (1'h0); (forvar324 < (3'h5)); forvar324 = (forvar324 + (1'h1)))
            begin
              reg325 <= ((~$unsigned(reg278)) | (7'h4c));
              reg326 = reg320;
              reg327 <= ($unsigned((reg282[(3'h4):(2'h3)] ?
                  {reg301[(3'h5):(3'h5)]} : {(wire226 * reg246)})) | $signed((-(&(reg253 | reg303)))));
              reg328 <= reg262;
              reg329 <= reg303[(4'he):(2'h3)];
              reg330 <= ({(7'h58), reg264} ?
                  $signed($unsigned($signed((^reg317)))) : $unsigned({((reg238 <<< (8'h9e)) ?
                          $signed(wire292) : ((8'hb7) || reg316)),
                      reg304[(1'h1):(1'h1)],
                      reg242[(3'h4):(2'h2)]}));
            end
          if ((+reg281[(5'h17):(4'ha)]))
            begin
              reg331 <= (8'hb2);
              reg332 <= {reg327};
              reg333 = reg322;
              reg334 <= reg231[(2'h3):(2'h2)];
              reg335 <= reg257;
              reg336 <= (~&(8'hb4));
            end
          else
            begin
              reg333 = reg320;
              reg334 <= $signed({reg240[(2'h2):(1'h1)],
                  (reg311[(1'h1):(1'h1)] ?
                      (!reg242) : ((wire228 >= (8'h9e)) ? reg300 : reg316))});
              reg335 <= wire226[(4'he):(4'h9)];
              reg336 <= (reg316 ?
                  (^(($unsigned((8'haa)) ?
                          (reg272 != reg329) : wire229[(4'ha):(4'h8)]) ?
                      $signed((reg320 + reg334)) : reg333[(5'h1c):(3'h4)])) : {$signed($signed($unsigned(forvar323)))});
              reg337 = reg301;
            end
          if (((($unsigned((reg287 < reg311)) ?
                  ((reg325 == reg326) ?
                      (reg304 ?
                          reg280 : reg247) : (forvar324 & reg296)) : ($unsigned(reg334) | forvar321)) ?
              ($signed(reg300[(3'h5):(1'h1)]) ?
                  reg303 : {(reg240 ? reg328 : reg273),
                      $unsigned(reg302),
                      reg333[(5'h11):(4'h9)]}) : reg250) >>> ({$signed((reg282 > wire291))} ?
              ((reg330[(2'h3):(2'h2)] ?
                  $signed(reg242) : reg329) - (&reg246)) : reg264[(2'h2):(2'h2)])))
            begin
              reg338 = ($signed(reg278) ?
                  reg239[(4'hb):(1'h1)] : reg331[(4'hd):(4'h8)]);
              reg339 = reg239[(4'h8):(3'h7)];
              reg340 = reg243;
              reg341 = (($signed($signed(reg252)) != reg239[(3'h6):(2'h3)]) ?
                  $signed({(reg262[(3'h4):(2'h3)] >>> (&reg240)),
                      reg329[(5'h18):(3'h7)]}) : (+(!$signed($unsigned(reg332)))));
            end
          else
            begin
              reg338 = $unsigned($signed($unsigned(reg327[(5'h10):(3'h7)])));
              reg342 <= ((($signed($signed(reg303)) * (^(~^reg231))) ?
                  $unsigned(wire319) : $signed($signed($signed(forvar321)))) <<< ((((reg288 ?
                      reg312 : reg240) ?
                  $unsigned(reg338) : (reg303 ?
                      reg243 : reg279)) + (|$unsigned(reg282))) ~^ (reg247 ?
                  ($unsigned(reg246) ?
                      {(7'h50),
                          reg252,
                          (8'hba)} : reg326) : $unsigned($unsigned((8'hb8))))));
              reg343 <= (reg304 ?
                  $signed($unsigned(({reg331,
                      reg317} >>> (!wire293)))) : reg242[(3'h7):(2'h3)]);
              reg344 = $signed(forvar323[(1'h0):(1'h0)]);
              reg345 <= {$signed((7'h56)), reg240, reg329[(4'ha):(2'h3)]};
              reg346 = reg337;
            end
          reg347 = wire225[(3'h6):(2'h2)];
          if (reg240)
            begin
              reg348 <= (({(reg250[(3'h4):(2'h2)] ?
                          reg329 : {reg300, reg238, reg304}),
                      $unsigned((~|(7'h55))),
                      (-$unsigned(reg280))} ?
                  reg337[(4'h8):(3'h6)] : wire225[(2'h2):(2'h2)]) ~^ ((reg307[(2'h3):(1'h1)] ?
                  reg326 : reg332[(5'h13):(1'h0)]) == reg341));
              reg349 = {{{$unsigned({reg250, reg243, reg247}),
                          reg239[(2'h2):(1'h0)]},
                      $unsigned($signed(reg329[(5'h18):(5'h15)])),
                      reg346[(2'h2):(2'h2)]},
                  (7'h47)};
              reg350 = ($unsigned(reg330[(3'h7):(1'h0)]) * (8'h9c));
              reg351 <= (reg349[(1'h1):(1'h0)] ?
                  $signed((8'hac)) : {(reg231[(3'h5):(3'h5)] ?
                          (~^{wire226, reg288, reg327}) : reg281)});
              reg352 = $signed($signed($unsigned($unsigned($signed(reg351)))));
              reg353 <= ($signed((reg281 * (reg335 ?
                      reg287 : (reg351 >> (7'h53))))) ?
                  reg340[(5'h19):(5'h12)] : reg328);
            end
          else
            begin
              reg349 = wire225;
              reg350 = (|(&wire228));
            end
          for (forvar354 = (1'h0); (forvar354 < (3'h6)); forvar354 = (forvar354 + (1'h1)))
            begin
              reg355 <= reg322[(5'h13):(1'h1)];
              reg356 = ({((~^$unsigned((7'h46))) > reg296[(4'he):(2'h3)])} ?
                  $signed((reg329 == ((~reg349) || (reg287 != (8'ha9))))) : $unsigned($unsigned(reg336[(5'h1a):(4'hd)])));
              reg357 = $signed((~|(|((-reg257) ?
                  (reg345 ? reg345 : wire225) : $signed((7'h56))))));
              reg358 <= {reg242, $unsigned(wire291[(1'h1):(1'h1)]), reg350};
              reg359 = (wire227 ? wire293 : $signed({reg343[(5'h19):(2'h3)]}));
              reg360 = (reg320[(4'hb):(4'h9)] != {wire228,
                  (8'ha7),
                  $signed(reg274[(2'h3):(1'h1)])});
            end
        end
      for (forvar361 = (1'h0); (forvar361 < (1'h1)); forvar361 = (forvar361 + (1'h1)))
        begin
          if ($unsigned(reg335[(3'h4):(1'h1)]))
            begin
              reg362 <= (reg339[(3'h5):(1'h1)] ?
                  ($unsigned({$unsigned((7'h48)), $signed(reg280)}) ?
                      (($unsigned(reg316) ? reg349[(2'h2):(1'h0)] : reg358) ?
                          (reg345[(3'h6):(3'h6)] ?
                              (~|reg231) : $unsigned(reg355)) : $signed($unsigned(reg316))) : (((~reg284) ?
                          (reg348 < forvar324) : $unsigned((8'h9e))) << (!$unsigned(wire293)))) : $unsigned(reg231[(3'h7):(3'h5)]));
              reg363 = (reg355 ? $signed(reg296[(4'h8):(3'h7)]) : reg278);
              reg364 = reg358[(4'h8):(1'h1)];
              reg365 = ($signed($unsigned({$unsigned(reg311),
                  (~&reg301),
                  (wire229 ? (7'h4a) : reg248)})) * (~^reg343));
              reg366 = ((^~($unsigned(wire227[(1'h0):(1'h0)]) ?
                  wire293[(1'h1):(1'h1)] : $unsigned((+reg238)))) && {$unsigned($signed(reg331[(4'h9):(3'h5)]))});
            end
          else
            begin
              reg363 = {{$unsigned(((reg316 & reg238) ?
                          $signed((7'h43)) : (forvar361 > reg239))),
                      $signed($unsigned($unsigned((8'hb6)))),
                      $signed((^(~&reg366)))},
                  (~|$unsigned((reg334 ?
                      $unsigned(reg262) : {reg304, reg364})))};
            end
        end
      if ((~reg300))
        begin
          for (forvar367 = (1'h0); (forvar367 < (1'h1)); forvar367 = (forvar367 + (1'h1)))
            begin
              reg368 = (reg246 ?
                  $signed(reg287[(2'h2):(1'h1)]) : $signed(($unsigned($unsigned((7'h49))) ^ {(reg336 ?
                          reg362 : reg253),
                      (~&reg348),
                      (~|reg366)})));
              reg369 = $unsigned({(~(&(reg349 ? reg357 : (8'ha3)))),
                  ((-(wire319 ? reg322 : reg333)) ?
                      ((-reg272) & reg350) : {{wire292, reg277, reg231},
                          (~&forvar354)})});
              reg370 = reg295;
              reg371 <= $unsigned(reg231);
            end
          reg372 = reg347;
          reg373 = reg253;
        end
      else
        begin
          for (forvar367 = (1'h0); (forvar367 < (2'h3)); forvar367 = (forvar367 + (1'h1)))
            begin
              reg371 <= (((-($unsigned(reg329) || reg358[(1'h0):(1'h0)])) >= reg356[(3'h7):(2'h2)]) ?
                  {reg344[(1'h0):(1'h0)],
                      (reg350[(3'h7):(3'h5)] ?
                          (((7'h58) >= wire229) ?
                              {reg340,
                                  reg342} : (^reg348)) : ((&reg371) ^ (~&reg332))),
                      ((^(&reg303)) <<< $unsigned((reg274 & wire228)))} : forvar354);
            end
          reg372 = {reg317[(3'h4):(2'h2)]};
          reg373 = (&$unsigned((8'hb2)));
          reg374 = (-(wire291 ? (7'h48) : (~(~^reg364[(3'h4):(1'h0)]))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar375 = (1'h0); (forvar375 < (1'h1)); forvar375 = (forvar375 + (1'h1)))
        begin
          reg376 = {($unsigned((+$unsigned(reg327))) > reg320),
              (7'h4f),
              wire292};
          if ($signed(reg330[(5'h1f):(3'h4)]))
            begin
              reg377 = $signed((((((7'h47) ?
                      wire228 : wire292) ^~ (wire226 ^~ reg362)) ?
                  $unsigned(reg316[(5'h1b):(5'h1b)]) : ((reg248 ?
                          reg284 : reg307) ?
                      $signed(reg248) : $signed(reg274))) << reg353));
              reg378 <= (~^((8'hb4) ?
                  (~(^~(~reg250))) : reg246[(5'h1c):(4'hf)]));
              reg379 <= reg312[(3'h5):(1'h0)];
            end
          else
            begin
              reg378 <= ((|(({reg248} ~^ $signed(reg332)) ?
                      ((&reg334) <<< $signed(reg371)) : ($unsigned(reg253) ?
                          (reg273 >> reg300) : (&reg327)))) ?
                  $signed({(~^(reg329 ? reg296 : reg316)),
                      $unsigned(wire226)}) : (reg379[(4'hf):(2'h3)] ~^ {reg242}));
              reg380 = (!(^reg301));
              reg381 <= (((-(reg231 & reg274[(4'ha):(2'h2)])) - wire319[(2'h2):(2'h2)]) <= (~^($unsigned((reg232 != reg302)) ?
                  (reg278 ? reg311 : {reg296}) : (-(^~(7'h47))))));
              reg382 = $signed(reg287[(3'h5):(3'h5)]);
              reg383 = $signed(reg331[(4'h9):(2'h3)]);
              reg384 <= reg345;
            end
          reg385 <= (((reg288 ? $signed(reg325[(3'h7):(3'h6)]) : reg335) ?
              (((reg250 ?
                  reg231 : reg343) == reg329[(5'h14):(4'hd)]) ~^ wire229) : (-$signed((reg282 ?
                  reg273 : reg288)))) ^ (((8'h9c) | reg331) && reg362[(5'h16):(3'h4)]));
          for (forvar386 = (1'h0); (forvar386 < (3'h6)); forvar386 = (forvar386 + (1'h1)))
            begin
              reg387 = {(~&(reg311 ?
                      $signed((!reg320)) : (forvar386[(1'h0):(1'h0)] ?
                          (~|wire227) : (reg239 & reg303)))),
                  $unsigned($unsigned({{reg247, reg376},
                      $signed(reg280),
                      {wire227}}))};
              reg388 <= reg381[(4'he):(4'hd)];
              reg389 = wire229[(3'h4):(1'h1)];
              reg390 <= reg304;
              reg391 <= {reg296,
                  ($signed((~^$signed((8'hb3)))) ?
                      reg327[(3'h6):(3'h6)] : {$unsigned((~^reg320))})};
              reg392 <= {reg355[(4'hd):(3'h4)],
                  (|(reg382[(5'h12):(4'h8)] ?
                      $unsigned($signed(wire229)) : reg257)),
                  (|{$unsigned(((7'h56) ? reg331 : reg302)),
                      reg383[(4'h8):(2'h3)]})};
            end
          reg393 = {(({(reg301 ? forvar375 : reg388),
                      wire225,
                      {reg329}} != $unsigned((forvar386 != reg273))) ?
                  ($signed((!(8'h9e))) ?
                      ((reg314 >> reg300) ?
                          (&wire226) : $unsigned(reg392)) : $unsigned((!reg355))) : (&$signed($signed(reg238)))),
              wire227[(4'h9):(3'h5)]};
          reg394 <= $signed((reg278[(5'h15):(3'h7)] ^ (|reg343)));
        end
      reg395 = ((reg385 == $unsigned(reg362[(3'h6):(3'h6)])) ?
          ($unsigned($unsigned(reg240[(1'h1):(1'h1)])) <= reg282) : reg378);
      reg396 = (~&(8'h9e));
      if (((~|((reg246[(4'h8):(3'h5)] ?
          (!reg336) : reg379[(4'hc):(2'h2)]) <<< (&(&wire226)))) <= ((^((^~reg384) > ((7'h52) ~^ reg240))) ?
          (reg343[(4'hd):(4'hb)] ?
              reg242 : (!reg325[(4'h9):(3'h6)])) : reg351)))
        begin
          reg397 <= $signed(($signed($signed((~(8'hb2)))) ?
              $unsigned($signed((reg380 ?
                  reg396 : reg351))) : (($unsigned((7'h55)) ?
                  $unsigned(reg383) : (~|wire225)) ^~ $signed((!reg331)))));
          for (forvar398 = (1'h0); (forvar398 < (1'h1)); forvar398 = (forvar398 + (1'h1)))
            begin
              reg399 = ($unsigned({((reg247 * reg384) ^ (7'h50)),
                      {reg307},
                      reg257[(3'h5):(3'h4)]}) ?
                  $unsigned(($signed(reg377) && (~&(reg320 ?
                      reg277 : reg389)))) : (reg378[(1'h0):(1'h0)] ?
                      forvar398[(3'h6):(2'h2)] : (reg316[(5'h16):(4'hd)] ?
                          (^~reg231[(3'h5):(2'h2)]) : ((!reg262) ?
                              (^~forvar398) : (reg336 ? reg329 : reg281)))));
              reg400 <= $unsigned(reg282[(3'h7):(2'h2)]);
              reg401 <= ($unsigned((({reg325, reg239, reg253} * (~reg325)) ?
                  $unsigned($unsigned(wire292)) : (~|reg376))) >= ($signed($unsigned((~^reg351))) ?
                  (^~reg394[(4'hf):(3'h6)]) : reg383[(3'h4):(2'h2)]));
              reg402 = (((8'h9c) * reg299) < (7'h44));
              reg403 <= reg384[(1'h1):(1'h0)];
              reg404 <= (((|((7'h40) ?
                      {(8'ha3),
                          (7'h57),
                          (8'hb7)} : (~^forvar398))) != (reg358[(2'h2):(1'h0)] ?
                      {$signed(reg400)} : $unsigned(reg280[(4'hb):(2'h3)]))) ?
                  reg389[(4'hf):(1'h0)] : $unsigned({reg232,
                      $signed({reg272, reg376})}));
              reg405 <= ((($signed({reg381, reg343, (8'ha0)}) ?
                          $unsigned((reg232 <= reg399)) : {$unsigned(reg380)}) ?
                      (($unsigned(reg252) ?
                              (+(7'h44)) : reg395[(3'h4):(3'h4)]) ?
                          $unsigned((reg402 ?
                              (7'h4d) : forvar375)) : $unsigned($unsigned(reg379))) : $signed((reg312 ?
                          reg343[(5'h16):(5'h15)] : ((7'h56) >= reg257)))) ?
                  $unsigned($unsigned($signed((reg264 <<< reg362)))) : (^$signed((8'hbb))));
            end
          reg406 <= $unsigned(((!(((8'hb4) ? reg262 : reg299) ?
              reg335[(1'h1):(1'h1)] : $signed((8'haa)))) >>> (($unsigned(reg401) ?
                  (&reg358) : ((7'h41) << reg329)) ?
              ((~&reg288) || (reg345 <<< reg257)) : $unsigned(reg264[(2'h3):(1'h1)]))));
          reg407 = reg383;
          if ($signed({(reg317[(3'h5):(2'h3)] ^~ ($signed(reg401) != reg392)),
              $signed($unsigned($unsigned(reg314))),
              $signed(reg250)}))
            begin
              reg408 <= $unsigned(reg395);
              reg409 <= reg334[(1'h0):(1'h0)];
              reg410 <= $unsigned(reg332);
              reg411 = {$signed(reg348),
                  $signed($unsigned({$signed(reg377),
                      (reg257 & reg330),
                      (reg343 ? wire292 : reg278)})),
                  reg336[(4'he):(4'h8)]};
              reg412 <= reg253;
              reg413 <= (~|$signed($unsigned({wire228[(3'h6):(2'h2)],
                  $unsigned(reg411),
                  $unsigned(reg382)})));
              reg414 = (reg381 - (7'h51));
            end
          else
            begin
              reg411 = reg401[(2'h3):(1'h1)];
              reg412 <= $signed(reg303);
              reg413 <= (8'haf);
              reg414 = (($signed(reg376) + (~&((wire227 ? reg302 : reg311) ?
                      reg316 : (~|reg264)))) ?
                  reg288 : (reg396[(5'h15):(1'h0)] ?
                      reg317[(3'h6):(2'h3)] : $signed($unsigned((reg279 ?
                          (8'ha0) : reg240)))));
              reg415 <= {(~((+reg301) ^ ($unsigned(reg376) <= reg320[(4'hb):(4'h8)])))};
              reg416 = (|$signed((!(8'h9e))));
              reg417 <= wire225;
            end
        end
      else
        begin
          if (reg314)
            begin
              reg397 <= $signed(reg389[(4'h8):(3'h6)]);
            end
          else
            begin
              reg397 <= reg274;
              reg398 = {$signed($signed((7'h52))),
                  {$unsigned($unsigned(reg257)),
                      reg288[(5'h12):(4'ha)],
                      reg351}};
              reg400 <= reg403;
            end
          reg401 <= $unsigned((reg303[(5'h16):(1'h0)] ^ $unsigned(reg325[(3'h5):(3'h4)])));
          for (forvar402 = (1'h0); (forvar402 < (1'h1)); forvar402 = (forvar402 + (1'h1)))
            begin
              reg407 = ($signed((+$unsigned(reg395))) ^ $unsigned((((reg343 == reg325) <<< reg343) >= {(reg334 > reg342),
                  (-wire225)})));
              reg408 <= $unsigned($unsigned(($unsigned((reg332 ?
                      reg404 : wire226)) ?
                  $unsigned((reg279 > reg330)) : $signed((reg381 > reg397)))));
              reg411 = $unsigned($signed((+$signed(reg279[(4'hb):(4'hb)]))));
              reg412 <= (~|$unsigned(($unsigned($signed(reg383)) ?
                  reg405 : $unsigned($unsigned(reg296)))));
              reg414 = $unsigned({$signed(($signed(reg246) ?
                      {reg399, reg382, reg327} : (+wire319))),
                  ($unsigned((^~(8'ha1))) + reg405)});
            end
          if (reg417[(4'h9):(3'h4)])
            begin
              reg416 = ((8'hbc) ~^ reg320);
            end
          else
            begin
              reg416 = (reg395[(3'h4):(3'h4)] ?
                  $signed((~&$signed((~|reg231)))) : (((^~reg407) ?
                          reg317 : $unsigned(reg299)) ?
                      reg414[(3'h5):(2'h2)] : (~|((^reg274) || (reg355 ?
                          reg396 : (8'ha4))))));
              reg418 = (&reg331);
              reg419 = $unsigned(wire227);
              reg420 <= ((~|$signed((~|(reg405 ?
                  (7'h55) : reg302)))) < (~|(8'hb7)));
            end
          reg421 <= {$signed(($signed({(7'h4e), forvar386}) ?
                  reg331 : (wire293[(2'h2):(2'h2)] < wire319[(1'h0):(1'h0)]))),
              (($unsigned(reg328[(4'hd):(3'h5)]) & ($signed(wire292) ~^ (8'hb3))) ?
                  (~^$signed($signed(reg316))) : (wire229[(3'h6):(3'h5)] <= $unsigned($signed((7'h45)))))};
          reg422 = reg414;
        end
      reg423 <= $signed({($unsigned((reg351 != reg247)) <<< $unsigned((reg311 ?
              reg328 : (8'hb3)))),
          (-forvar386[(3'h4):(2'h3)])});
      reg424 = reg316[(4'he):(1'h1)];
      if ($signed($signed(reg287)))
        begin
          for (forvar425 = (1'h0); (forvar425 < (2'h3)); forvar425 = (forvar425 + (1'h1)))
            begin
              reg426 <= $unsigned($unsigned(wire228));
              reg427 = {$unsigned((^$unsigned($unsigned((7'h58))))),
                  $unsigned(reg332[(2'h3):(1'h0)]),
                  reg400};
              reg428 = (8'hb5);
            end
          for (forvar429 = (1'h0); (forvar429 < (3'h6)); forvar429 = (forvar429 + (1'h1)))
            begin
              reg430 <= (reg325[(3'h6):(1'h0)] || $signed(($unsigned((reg232 != reg393)) ?
                  reg278 : reg394)));
            end
          reg431 <= (reg273 ?
              ({((reg400 ^~ (8'hb8)) ?
                          (reg240 ? reg342 : reg393) : (reg388 ?
                              reg231 : (8'hac)))} ?
                  ({$unsigned(reg273),
                      $signed(wire293),
                      (~reg277)} | ({forvar429} ?
                      (7'h42) : reg335)) : (~|((-reg424) == (~^reg428)))) : (((~(reg430 * reg240)) > reg362) << reg396[(5'h18):(5'h14)]));
          reg432 <= ({((~&$unsigned(reg240)) == $signed((reg430 ?
                  (8'ha8) : forvar425))),
              $signed($signed(reg243[(4'hc):(4'h8)])),
              (reg274[(4'hb):(1'h0)] && $signed({(8'ha3), reg281}))} < reg288);
          reg433 = $signed($signed(reg262[(4'h8):(1'h1)]));
        end
      else
        begin
          reg425 = reg311;
        end
    end
  module434 #() modinst1998 (wire1997, clk, reg253, reg328, reg336, reg362, reg307);
  assign wire1999 = reg279;
  assign wire2000 = reg288;
  always
    @(posedge clk) begin
      if (wire227[(1'h0):(1'h0)])
        begin
          reg2001 <= (({$unsigned(reg379)} ?
              wire226[(4'hf):(1'h0)] : {{(~&reg404)}}) < ($signed($unsigned((reg426 ?
              reg277 : reg409))) << $signed($unsigned(reg401))));
          reg2002 <= (($unsigned(wire229[(4'ha):(3'h7)]) ?
              reg430[(3'h4):(1'h0)] : ($signed($signed(reg327)) ?
                  ((reg232 ? (8'haa) : reg327) ?
                      $unsigned(wire227) : $signed((8'ha9))) : {{(8'hba)},
                      (wire2000 ?
                          (8'hb7) : reg273)})) > reg262[(5'h1e):(5'h1b)]);
          if ($signed($signed($unsigned((7'h49)))))
            begin
              reg2003 <= (!$signed(((-reg281[(2'h3):(1'h1)]) <= $signed((reg336 >>> reg317)))));
              reg2004 = ($unsigned(reg248) ?
                  ({(((7'h53) >>> reg278) ? reg348 : reg384),
                          ($unsigned(reg250) * ((8'h9c) >= reg353)),
                          (reg295 == (reg378 ? reg392 : reg238))} ?
                      (!$signed((reg336 ?
                          reg423 : reg280))) : (8'h9d)) : reg330[(4'hb):(2'h3)]);
              reg2005 <= (8'hba);
              reg2006 <= (reg345[(3'h6):(3'h6)] && {({(~|reg392),
                          $signed(reg239)} ?
                      reg330 : reg328),
                  wire1999});
              reg2007 = reg355[(4'h8):(3'h4)];
              reg2008 <= $unsigned(($signed((|{reg296, (8'ha6)})) ?
                  ((^~(~|reg287)) | {(-reg2003)}) : $signed(($unsigned(reg410) < reg246[(4'hc):(2'h2)]))));
              reg2009 <= $signed($signed($signed(((-wire1997) - reg246[(2'h2):(2'h2)]))));
            end
          else
            begin
              reg2004 = {$unsigned(reg329),
                  $signed($signed((reg426[(2'h3):(1'h1)] ?
                      (reg379 & (7'h46)) : reg262[(5'h13):(4'hb)]))),
                  $unsigned({((~&reg362) ? reg238[(3'h5):(1'h0)] : (~|reg320)),
                      $signed(reg385),
                      (|(~&reg406))})};
              reg2007 = reg2008[(2'h3):(1'h0)];
              reg2008 <= {$signed({$unsigned((reg431 < (8'hbf))),
                      $unsigned((reg404 ? reg317 : reg353)),
                      $unsigned(reg242)}),
                  reg329,
                  ({$signed((reg351 ? reg281 : reg401)),
                          (&reg278),
                          ($signed(reg417) >>> reg336[(1'h1):(1'h0)])} ?
                      reg345 : reg390[(3'h6):(3'h4)])};
              reg2009 <= {(&($unsigned($unsigned(reg336)) < $signed((reg2004 ^~ reg262))))};
              reg2010 = ((-reg302[(1'h0):(1'h0)]) ?
                  (|($signed(reg264[(1'h0):(1'h0)]) < reg371[(3'h6):(3'h6)])) : ((8'ha4) ?
                      ((reg371 ?
                          (^reg351) : (reg299 < reg2006)) <<< reg385) : (((^reg358) ?
                          $signed(reg410) : (reg334 <= reg242)) != reg300)));
              reg2011 <= $unsigned(wire319);
              reg2012 <= (~|$signed((&$signed(wire2000))));
            end
        end
      else
        begin
          reg2004 = reg253;
          reg2005 <= (reg2002[(2'h3):(1'h0)] ?
              (($unsigned($unsigned((8'ha0))) ^~ (reg379 ?
                  (7'h40) : (+wire225))) | reg351[(5'h13):(2'h2)]) : ($unsigned(reg2012[(4'hd):(3'h6)]) & $signed(($signed(wire1999) ?
                  (reg2007 ? reg342 : (8'ha6)) : $unsigned(reg332)))));
          if (reg302)
            begin
              reg2006 <= reg307;
              reg2008 <= (8'hb4);
              reg2009 <= (-(^((~&(-reg394)) ?
                  ((wire292 ? reg371 : reg390) ?
                      $unsigned(wire292) : $signed(reg358)) : (^$unsigned((7'h45))))));
              reg2011 <= $unsigned((!(|((reg272 ?
                  reg303 : reg378) < $unsigned(reg401)))));
            end
          else
            begin
              reg2007 = {$signed({reg381[(4'he):(4'h8)],
                      reg317[(3'h7):(3'h5)]}),
                  ((!reg312) ? reg400[(4'ha):(2'h3)] : reg250),
                  (~|reg2009[(3'h5):(1'h0)])};
              reg2008 <= $unsigned({(8'ha7),
                  (reg281 > {(reg238 ? reg242 : wire227)})});
              reg2009 <= ((reg385[(4'h8):(4'h8)] ?
                  reg384[(5'h11):(2'h2)] : reg2002[(5'h12):(5'h12)]) == $unsigned(reg328));
              reg2010 = reg307[(1'h0):(1'h0)];
            end
          if ((8'hb0))
            begin
              reg2013 = reg264[(2'h2):(1'h1)];
              reg2014 <= wire1999;
              reg2015 <= reg282;
              reg2016 = $unsigned(reg288);
              reg2017 <= $unsigned(($unsigned(reg264) ?
                  reg320[(4'he):(4'ha)] : $unsigned($signed((+reg257)))));
              reg2018 = $unsigned((^~$unsigned(((~^(8'hae)) ?
                  $unsigned(reg415) : reg362[(3'h5):(1'h0)]))));
              reg2019 = reg388;
            end
          else
            begin
              reg2012 <= reg327[(5'h12):(2'h2)];
              reg2013 = $unsigned(((($signed(reg331) == $unsigned(reg295)) ?
                      (!reg420) : ($signed(reg2009) ?
                          $unsigned(reg302) : reg390[(4'h8):(3'h7)])) ?
                  reg2005[(5'h11):(1'h0)] : reg331[(5'h12):(5'h10)]));
            end
          if (reg2012)
            begin
              reg2020 <= ($unsigned(reg345[(3'h6):(3'h5)]) || (-$unsigned($unsigned({reg314,
                  reg385}))));
              reg2021 = $signed((^~reg2008));
              reg2022 <= reg248[(4'hb):(4'h9)];
              reg2023 = ($unsigned((^wire227[(1'h0):(1'h0)])) >> $signed($signed(reg288)));
              reg2024 <= (7'h52);
            end
          else
            begin
              reg2021 = ($signed((reg2021 ?
                      $signed($signed(reg2023)) : reg299)) ?
                  ($unsigned(reg325) ?
                      $unsigned((8'ha5)) : wire229[(5'h16):(2'h2)]) : ($unsigned((^~$unsigned(reg381))) ~^ reg358[(3'h7):(1'h1)]));
              reg2023 = wire293[(1'h0):(1'h0)];
            end
          for (forvar2025 = (1'h0); (forvar2025 < (2'h3)); forvar2025 = (forvar2025 + (1'h1)))
            begin
              reg2026 = {reg327};
              reg2027 = $unsigned(({($signed(reg303) <= reg327[(1'h0):(1'h0)]),
                      reg253[(4'h9):(1'h0)],
                      ($signed(reg401) ? (~reg426) : $signed(reg2021))} ?
                  reg426[(3'h4):(1'h1)] : reg273[(3'h5):(1'h1)]));
              reg2028 = $unsigned((~|reg300));
              reg2029 <= $signed($unsigned((($signed((8'h9c)) <<< $unsigned(reg299)) >= {reg423[(3'h6):(3'h5)],
                  {reg287},
                  $unsigned(reg231)})));
            end
          for (forvar2030 = (1'h0); (forvar2030 < (1'h1)); forvar2030 = (forvar2030 + (1'h1)))
            begin
              reg2031 <= $unsigned(reg391);
              reg2032 = $unsigned(reg397[(2'h3):(2'h3)]);
            end
        end
      if (({$signed(((reg316 >>> (8'h9e)) || reg240)),
          {reg2021},
          ((reg247[(4'he):(4'h8)] ? reg2028 : $signed(reg239)) ?
              (~|(!reg336)) : (reg403 & wire291))} & reg279[(4'h9):(3'h4)]))
        begin
          reg2033 = ($signed(reg403[(5'h15):(4'h9)]) ?
              (((^(+reg2024)) << reg304) ~^ (|(8'hbf))) : $unsigned(($signed((reg240 > reg332)) > ((forvar2030 ?
                  reg314 : reg2031) << reg2020))));
          reg2034 = forvar2030;
          if ($signed((^reg295[(1'h0):(1'h0)])))
            begin
              reg2035 <= (7'h45);
              reg2036 <= $unsigned(($unsigned(reg381) ?
                  $unsigned(($unsigned(reg295) ?
                      reg317[(3'h7):(3'h7)] : wire319)) : (((+reg320) ?
                      ((7'h44) ?
                          reg412 : reg2014) : reg243) || reg295[(3'h6):(1'h0)])));
              reg2037 = {$unsigned(((~&reg246) ?
                      (reg312 | wire228[(3'h5):(2'h3)]) : reg421[(4'hb):(2'h2)])),
                  $unsigned({reg343}),
                  (~|({(reg2022 ? reg299 : reg231),
                          $unsigned(reg2020),
                          ((7'h4b) >= reg257)} ?
                      {reg316, (reg2029 ? (8'hbe) : (7'h58))} : (~|((8'ha9) ?
                          reg302 : reg311))))};
              reg2038 = {((reg430[(2'h2):(1'h0)] ?
                          reg264[(1'h0):(1'h0)] : ({reg2020,
                              reg430,
                              reg2012} ^ (^~reg403))) ?
                      (~(~|$unsigned(reg2008))) : {($signed(reg432) ?
                              reg432 : reg2013),
                          ({(7'h55)} << $unsigned(reg2037)),
                          $signed((7'h55))}),
                  $signed($signed((reg2019 ?
                      (reg331 ? reg299 : reg279) : reg392))),
                  $signed({reg432, $signed((reg2011 > wire1997))})};
              reg2039 <= $unsigned(reg2010);
            end
          else
            begin
              reg2035 <= reg2033[(5'h15):(2'h3)];
              reg2037 = ((8'h9d) ?
                  ((($signed((8'hb1)) || (reg262 >> reg2015)) > reg2020) && ((&$signed(reg400)) ?
                      (~&reg2008[(1'h1):(1'h0)]) : (reg432 ?
                          {(7'h45)} : $unsigned(reg353)))) : ({(~reg353),
                      reg242,
                      {$unsigned(reg351)}} - ((!reg2034[(3'h7):(3'h4)]) != $signed($unsigned(reg274)))));
            end
        end
      else
        begin
          reg2035 <= reg287[(4'hf):(4'hb)];
          if ({$signed(((~reg2011) <= ($unsigned(forvar2030) == $unsigned(reg2006)))),
              $signed({(~^reg2031[(4'h8):(1'h1)]),
                  (~&$unsigned(reg2034)),
                  reg394}),
              reg247[(5'h12):(4'he)]})
            begin
              reg2037 = $unsigned(({({reg317, reg296, (7'h4b)} ?
                      (reg282 != (8'ha4)) : ((8'hb5) ? reg2006 : reg2014)),
                  $unsigned((wire229 < reg2037)),
                  $unsigned((reg231 ~^ reg272))} ~^ (~reg325)));
            end
          else
            begin
              reg2037 = ((reg238 ?
                  ($signed((7'h4c)) * (7'h51)) : $unsigned(wire292[(3'h6):(2'h3)])) | $unsigned((reg2035 <= (^reg2009))));
              reg2038 = ((($signed({reg317,
                          reg2012,
                          reg2037}) != $unsigned((7'h55))) ?
                      $signed({reg2021,
                          $unsigned(reg2003),
                          (~^reg2024)}) : ($unsigned($unsigned(reg331)) ?
                          (~$signed(reg378)) : ((reg262 != reg371) << reg388))) ?
                  $signed((($unsigned((8'hab)) != $unsigned(reg2002)) != (~^(reg413 > reg2011)))) : $signed(($unsigned($unsigned(reg320)) ?
                      reg378[(2'h2):(2'h2)] : ((7'h49) <<< reg252))));
              reg2039 <= reg295[(2'h2):(1'h1)];
              reg2040 = ((~&(({(8'ha7),
                          wire229,
                          reg246} >> reg2009[(1'h1):(1'h1)]) ?
                      $signed((reg279 ? wire227 : wire319)) : {$signed(reg262),
                          $signed(reg296)})) ?
                  $unsigned((reg2013 ?
                      (reg332 ?
                          $signed(reg345) : (wire292 ?
                              wire1999 : reg301)) : $signed((reg406 ?
                          reg311 : reg343)))) : (~({reg412[(1'h0):(1'h0)]} ?
                      wire293 : reg232)));
              reg2041 <= (7'h56);
              reg2042 <= reg2022;
              reg2043 = (7'h45);
            end
          reg2044 <= (|(wire291[(1'h1):(1'h0)] ?
              {$signed((reg2011 <= reg280)),
                  (|$signed(reg2042))} : {(^~(reg330 <= wire227)),
                  $unsigned(reg358[(2'h3):(1'h1)])}));
        end
      if ((|reg2033))
        begin
          reg2045 <= $signed((8'ha0));
          reg2046 <= (-(~$signed(reg378[(2'h2):(1'h1)])));
          if ({(7'h50), reg296})
            begin
              reg2047 = $signed((~&{(!reg330)}));
              reg2048 = reg358[(3'h6):(3'h4)];
              reg2049 <= ({$signed($unsigned(((8'had) <= reg371))),
                  (~$unsigned(reg2016)),
                  (-((^~reg2034) ?
                      $unsigned(reg2032) : {(8'ha3),
                          reg2007}))} | ($unsigned((~|((7'h4c) ?
                  reg400 : reg417))) | (~^(^~$unsigned(reg2010)))));
              reg2050 = $signed($unsigned({(+reg304[(1'h0):(1'h0)])}));
              reg2051 = $signed($signed(((-$signed(wire227)) <<< $signed((reg430 ?
                  reg404 : (7'h40))))));
              reg2052 = (7'h4c);
            end
          else
            begin
              reg2047 = $signed(((+(&(wire227 ?
                  (8'h9f) : (8'haf)))) != reg329));
              reg2049 <= $signed(wire291);
            end
          reg2053 = reg362[(5'h1a):(3'h4)];
          if (reg415[(3'h6):(3'h6)])
            begin
              reg2054 <= {$signed($signed($unsigned((reg334 ?
                      (7'h4f) : reg248))))};
              reg2055 = reg335;
              reg2056 <= reg430[(2'h3):(2'h3)];
              reg2057 = reg2031;
              reg2058 <= (reg2051 ?
                  $signed($unsigned($unsigned((reg301 ?
                      reg2053 : (7'h50))))) : reg2053[(1'h1):(1'h1)]);
              reg2059 = $signed(reg2016);
              reg2060 <= $unsigned($signed((7'h43)));
            end
          else
            begin
              reg2055 = $unsigned((((^~forvar2025) != ($signed(reg246) ?
                  $signed((8'hbf)) : (reg430 == reg2008))) | (~^$unsigned($unsigned(reg262)))));
              reg2056 <= reg250[(1'h1):(1'h1)];
              reg2058 <= $unsigned((~(~|reg2049[(4'ha):(3'h5)])));
            end
          reg2061 = $signed(reg327);
          reg2062 <= reg421;
        end
      else
        begin
          if (reg2059[(1'h1):(1'h1)])
            begin
              reg2045 <= ((-(|((reg409 & reg2007) ?
                      (7'h55) : reg327[(4'h8):(3'h4)]))) ?
                  reg2008 : (~^$signed(reg2023)));
              reg2047 = (((reg2028 & {$unsigned(reg2051),
                          reg355[(3'h7):(2'h3)]}) ?
                      wire2000[(4'hd):(2'h2)] : ($unsigned($signed(reg274)) ?
                          $signed($signed(reg2005)) : ((~|reg2004) ?
                              (8'hb7) : (reg343 ? reg381 : (7'h58))))) ?
                  (reg2034[(4'hd):(1'h1)] << (+$unsigned((reg2028 ?
                      reg253 : reg317)))) : (!reg362[(5'h11):(3'h7)]));
              reg2048 = $signed(reg281);
              reg2049 <= reg351[(4'he):(2'h2)];
              reg2050 = {(~|$unsigned((~&reg2045))),
                  $unsigned(reg273[(4'hc):(1'h1)]),
                  (8'ha0)};
              reg2054 <= reg2027[(5'h1a):(5'h12)];
              reg2055 = reg2035;
            end
          else
            begin
              reg2047 = reg2022;
              reg2049 <= {($signed($unsigned(reg2034[(4'hd):(4'ha)])) <= $signed((+$unsigned(reg2012)))),
                  {$signed(reg2039),
                      {(|$signed(reg355))},
                      ((7'h4e) ?
                          ((reg397 * reg2058) <<< (!reg342)) : $signed((reg2004 ^~ reg2062)))}};
              reg2054 <= ($unsigned($signed(((+wire225) ?
                  reg2005[(5'h15):(5'h12)] : (reg408 + (7'h4a))))) != {(&$signed(((8'hb9) ?
                      reg2018 : (8'ha3))))});
              reg2055 = $signed(reg2027[(4'ha):(4'h9)]);
            end
          reg2056 <= reg420[(5'h11):(1'h1)];
        end
      reg2063 <= {reg391,
          {({reg328[(3'h6):(1'h0)],
                  (reg2059 != reg2052)} > (~wire319[(1'h1):(1'h0)])),
              $signed($signed(reg2001[(4'he):(4'hc)]))},
          ((reg2024 ? $unsigned((&reg2020)) : $unsigned($signed(reg311))) ?
              (reg274[(3'h5):(2'h3)] ?
                  $unsigned(reg2048[(3'h6):(1'h1)]) : (-{reg2060,
                      reg426,
                      reg320})) : reg336[(5'h1e):(4'hb)])};
      if ((reg311[(4'h8):(3'h7)] ?
          ($unsigned(reg2007) ?
              $unsigned(({(8'hb4)} ?
                  ((7'h50) << (8'hb4)) : (forvar2030 * reg2004))) : ($signed((forvar2025 ?
                      reg231 : reg362)) ?
                  (-(reg273 <<< reg303)) : (((8'h9c) ?
                      reg408 : reg400) ^ reg238[(3'h4):(3'h4)]))) : $unsigned($unsigned($unsigned((&reg2018))))))
        begin
          reg2064 <= (reg242 ?
              (+$signed((-$unsigned(reg335)))) : $signed($signed({(&reg288),
                  reg348})));
          for (forvar2065 = (1'h0); (forvar2065 < (3'h5)); forvar2065 = (forvar2065 + (1'h1)))
            begin
              reg2066 <= ({reg2007,
                      (wire293[(1'h1):(1'h1)] >= ($signed((7'h41)) & reg2053[(3'h7):(3'h6)]))} ?
                  $signed(((^~{reg325,
                      reg328,
                      reg274}) << reg2011)) : $unsigned({(&$signed(reg2050)),
                      $signed(reg307[(2'h3):(2'h2)]),
                      reg328[(4'hd):(2'h2)]}));
              reg2067 <= $unsigned(($unsigned(reg2062[(5'h10):(1'h1)]) == $signed(({wire227,
                      reg274,
                      reg2045} ?
                  $unsigned(wire1999) : (reg385 <= (8'hb8))))));
              reg2068 = $signed($signed($signed((+reg314[(3'h4):(2'h3)]))));
              reg2069 = reg2054[(1'h1):(1'h1)];
              reg2070 = (&((((reg274 * forvar2065) ?
                      reg408[(4'hc):(3'h6)] : ((8'hbd) ~^ reg2046)) < wire225) ?
                  ((reg2039 ^~ $signed(reg420)) ?
                      {reg2067[(2'h3):(1'h0)],
                          (reg409 ?
                              reg295 : reg2002)} : (^~reg2006[(5'h15):(4'ha)])) : reg232));
              reg2071 <= reg371[(3'h5):(1'h0)];
              reg2072 <= wire1999[(3'h6):(2'h2)];
            end
          for (forvar2073 = (1'h0); (forvar2073 < (1'h1)); forvar2073 = (forvar2073 + (1'h1)))
            begin
              reg2074 <= $unsigned((reg252 ?
                  {((&reg232) << $unsigned(wire319)),
                      $unsigned(wire1999),
                      ($unsigned(reg2027) - (reg2012 ?
                          reg2061 : reg408))} : {reg385[(3'h5):(3'h5)],
                      reg405,
                      reg2005}));
              reg2075 = (^~reg332);
              reg2076 <= $unsigned($signed($unsigned((~&reg2038[(1'h1):(1'h0)]))));
              reg2077 = $unsigned($signed((^reg332)));
              reg2078 <= reg2070;
              reg2079 <= reg406;
            end
          reg2080 <= $signed(reg2028[(2'h3):(1'h1)]);
          for (forvar2081 = (1'h0); (forvar2081 < (1'h1)); forvar2081 = (forvar2081 + (1'h1)))
            begin
              reg2082 <= reg2067;
            end
        end
      else
        begin
          for (forvar2064 = (1'h0); (forvar2064 < (2'h2)); forvar2064 = (forvar2064 + (1'h1)))
            begin
              reg2065 <= reg362;
              reg2066 <= (^$unsigned($signed(((reg232 ^ wire292) >= $signed(reg404)))));
              reg2068 = $signed(reg2078[(5'h18):(1'h0)]);
              reg2071 <= (+reg278);
              reg2073 = (reg355[(1'h1):(1'h0)] > (^(($signed(wire1999) == reg2038[(1'h0):(1'h0)]) ^ ((~|reg2031) >>> (reg252 | reg362)))));
              reg2075 = (~^$signed($signed(((reg2044 ~^ (7'h45)) ?
                  $signed(reg2078) : $unsigned(reg2012)))));
            end
          for (forvar2076 = (1'h0); (forvar2076 < (2'h3)); forvar2076 = (forvar2076 + (1'h1)))
            begin
              reg2077 = $signed($unsigned((-$unsigned($signed(reg403)))));
              reg2081 = (|($unsigned(reg242[(3'h7):(2'h2)]) || $signed(reg421[(5'h1c):(5'h13)])));
              reg2082 <= reg2024;
              reg2083 <= $unsigned(reg431);
              reg2084 <= (+reg232);
              reg2085 <= (|(reg284[(4'hb):(2'h2)] ?
                  reg412[(2'h3):(1'h0)] : reg2035));
            end
          for (forvar2086 = (1'h0); (forvar2086 < (1'h1)); forvar2086 = (forvar2086 + (1'h1)))
            begin
              reg2087 = $signed((|reg2035));
              reg2088 = {reg2056[(4'h8):(3'h6)],
                  (((|(reg2010 ^~ (8'hbd))) ?
                          $signed($unsigned(reg2012)) : (-((7'h56) > reg277))) ?
                      (~^reg252) : ($signed({reg329, reg423, reg2056}) ?
                          reg280[(3'h4):(1'h1)] : reg2069[(4'ha):(4'h9)]))};
              reg2089 <= reg2073;
              reg2090 = ((reg272 ? (+reg351) : (7'h57)) ?
                  reg394[(5'h11):(4'he)] : $unsigned($unsigned((7'h4d))));
              reg2091 = ($signed(reg299) * $unsigned((reg2002 ?
                  (reg2051[(5'h10):(4'he)] ?
                      reg334 : (reg282 < reg246)) : $signed($unsigned(reg413)))));
              reg2092 = (($unsigned(($signed(reg295) ^~ reg327[(4'he):(1'h1)])) ?
                      reg417 : {(~(reg2071 * (8'hb8)))}) ?
                  ((reg2018[(4'hf):(4'hf)] <<< $unsigned((reg426 ~^ reg247))) | forvar2030[(5'h1c):(2'h3)]) : ((reg430 ?
                      ($signed(reg2016) >= {reg2021,
                          (8'h9f),
                          reg247}) : reg277) & (reg421[(5'h1c):(4'hb)] ^~ (~reg2001[(2'h3):(1'h0)]))));
              reg2093 <= (({reg2012[(5'h10):(4'hd)],
                      $unsigned((|reg2083))} >> ($signed((+reg408)) <= reg272)) ?
                  reg412[(2'h2):(2'h2)] : $unsigned((!$unsigned((reg2084 * reg2052)))));
            end
          for (forvar2094 = (1'h0); (forvar2094 < (2'h3)); forvar2094 = (forvar2094 + (1'h1)))
            begin
              reg2095 = ({reg2033,
                      ((reg2074 <= (7'h42)) ?
                          $unsigned((+reg2039)) : (^~(reg378 ?
                              reg2044 : reg2047)))} ?
                  {$signed((reg2033[(3'h7):(2'h2)] <= ((8'ha8) < forvar2094))),
                      (reg390[(3'h6):(1'h0)] ?
                          ((~reg272) >= (reg2017 <<< (7'h45))) : $signed((reg252 < reg257))),
                      reg421[(5'h1d):(3'h5)]} : (reg284[(5'h11):(4'hf)] ?
                      forvar2094 : ($signed($signed(reg2012)) ?
                          $signed(reg342) : (((8'ha7) ? forvar2030 : reg2090) ?
                              reg2022 : ((8'h9c) || (7'h58))))));
            end
          reg2096 <= $signed(reg334);
        end
      reg2097 = ((&reg2084) >>> reg2070);
    end
  assign wire2098 = $signed({$unsigned((8'ha2)),
                        (^~(((8'hb8) ? reg334 : reg334) != (reg2029 ?
                            reg351 : reg335))),
                        ((reg281 || $unsigned(reg2031)) <<< reg2079[(3'h4):(1'h0)])});
  always
    @(posedge clk) begin
      reg2099 = (((reg242[(1'h0):(1'h0)] >> (8'hb4)) | reg320) ?
          $signed((&(!reg353[(1'h0):(1'h0)]))) : (~^reg2084));
      if ((^(reg2060[(2'h3):(1'h0)] <= $unsigned(($unsigned(reg2002) ?
          (reg331 <= (8'hb1)) : reg2058[(3'h4):(2'h3)])))))
        begin
          for (forvar2100 = (1'h0); (forvar2100 < (1'h1)); forvar2100 = (forvar2100 + (1'h1)))
            begin
              reg2101 <= ($unsigned((($signed((8'hb2)) ?
                  $signed(reg2084) : $unsigned(wire1999)) & (&{reg391}))) ^ ((reg243 ?
                      reg296 : reg2020[(4'h8):(3'h7)]) ?
                  (!wire2000) : (8'hba)));
              reg2102 <= $signed((+reg240));
            end
          if ((~^$unsigned((~$unsigned(reg243[(3'h6):(2'h2)])))))
            begin
              reg2103 = reg307;
              reg2104 <= $unsigned({reg403[(1'h1):(1'h0)],
                  (({reg2020, reg257, (7'h57)} ?
                      (wire228 ?
                          reg253 : reg381) : $unsigned(reg394)) & reg358),
                  (!(-$unsigned(reg281)))});
              reg2105 = (&reg279);
              reg2106 <= $unsigned((($signed(reg2065) > reg2062[(4'hf):(4'hf)]) ?
                  reg390 : reg2082));
              reg2107 <= reg2045[(2'h3):(1'h1)];
              reg2108 <= (+(^wire291[(1'h1):(1'h0)]));
            end
          else
            begin
              reg2103 = ($signed($unsigned((7'h51))) && reg420);
              reg2105 = ((reg252[(4'he):(1'h0)] ?
                  reg307 : ($signed((reg242 && (7'h52))) ?
                      reg2065 : (8'ha7))) & (reg2108 ?
                  $signed((8'hb9)) : wire227));
              reg2106 <= (!(~|$unsigned(reg2063[(1'h0):(1'h0)])));
              reg2109 = $unsigned($signed(($unsigned((reg280 ?
                  (8'ha9) : (7'h40))) <= $unsigned((reg358 ?
                  reg384 : reg2089)))));
              reg2110 = $unsigned((&$unsigned(((+reg343) ~^ {reg248}))));
              reg2111 <= $signed(wire225[(3'h7):(2'h3)]);
              reg2112 <= {(((~|(reg355 ? reg2002 : wire292)) ?
                          reg2011[(4'h8):(1'h1)] : reg252) ?
                      (&reg278[(4'h9):(4'h9)]) : $unsigned(((^~reg2049) ?
                          (^reg2058) : reg2110[(1'h1):(1'h0)])))};
            end
          if ((~&reg2031))
            begin
              reg2113 = reg2020[(1'h1):(1'h1)];
            end
          else
            begin
              reg2114 <= ((&((7'h4e) >= ((reg2015 ? reg332 : reg2039) ?
                  (&reg2083) : reg238))) || (7'h4b));
            end
          reg2115 <= reg2096[(4'h8):(2'h2)];
          reg2116 <= (^~$signed((reg2112 * ((~^reg401) <= (!reg2002)))));
        end
      else
        begin
          reg2100 <= (^~reg430[(2'h3):(2'h2)]);
          reg2103 = reg2106;
          reg2105 = {$unsigned(($signed((reg342 ?
                  (8'h9c) : reg2113)) | ((reg413 ? wire225 : reg317) ?
                  reg279 : $signed(wire2000)))),
              reg358};
          for (forvar2106 = (1'h0); (forvar2106 < (3'h6)); forvar2106 = (forvar2106 + (1'h1)))
            begin
              reg2107 <= reg432;
              reg2108 <= $unsigned(reg2014);
              reg2109 = $signed($signed($signed(reg253)));
              reg2110 = reg358[(2'h3):(2'h3)];
              reg2111 <= (-reg2002);
            end
        end
    end
  always
    @(posedge clk) begin
      reg2117 = ((reg2076[(2'h3):(2'h2)] ?
              reg295 : (&((8'had) ?
                  (~&reg2111) : (wire229 ? (7'h48) : reg2063)))) ?
          {$signed(reg401[(1'h1):(1'h1)])} : $signed(reg381));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module91  (y, clk, wire96, wire95, wire94, wire93, wire92);
  output wire [(32'h41):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire96;
  input wire signed [(5'h19):(1'h0)] wire95;
  input wire [(4'hc):(1'h0)] wire94;
  input wire [(5'h19):(1'h0)] wire93;
  input wire signed [(4'hc):(1'h0)] wire92;
  wire [(3'h6):(1'h0)] wire220;
  wire signed [(5'h18):(1'h0)] wire99;
  wire signed [(3'h7):(1'h0)] wire98;
  wire [(5'h1b):(1'h0)] wire97;
  assign y = {wire220, wire99, wire98, wire97, (1'h0)};
  assign wire97 = (($unsigned((wire96 >>> $signed(wire92))) ?
                          {wire93[(1'h1):(1'h1)]} : (~^(&(wire95 - wire93)))) ?
                      (8'ha6) : {wire94, (wire93[(5'h14):(3'h5)] << wire95)});
  assign wire98 = wire93;
  assign wire99 = $unsigned($signed(((7'h40) < (wire93[(4'hb):(1'h1)] || $unsigned(wire95)))));
  module100 #() modinst221 (wire220, clk, wire99, wire94, wire97, wire95, wire92, wire96);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module100
#(parameter param218 = ((~^({((7'h42) ? (8'hb2) : (7'h4c)), ((8'hbb) ? (8'hb2) : (7'h56)), ((8'hba) ? (8'ha1) : (8'hbb))} > {{(8'hae)}, ((7'h42) | (8'hbc)), (^(8'hb5))})) ? {(({(8'hb7), (7'h54), (8'h9f)} >= ((8'ha1) ^ (7'h4e))) - (8'hbd))} : ((8'h9c) ^ (~&(-{(8'haa), (8'hbc)})))), 
parameter param219 = param218)
(y, clk, wire106, wire105, wire104, wire103, wire102, wire101);
  output wire [(32'h774):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h18):(1'h0)] wire106;
  input wire [(3'h7):(1'h0)] wire105;
  input wire [(5'h1b):(1'h0)] wire104;
  input wire [(5'h19):(1'h0)] wire103;
  input wire signed [(4'hc):(1'h0)] wire102;
  input wire [(2'h2):(1'h0)] wire101;
  wire signed [(4'hc):(1'h0)] wire217;
  wire signed [(5'h13):(1'h0)] wire216;
  wire [(4'hf):(1'h0)] wire215;
  wire signed [(4'hc):(1'h0)] wire214;
  wire [(5'h15):(1'h0)] wire196;
  wire [(2'h2):(1'h0)] wire107;
  reg signed [(4'hc):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg212 = (1'h0);
  reg [(5'h1c):(1'h0)] reg208 = (1'h0);
  reg signed [(4'he):(1'h0)] reg207 = (1'h0);
  reg [(3'h5):(1'h0)] reg206 = (1'h0);
  reg [(5'h12):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg197 = (1'h0);
  reg [(2'h2):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg191 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg189 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg186 = (1'h0);
  reg [(4'hc):(1'h0)] reg185 = (1'h0);
  reg [(5'h1a):(1'h0)] reg182 = (1'h0);
  reg [(5'h1c):(1'h0)] reg180 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg178 = (1'h0);
  reg [(5'h16):(1'h0)] reg175 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg172 = (1'h0);
  reg [(5'h12):(1'h0)] reg170 = (1'h0);
  reg [(2'h3):(1'h0)] reg169 = (1'h0);
  reg [(4'ha):(1'h0)] reg167 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg164 = (1'h0);
  reg [(5'h14):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg159 = (1'h0);
  reg [(3'h6):(1'h0)] reg157 = (1'h0);
  reg [(4'ha):(1'h0)] reg155 = (1'h0);
  reg [(5'h16):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg152 = (1'h0);
  reg [(5'h1c):(1'h0)] reg148 = (1'h0);
  reg [(5'h10):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg138 = (1'h0);
  reg [(5'h1b):(1'h0)] reg136 = (1'h0);
  reg [(5'h1d):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg132 = (1'h0);
  reg [(5'h1f):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg126 = (1'h0);
  reg [(5'h16):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg123 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg122 = (1'h0);
  reg [(5'h11):(1'h0)] reg118 = (1'h0);
  reg [(5'h1d):(1'h0)] reg117 = (1'h0);
  reg [(5'h11):(1'h0)] reg113 = (1'h0);
  reg [(4'he):(1'h0)] reg110 = (1'h0);
  reg [(5'h18):(1'h0)] reg108 = (1'h0);
  reg [(4'hb):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg210 = (1'h0);
  reg [(5'h12):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg205 = (1'h0);
  reg [(5'h19):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg202 = (1'h0);
  reg [(5'h13):(1'h0)] reg201 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar199 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar198 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg193 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg192 = (1'h0);
  reg [(5'h17):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar188 = (1'h0);
  reg [(4'hf):(1'h0)] reg184 = (1'h0);
  reg [(4'ha):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg181 = (1'h0);
  reg [(4'h8):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg177 = (1'h0);
  reg [(4'hf):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg174 = (1'h0);
  reg [(4'hb):(1'h0)] reg171 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar168 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar166 = (1'h0);
  reg [(5'h11):(1'h0)] forvar165 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg163 = (1'h0);
  reg [(5'h1e):(1'h0)] reg162 = (1'h0);
  reg [(5'h13):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg158 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg154 = (1'h0);
  reg [(5'h10):(1'h0)] reg151 = (1'h0);
  reg [(4'he):(1'h0)] reg150 = (1'h0);
  reg [(4'ha):(1'h0)] reg149 = (1'h0);
  reg [(3'h5):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg145 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg144 = (1'h0);
  reg [(3'h7):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar142 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg141 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg137 = (1'h0);
  reg [(4'he):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar133 = (1'h0);
  reg [(5'h17):(1'h0)] reg129 = (1'h0);
  reg [(4'hd):(1'h0)] reg128 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg127 = (1'h0);
  reg [(3'h4):(1'h0)] forvar124 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg121 = (1'h0);
  reg [(4'h8):(1'h0)] reg120 = (1'h0);
  reg [(4'he):(1'h0)] forvar119 = (1'h0);
  reg [(4'ha):(1'h0)] reg116 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg115 = (1'h0);
  reg [(4'h9):(1'h0)] reg114 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg112 = (1'h0);
  reg [(5'h1f):(1'h0)] reg111 = (1'h0);
  reg [(4'ha):(1'h0)] forvar109 = (1'h0);
  assign y = {wire217,
                 wire216,
                 wire215,
                 wire214,
                 wire196,
                 wire107,
                 reg213,
                 reg212,
                 reg208,
                 reg207,
                 reg206,
                 reg204,
                 reg197,
                 reg195,
                 reg194,
                 reg191,
                 reg189,
                 reg187,
                 reg186,
                 reg185,
                 reg182,
                 reg180,
                 reg178,
                 reg175,
                 reg173,
                 reg172,
                 reg170,
                 reg169,
                 reg167,
                 reg164,
                 reg160,
                 reg159,
                 reg157,
                 reg155,
                 reg153,
                 reg152,
                 reg148,
                 reg147,
                 reg139,
                 reg138,
                 reg136,
                 reg135,
                 reg132,
                 reg131,
                 reg130,
                 reg126,
                 reg125,
                 reg123,
                 reg122,
                 reg118,
                 reg117,
                 reg113,
                 reg110,
                 reg108,
                 reg211,
                 reg210,
                 reg209,
                 reg205,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 forvar199,
                 forvar198,
                 reg193,
                 reg192,
                 reg190,
                 forvar188,
                 reg184,
                 reg183,
                 reg181,
                 reg179,
                 reg177,
                 reg176,
                 reg174,
                 reg171,
                 forvar168,
                 forvar166,
                 forvar165,
                 reg163,
                 reg162,
                 reg161,
                 reg158,
                 reg156,
                 reg154,
                 reg151,
                 reg150,
                 reg149,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 forvar142,
                 reg141,
                 reg140,
                 reg137,
                 reg134,
                 forvar133,
                 reg129,
                 reg128,
                 reg127,
                 forvar124,
                 reg121,
                 reg120,
                 forvar119,
                 reg116,
                 reg115,
                 reg114,
                 reg112,
                 reg111,
                 forvar109,
                 (1'h0)};
  assign wire107 = {wire105[(3'h7):(2'h2)],
                       (&($signed(wire104) - (wire106 ?
                           wire104[(5'h14):(5'h14)] : (wire101 ?
                               wire102 : wire103)))),
                       (~|wire106[(4'hf):(4'hc)])};
  always
    @(posedge clk) begin
      reg108 <= $unsigned($signed($signed({$signed(wire107),
          ((7'h56) ? wire106 : (7'h4a))})));
      for (forvar109 = (1'h0); (forvar109 < (3'h6)); forvar109 = (forvar109 + (1'h1)))
        begin
          if ({((&(((8'ha8) && wire105) + (~|(8'hae)))) ?
                  wire103 : (((forvar109 ? wire104 : wire106) ?
                          $unsigned(reg108) : (~^wire107)) ?
                      (^~{wire101}) : ((wire106 - wire107) + $signed(forvar109)))),
              $signed(((wire104 ?
                  wire104 : (~&wire102)) * $unsigned((!(7'h54))))),
              (((|$signed(forvar109)) ~^ wire106) ^~ {($unsigned(reg108) >> $unsigned(forvar109)),
                  (wire103[(4'hb):(4'h9)] > (7'h4d)),
                  (&$unsigned(forvar109))})})
            begin
              reg110 <= $signed((reg108 ?
                  ((wire103[(4'hf):(3'h7)] ?
                          wire102[(3'h6):(1'h0)] : $signed(wire107)) ?
                      (|((7'h41) ?
                          (8'hbb) : wire103)) : $signed((reg108 <<< wire101))) : $unsigned(wire106)));
            end
          else
            begin
              reg110 <= reg110[(4'he):(4'h8)];
              reg111 = (^~reg110);
              reg112 = $signed($unsigned(wire101[(1'h1):(1'h1)]));
              reg113 <= $signed($signed(reg111));
              reg114 = (^((~|((~(7'h4d)) ?
                  wire103[(5'h11):(2'h3)] : (-reg113))) - reg110));
              reg115 = (reg114[(3'h4):(2'h3)] * forvar109);
              reg116 = ($unsigned(reg112[(1'h1):(1'h0)]) || {$signed($signed((~^(8'ha5)))),
                  reg115});
            end
          reg117 <= (reg115 ?
              $signed(((+(|forvar109)) ?
                  ((8'h9c) ~^ reg111[(3'h7):(1'h1)]) : (wire105 || {(8'hb8),
                      reg108,
                      reg108}))) : reg108[(5'h10):(4'hd)]);
          reg118 <= $signed(($unsigned({reg115}) ?
              (reg116[(3'h7):(1'h0)] << $signed((wire104 >>> forvar109))) : ((~|(^~wire101)) - reg111)));
          for (forvar119 = (1'h0); (forvar119 < (1'h0)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg120 = (7'h4c);
              reg121 = $unsigned(reg120[(3'h6):(3'h4)]);
              reg122 <= reg112[(4'h9):(1'h0)];
              reg123 <= (7'h58);
            end
          for (forvar124 = (1'h0); (forvar124 < (1'h1)); forvar124 = (forvar124 + (1'h1)))
            begin
              reg125 <= {reg120,
                  (wire103[(4'ha):(1'h0)] & $unsigned(($signed(wire104) >> (!reg123))))};
              reg126 <= $signed(wire102);
              reg127 = ($signed(($unsigned($unsigned(reg118)) ?
                      forvar109[(4'h8):(4'h8)] : $signed($signed(reg125)))) ?
                  $signed((~(reg126 ?
                      $signed(wire101) : $signed(forvar119)))) : ($signed(reg113) << ((~|((8'hba) ?
                      wire101 : (8'haf))) <<< (~(7'h47)))));
              reg128 = $signed(wire106[(5'h15):(5'h13)]);
              reg129 = (forvar124[(3'h4):(2'h3)] | (reg123[(5'h16):(5'h13)] ?
                  $signed({((8'had) * reg116)}) : $unsigned(((wire104 ^ reg123) != (reg125 ?
                      reg128 : reg114)))));
              reg130 <= (-{reg110[(4'hd):(4'hd)],
                  (((wire104 ? wire107 : reg128) <<< (reg112 ?
                      reg120 : wire103)) || ({reg114, (7'h48)} ?
                      $signed(reg122) : (^reg113)))});
              reg131 <= (+(~&wire107[(2'h2):(1'h0)]));
            end
          reg132 <= reg114;
        end
      for (forvar133 = (1'h0); (forvar133 < (3'h6)); forvar133 = (forvar133 + (1'h1)))
        begin
          reg134 = $unsigned(({$unsigned({wire103}),
                  $signed(reg108[(1'h1):(1'h1)]),
                  reg113[(4'hb):(4'ha)]} ?
              wire107 : $unsigned(((reg108 || (8'haf)) <= $unsigned((7'h4b))))));
          reg135 <= ((forvar124[(3'h4):(3'h4)] ?
              {forvar124,
                  ($unsigned((7'h46)) << wire104),
                  {$unsigned(wire102),
                      wire107[(2'h2):(2'h2)]}} : $unsigned(({forvar133,
                      reg120} ?
                  {reg134,
                      forvar119} : $signed(reg131)))) >>> (forvar109[(3'h7):(3'h7)] ?
              ($unsigned(reg127[(4'h8):(3'h4)]) ?
                  (^~$signed(reg121)) : $signed($unsigned(reg112))) : ((-$signed(reg125)) < (+(~&reg108)))));
          if ($unsigned(reg122))
            begin
              reg136 <= reg123[(3'h4):(2'h2)];
              reg137 = reg121[(4'he):(4'hd)];
              reg138 <= reg127;
              reg139 <= $unsigned(reg137);
              reg140 = forvar133[(4'hb):(4'h9)];
            end
          else
            begin
              reg137 = ((-$signed(($signed(reg110) < $signed(reg137)))) >> (|{{{reg127},
                      (reg114 - reg125),
                      (reg110 <<< (7'h55))}}));
              reg140 = ($signed(reg127) && ({$unsigned({forvar124,
                      reg129,
                      reg110}),
                  reg115[(3'h5):(3'h5)]} <= reg126));
              reg141 = $unsigned(forvar133[(5'h1d):(2'h3)]);
            end
          for (forvar142 = (1'h0); (forvar142 < (1'h0)); forvar142 = (forvar142 + (1'h1)))
            begin
              reg143 = $signed(wire103[(5'h17):(5'h15)]);
              reg144 = reg110;
              reg145 = (^(^reg136));
              reg146 = reg144[(2'h3):(1'h0)];
            end
          if ((reg135[(5'h14):(5'h11)] * reg135))
            begin
              reg147 <= (-$signed(({(reg114 ? wire106 : reg113),
                  (reg137 << (8'ha6))} > reg145[(5'h14):(4'hb)])));
              reg148 <= reg113;
              reg149 = $signed(reg108);
              reg150 = reg132[(2'h3):(2'h3)];
            end
          else
            begin
              reg149 = reg128[(4'h8):(3'h4)];
              reg150 = (reg141[(1'h1):(1'h1)] ?
                  ($unsigned($unsigned(forvar119)) ?
                      ($signed((~^reg138)) ?
                          (~^{reg145, reg121}) : {(|reg111),
                              reg135[(1'h0):(1'h0)]}) : $signed($unsigned((~reg111)))) : {(reg134[(4'he):(4'ha)] <<< reg117[(2'h3):(1'h1)]),
                      wire103[(4'hf):(2'h3)],
                      reg128});
              reg151 = reg150;
              reg152 <= (+(|$unsigned($signed((reg117 ? reg123 : reg118)))));
              reg153 <= ($signed($unsigned($signed((reg115 + (7'h46))))) + (reg114 ~^ $signed(((reg126 ?
                  reg141 : reg108) << (~|reg110)))));
            end
          if ((reg114[(3'h6):(2'h3)] ?
              $signed($signed($unsigned(forvar119))) : wire101))
            begin
              reg154 = $signed({reg113, wire101[(2'h2):(2'h2)]});
              reg155 <= $unsigned({reg132, reg118[(2'h3):(2'h2)]});
              reg156 = ({wire102[(3'h5):(3'h4)]} ?
                  ($signed(((reg120 || reg117) != reg115)) + reg108[(5'h15):(5'h10)]) : (|reg152));
              reg157 <= $unsigned(reg154[(2'h2):(1'h1)]);
              reg158 = ((((&reg127[(4'ha):(3'h5)]) ?
                      reg152[(5'h18):(4'hd)] : reg144[(3'h5):(1'h0)]) ?
                  reg118[(3'h4):(1'h0)] : (reg110 ?
                      $unsigned((reg115 <= (7'h4c))) : ((reg114 ?
                              reg138 : reg150) ?
                          (7'h53) : $unsigned(reg155)))) > (($signed(reg108) ?
                      $signed({reg154, (7'h46), wire104}) : reg154) ?
                  $unsigned(($unsigned(reg123) > reg123[(3'h6):(1'h1)])) : forvar142[(3'h5):(3'h4)]));
              reg159 <= (wire104[(1'h0):(1'h0)] ?
                  $signed(((&(reg150 ~^ reg145)) ?
                      (+(reg129 ^~ reg147)) : $unsigned($signed((7'h53))))) : $signed($signed($signed(reg117[(3'h7):(3'h6)]))));
              reg160 <= (reg159[(2'h3):(2'h2)] ?
                  reg132 : (|(-($signed(reg150) ?
                      $signed(reg144) : $signed(reg136)))));
            end
          else
            begin
              reg154 = $unsigned((($unsigned(reg154[(3'h6):(2'h2)]) ^ (((7'h41) - (7'h47)) ?
                  (~|reg132) : reg159)) - reg157));
              reg155 <= $signed(reg159[(5'h17):(3'h7)]);
              reg157 <= reg160;
              reg159 <= reg141;
              reg161 = $unsigned((-{reg139[(1'h0):(1'h0)]}));
              reg162 = (reg153[(5'h12):(4'hd)] ? (8'hbb) : reg114);
            end
        end
      reg163 = (((((+(7'h51)) ?
          (reg159 ?
              forvar142 : reg160) : $signed(reg134)) << reg153) + (reg141 ?
          $signed(reg147[(2'h3):(2'h3)]) : {(reg113 + forvar133)})) ^~ (-(wire103 ?
          ($unsigned(reg121) ? $unsigned(reg132) : {reg114}) : reg158)));
      reg164 <= (!({$unsigned($signed(reg146)),
              $signed(reg145),
              $signed((reg138 ? wire103 : reg151))} ?
          $signed($signed((reg162 > reg147))) : (reg120 ?
              (((7'h4f) ? reg135 : reg128) ?
                  (^~reg155) : reg145[(3'h7):(1'h1)]) : reg112)));
      for (forvar165 = (1'h0); (forvar165 < (1'h1)); forvar165 = (forvar165 + (1'h1)))
        begin
          for (forvar166 = (1'h0); (forvar166 < (3'h4)); forvar166 = (forvar166 + (1'h1)))
            begin
              reg167 <= wire104[(5'h17):(5'h10)];
            end
          for (forvar168 = (1'h0); (forvar168 < (2'h2)); forvar168 = (forvar168 + (1'h1)))
            begin
              reg169 <= {reg163};
              reg170 <= reg138;
              reg171 = reg115;
              reg172 <= reg112[(3'h4):(1'h0)];
              reg173 <= wire104;
            end
          if (reg140[(2'h2):(1'h1)])
            begin
              reg174 = (+reg144);
              reg175 <= ((+reg152[(4'he):(2'h3)]) ^ wire105[(3'h7):(2'h2)]);
              reg176 = reg129[(4'ha):(1'h1)];
              reg177 = wire107[(1'h1):(1'h0)];
            end
          else
            begin
              reg175 <= reg120;
              reg178 <= reg157;
              reg179 = ($unsigned((reg138[(5'h15):(5'h12)] ?
                  {wire104} : $signed($unsigned(reg173)))) || (($unsigned($unsigned(reg110)) ?
                  $signed($signed(reg130)) : ($unsigned(wire104) < (&(8'hbf)))) != reg141));
              reg180 <= (forvar133[(4'hf):(2'h3)] ?
                  reg167 : (reg149 ? reg139 : (8'h9e)));
            end
          if ((+(reg108 ?
              reg135[(5'h19):(5'h18)] : ($unsigned($unsigned((8'hba))) <<< reg167))))
            begin
              reg181 = reg146[(2'h2):(2'h2)];
              reg182 <= reg122;
              reg183 = ($signed((({reg146, reg148} & {(7'h51),
                      reg110,
                      reg118}) ?
                  forvar142[(5'h14):(5'h14)] : (~^$unsigned(forvar119)))) <= (8'h9e));
              reg184 = ($signed(reg162) ~^ (reg139 ~^ (8'ha8)));
            end
          else
            begin
              reg181 = (({(~^reg126[(2'h2):(1'h1)]),
                  reg120[(2'h2):(1'h0)]} * (reg173[(1'h1):(1'h1)] | $signed($unsigned((8'h9f))))) || {reg121[(3'h7):(2'h2)],
                  (reg108[(4'hb):(4'h9)] ?
                      $unsigned((reg134 ? reg121 : reg162)) : {$signed(wire106),
                          (reg154 > reg144)})});
              reg182 <= ((|reg118[(5'h10):(1'h0)]) ?
                  ($signed((+reg161)) & (reg173[(1'h1):(1'h0)] ?
                      (-(~reg132)) : (+{reg114,
                          reg162}))) : $unsigned((|$unsigned(wire105[(3'h5):(2'h2)]))));
              reg183 = {$unsigned((((wire102 ?
                          reg118 : (8'hb7)) >>> wire107[(1'h0):(1'h0)]) ?
                      reg139[(5'h19):(3'h6)] : (reg172 ?
                          reg123[(5'h10):(4'h9)] : {reg108, reg136, reg176}))),
                  (((+(reg110 * wire104)) ?
                          reg150[(4'hd):(3'h7)] : reg169[(2'h3):(1'h1)]) ?
                      reg177 : {(~^((8'hbb) ? reg157 : (7'h50))),
                          (reg111[(5'h1b):(4'h8)] ?
                              (reg141 ? reg115 : reg138) : ((8'ha1) ?
                                  reg178 : (8'h9d))),
                          $signed(((7'h49) ^~ (7'h4c)))})};
              reg185 <= (($signed((!(reg134 ? reg162 : wire106))) ?
                      reg181 : ($signed(reg137[(5'h13):(3'h4)]) + ($signed(reg156) ?
                          (wire107 & forvar166) : reg146))) ?
                  ((7'h43) >> $signed(((~^reg153) ?
                      (reg141 != reg184) : $unsigned(reg184)))) : (((~(^~forvar109)) ?
                      ($unsigned((7'h4a)) ?
                          $signed((7'h52)) : reg125[(4'hc):(1'h1)]) : {(reg134 != reg151)}) | (({reg156} ?
                          reg177[(4'he):(4'h8)] : reg164[(1'h0):(1'h0)]) ?
                      ((reg125 ?
                          forvar109 : reg140) << $signed(reg130)) : ((^(8'ha4)) ?
                          $unsigned(reg145) : reg143))));
              reg186 <= wire105;
              reg187 <= (~&($signed(reg116) || ($signed((reg130 ?
                      reg182 : wire107)) ?
                  reg184 : $unsigned({(8'hb6)}))));
            end
          for (forvar188 = (1'h0); (forvar188 < (3'h4)); forvar188 = (forvar188 + (1'h1)))
            begin
              reg189 <= reg111[(5'h11):(4'hf)];
              reg190 = reg164;
              reg191 <= (^$unsigned((reg157[(3'h4):(1'h1)] ?
                  ($unsigned(forvar142) ?
                      $signed(wire102) : (|reg176)) : ((reg131 ?
                      reg177 : (8'h9e)) < ((8'haa) ? reg149 : reg126)))));
              reg192 = $signed((8'hae));
              reg193 = $unsigned(($signed(reg112) ?
                  ($signed(forvar124[(1'h1):(1'h1)]) ?
                      (~|((8'ha7) >> reg117)) : (~&reg164)) : forvar188));
              reg194 <= reg150[(4'hd):(2'h3)];
              reg195 <= reg153[(5'h15):(4'h8)];
            end
        end
    end
  assign wire196 = (8'h9d);
  always
    @(posedge clk) begin
      reg197 <= {$signed((|reg185))};
      for (forvar198 = (1'h0); (forvar198 < (2'h3)); forvar198 = (forvar198 + (1'h1)))
        begin
          for (forvar199 = (1'h0); (forvar199 < (1'h0)); forvar199 = (forvar199 + (1'h1)))
            begin
              reg200 = reg125;
              reg201 = $signed($unsigned((reg187 ?
                  reg148[(1'h1):(1'h1)] : $unsigned({(8'h9e)}))));
              reg202 = $unsigned($unsigned((((|reg125) - wire106[(5'h13):(4'h8)]) ?
                  wire196[(4'h9):(3'h4)] : (8'hbe))));
            end
          reg203 = reg113[(3'h4):(1'h0)];
          if ($signed($signed(wire196)))
            begin
              reg204 <= ($unsigned($signed((&reg191))) < reg136);
              reg205 = $signed($unsigned(reg157[(2'h2):(1'h1)]));
              reg206 <= ({reg185[(4'hb):(3'h6)]} <= {(~&reg204[(3'h5):(1'h0)]),
                  reg135[(4'hf):(3'h6)]});
              reg207 <= reg130;
              reg208 <= ((((wire101 ?
                      reg132[(1'h1):(1'h0)] : (reg206 ?
                          (8'ha2) : reg130)) <= (reg152[(5'h12):(3'h5)] && reg202)) ?
                  $signed(($signed(reg182) ?
                      (!wire103) : reg113[(3'h4):(1'h0)])) : {(~&reg180[(3'h4):(1'h0)])}) ~^ $unsigned((forvar199 ^ ((reg139 ?
                  (7'h45) : reg123) * $unsigned((8'hb1))))));
            end
          else
            begin
              reg205 = (^~reg164);
              reg206 <= $signed(wire105);
              reg207 <= ((8'haa) ^ ($unsigned({(reg123 ? reg117 : reg170)}) ?
                  $unsigned($signed(reg132)) : (8'h9f)));
              reg209 = ((($signed(reg138[(4'hb):(2'h3)]) ?
                      reg130 : (~^$unsigned(reg180))) * $signed((~&reg200[(1'h0):(1'h0)]))) ?
                  ((($signed(reg147) >>> $signed(reg130)) ?
                          ($signed(reg126) ?
                              $signed(reg204) : reg185) : ($signed(reg118) ?
                              reg186[(2'h2):(2'h2)] : reg182[(4'hf):(3'h4)])) ?
                      $unsigned($signed($signed(reg191))) : $unsigned((reg138[(4'he):(3'h5)] ?
                          $unsigned(reg117) : reg194))) : $unsigned({(^~(~^reg148)),
                      $signed(reg125[(4'he):(4'hc)]),
                      {(reg125 >> reg197), (~reg178)}}));
              reg210 = $unsigned((reg167[(3'h5):(3'h5)] - reg182));
              reg211 = {$unsigned((((reg164 >= reg131) + {reg108}) > (+(!reg147)))),
                  ((~reg172[(3'h4):(1'h0)]) <= reg197[(3'h7):(2'h3)])};
            end
        end
      reg212 <= {(-reg202), reg187, wire106[(5'h18):(5'h14)]};
      reg213 <= (7'h4e);
    end
  assign wire214 = (($signed(((reg123 ? reg164 : reg213) ?
                           (reg208 ?
                               reg152 : reg138) : (wire107 != reg125))) <<< $unsigned(wire196[(2'h2):(1'h0)])) ?
                       (((reg136 ^ $unsigned(wire105)) ? reg157 : reg139) ?
                           (reg197[(4'hd):(4'hd)] ?
                               ($signed(reg187) && (reg186 && reg169)) : $signed(reg170[(3'h6):(1'h0)])) : {$signed(((8'ha9) ?
                                   reg139 : reg147))}) : (reg213 >= $signed((|$unsigned((8'haf))))));
  assign wire215 = (~|reg159[(5'h12):(5'h10)]);
  assign wire216 = (reg160 != $signed($signed((reg175 * (7'h4b)))));
  assign wire217 = $unsigned(reg138[(4'hf):(3'h4)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module434
#(parameter param1995 = (((({(8'hbb)} ? ((7'h4d) | (7'h4a)) : ((7'h58) > (7'h4b))) >> {{(8'ha9), (8'ha6), (8'ha5)}, ((7'h44) ? (8'ha5) : (7'h4b)), ((8'ha4) << (7'h54))}) ^~ (&((!(7'h43)) ? {(8'ha9), (7'h57), (8'hbe)} : (&(8'hb0))))) < ((&(-{(8'ha9), (7'h55), (8'hae)})) >>> {(&(~&(8'hba)))})), 
parameter param1996 = (param1995 & (((param1995 ? (!param1995) : (~param1995)) != param1995) <= ((~&(!param1995)) ? ({param1995, param1995} < {param1995, (8'h9e)}) : param1995))))
(y, clk, wire439, wire438, wire437, wire436, wire435);
  output wire [(32'h1f9e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire439;
  input wire signed [(5'h13):(1'h0)] wire438;
  input wire [(5'h14):(1'h0)] wire437;
  input wire signed [(4'h9):(1'h0)] wire436;
  input wire [(3'h4):(1'h0)] wire435;
  wire signed [(4'he):(1'h0)] wire1993;
  wire signed [(2'h2):(1'h0)] wire1992;
  wire [(5'h16):(1'h0)] wire1990;
  wire signed [(3'h7):(1'h0)] wire1478;
  wire [(3'h7):(1'h0)] wire1247;
  wire [(5'h14):(1'h0)] wire1246;
  wire [(4'hb):(1'h0)] wire1244;
  wire signed [(5'h16):(1'h0)] wire1059;
  wire signed [(5'h1f):(1'h0)] wire860;
  wire signed [(5'h13):(1'h0)] wire838;
  wire signed [(4'hc):(1'h0)] wire542;
  reg [(5'h1b):(1'h0)] reg1994 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1386 = (1'h0);
  reg [(5'h10):(1'h0)] reg1381 = (1'h0);
  reg [(2'h2):(1'h0)] reg1380 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1353 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1378 = (1'h0);
  reg [(4'hc):(1'h0)] reg1377 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1374 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1372 = (1'h0);
  reg [(5'h11):(1'h0)] reg1369 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1368 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1366 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1362 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1361 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1360 = (1'h0);
  reg [(5'h15):(1'h0)] reg1356 = (1'h0);
  reg [(2'h3):(1'h0)] reg1355 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1354 = (1'h0);
  reg [(5'h10):(1'h0)] reg1352 = (1'h0);
  reg [(4'hf):(1'h0)] reg1350 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1346 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1345 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1344 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1341 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1339 = (1'h0);
  reg [(3'h6):(1'h0)] reg1337 = (1'h0);
  reg [(4'h8):(1'h0)] reg1335 = (1'h0);
  reg [(4'hd):(1'h0)] reg1334 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1331 = (1'h0);
  reg [(5'h17):(1'h0)] reg1330 = (1'h0);
  reg [(3'h5):(1'h0)] reg1327 = (1'h0);
  reg [(5'h11):(1'h0)] reg1323 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1322 = (1'h0);
  reg [(5'h15):(1'h0)] reg1320 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1319 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1317 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1313 = (1'h0);
  reg [(5'h12):(1'h0)] reg1312 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1310 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1308 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1307 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1306 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1302 = (1'h0);
  reg [(5'h12):(1'h0)] reg1301 = (1'h0);
  reg [(4'h8):(1'h0)] reg1299 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1295 = (1'h0);
  reg [(5'h10):(1'h0)] reg1294 = (1'h0);
  reg [(4'hf):(1'h0)] reg1292 = (1'h0);
  reg [(3'h6):(1'h0)] reg1290 = (1'h0);
  reg [(4'hc):(1'h0)] reg1285 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1283 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1279 = (1'h0);
  reg [(3'h5):(1'h0)] reg1278 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1277 = (1'h0);
  reg [(3'h5):(1'h0)] reg1276 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1274 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1272 = (1'h0);
  reg [(2'h2):(1'h0)] reg1271 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1264 = (1'h0);
  reg [(5'h16):(1'h0)] reg1262 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1260 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1258 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1257 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1255 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1254 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1252 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1251 = (1'h0);
  reg [(2'h2):(1'h0)] reg1058 = (1'h0);
  reg [(5'h17):(1'h0)] reg1055 = (1'h0);
  reg [(4'he):(1'h0)] reg1051 = (1'h0);
  reg [(4'ha):(1'h0)] reg1049 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1047 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1046 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1041 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1040 = (1'h0);
  reg [(2'h2):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1037 = (1'h0);
  reg [(5'h12):(1'h0)] reg1036 = (1'h0);
  reg [(5'h13):(1'h0)] reg1033 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1031 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1030 = (1'h0);
  reg [(5'h14):(1'h0)] reg1027 = (1'h0);
  reg [(5'h14):(1'h0)] reg1022 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1021 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1020 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1017 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1016 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1004 = (1'h0);
  reg [(5'h11):(1'h0)] reg999 = (1'h0);
  reg [(5'h1b):(1'h0)] reg998 = (1'h0);
  reg [(5'h1e):(1'h0)] reg997 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg996 = (1'h0);
  reg [(5'h1d):(1'h0)] reg995 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg993 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg990 = (1'h0);
  reg [(5'h16):(1'h0)] reg989 = (1'h0);
  reg [(4'hd):(1'h0)] reg988 = (1'h0);
  reg [(2'h2):(1'h0)] reg985 = (1'h0);
  reg [(5'h19):(1'h0)] reg980 = (1'h0);
  reg [(3'h7):(1'h0)] reg978 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg977 = (1'h0);
  reg [(5'h1d):(1'h0)] reg976 = (1'h0);
  reg [(4'hf):(1'h0)] reg971 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg970 = (1'h0);
  reg [(5'h13):(1'h0)] reg968 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg963 = (1'h0);
  reg [(3'h5):(1'h0)] reg960 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg957 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg956 = (1'h0);
  reg [(4'hb):(1'h0)] reg951 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg950 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg949 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg945 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg942 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg941 = (1'h0);
  reg [(3'h4):(1'h0)] reg932 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg929 = (1'h0);
  reg [(5'h1d):(1'h0)] reg926 = (1'h0);
  reg [(5'h10):(1'h0)] reg919 = (1'h0);
  reg [(4'ha):(1'h0)] reg916 = (1'h0);
  reg [(2'h3):(1'h0)] reg910 = (1'h0);
  reg signed [(4'he):(1'h0)] reg909 = (1'h0);
  reg [(2'h3):(1'h0)] reg907 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg905 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg902 = (1'h0);
  reg [(4'h8):(1'h0)] reg900 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg898 = (1'h0);
  reg [(5'h14):(1'h0)] reg897 = (1'h0);
  reg [(4'hf):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg894 = (1'h0);
  reg [(3'h6):(1'h0)] reg891 = (1'h0);
  reg [(5'h17):(1'h0)] reg889 = (1'h0);
  reg [(5'h19):(1'h0)] reg888 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg887 = (1'h0);
  reg [(5'h1f):(1'h0)] reg885 = (1'h0);
  reg [(4'hd):(1'h0)] reg884 = (1'h0);
  reg [(5'h1b):(1'h0)] reg883 = (1'h0);
  reg [(4'h9):(1'h0)] reg878 = (1'h0);
  reg [(5'h1e):(1'h0)] reg877 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg876 = (1'h0);
  reg [(5'h15):(1'h0)] reg872 = (1'h0);
  reg signed [(4'he):(1'h0)] reg870 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg868 = (1'h0);
  reg [(5'h13):(1'h0)] reg867 = (1'h0);
  reg [(4'hb):(1'h0)] reg866 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg863 = (1'h0);
  reg [(5'h16):(1'h0)] reg861 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg857 = (1'h0);
  reg [(5'h11):(1'h0)] reg856 = (1'h0);
  reg [(5'h1f):(1'h0)] reg854 = (1'h0);
  reg [(4'hb):(1'h0)] reg850 = (1'h0);
  reg [(3'h6):(1'h0)] reg849 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg848 = (1'h0);
  reg [(4'hd):(1'h0)] reg845 = (1'h0);
  reg [(5'h19):(1'h0)] reg843 = (1'h0);
  reg [(3'h7):(1'h0)] reg842 = (1'h0);
  reg [(4'hf):(1'h0)] reg841 = (1'h0);
  reg [(4'hc):(1'h0)] reg840 = (1'h0);
  reg [(5'h11):(1'h0)] reg541 = (1'h0);
  reg [(3'h7):(1'h0)] reg537 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg536 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg533 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg530 = (1'h0);
  reg [(3'h6):(1'h0)] reg529 = (1'h0);
  reg [(3'h5):(1'h0)] reg528 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg524 = (1'h0);
  reg [(5'h10):(1'h0)] reg523 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg507 = (1'h0);
  reg [(5'h17):(1'h0)] reg521 = (1'h0);
  reg [(5'h1b):(1'h0)] reg520 = (1'h0);
  reg [(4'hf):(1'h0)] reg517 = (1'h0);
  reg [(5'h17):(1'h0)] reg516 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg514 = (1'h0);
  reg [(5'h14):(1'h0)] reg511 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg510 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg503 = (1'h0);
  reg [(4'h9):(1'h0)] reg502 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg498 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg495 = (1'h0);
  reg [(3'h6):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg491 = (1'h0);
  reg [(5'h1c):(1'h0)] reg489 = (1'h0);
  reg [(5'h18):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg485 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg484 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg482 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg480 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg479 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg478 = (1'h0);
  reg [(5'h14):(1'h0)] reg477 = (1'h0);
  reg [(3'h6):(1'h0)] reg476 = (1'h0);
  reg signed [(4'he):(1'h0)] reg473 = (1'h0);
  reg [(3'h5):(1'h0)] reg471 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg470 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg469 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg468 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg467 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg466 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg465 = (1'h0);
  reg [(5'h1f):(1'h0)] reg464 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg463 = (1'h0);
  reg [(5'h1e):(1'h0)] reg461 = (1'h0);
  reg [(5'h1c):(1'h0)] reg457 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg452 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg448 = (1'h0);
  reg signed [(4'he):(1'h0)] reg446 = (1'h0);
  reg [(3'h4):(1'h0)] reg444 = (1'h0);
  reg [(5'h18):(1'h0)] reg443 = (1'h0);
  reg [(5'h1d):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg441 = (1'h0);
  reg [(5'h13):(1'h0)] reg1385 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1384 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1383 = (1'h0);
  reg [(3'h6):(1'h0)] reg1382 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1371 = (1'h0);
  reg [(3'h6):(1'h0)] reg1363 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1379 = (1'h0);
  reg [(4'hf):(1'h0)] reg1376 = (1'h0);
  reg [(4'hb):(1'h0)] reg1375 = (1'h0);
  reg [(5'h18):(1'h0)] reg1373 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1371 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1370 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1367 = (1'h0);
  reg [(2'h2):(1'h0)] reg1365 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1364 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1363 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1359 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1358 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1357 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1353 = (1'h0);
  reg [(5'h12):(1'h0)] reg1351 = (1'h0);
  reg [(5'h10):(1'h0)] reg1349 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1348 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1347 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1343 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1342 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1340 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1338 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1336 = (1'h0);
  reg [(3'h6):(1'h0)] reg1333 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1332 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1329 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1328 = (1'h0);
  reg [(5'h18):(1'h0)] reg1328 = (1'h0);
  reg [(3'h4):(1'h0)] reg1326 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1325 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1324 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1321 = (1'h0);
  reg [(5'h15):(1'h0)] reg1318 = (1'h0);
  reg [(3'h4):(1'h0)] reg1316 = (1'h0);
  reg [(2'h2):(1'h0)] reg1315 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1314 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1311 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1309 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1305 = (1'h0);
  reg [(4'hd):(1'h0)] reg1304 = (1'h0);
  reg [(3'h7):(1'h0)] reg1303 = (1'h0);
  reg [(4'he):(1'h0)] reg1300 = (1'h0);
  reg [(2'h2):(1'h0)] reg1298 = (1'h0);
  reg [(5'h17):(1'h0)] reg1297 = (1'h0);
  reg [(4'he):(1'h0)] reg1296 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1293 = (1'h0);
  reg [(5'h19):(1'h0)] reg1291 = (1'h0);
  reg [(2'h2):(1'h0)] reg1289 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1288 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1287 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1286 = (1'h0);
  reg [(5'h10):(1'h0)] reg1284 = (1'h0);
  reg [(5'h12):(1'h0)] reg1282 = (1'h0);
  reg [(5'h16):(1'h0)] reg1281 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1280 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1275 = (1'h0);
  reg [(3'h7):(1'h0)] reg1273 = (1'h0);
  reg [(5'h15):(1'h0)] reg1270 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1269 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1268 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1267 = (1'h0);
  reg [(3'h4):(1'h0)] reg1266 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1265 = (1'h0);
  reg [(5'h17):(1'h0)] reg1263 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1261 = (1'h0);
  reg [(5'h14):(1'h0)] reg1259 = (1'h0);
  reg [(5'h10):(1'h0)] reg1256 = (1'h0);
  reg [(4'he):(1'h0)] reg1253 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1250 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1249 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1248 = (1'h0);
  reg [(4'h9):(1'h0)] reg1057 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1056 = (1'h0);
  reg [(5'h17):(1'h0)] reg1054 = (1'h0);
  reg [(4'he):(1'h0)] reg1053 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1052 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1050 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1048 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1045 = (1'h0);
  reg [(2'h2):(1'h0)] reg1044 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1043 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1039 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1042 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1039 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1038 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1010 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1035 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1034 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1032 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1029 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1028 = (1'h0);
  reg [(5'h11):(1'h0)] reg1026 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1025 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1024 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1023 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1019 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1018 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1015 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1014 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1013 = (1'h0);
  reg [(4'hb):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1011 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1010 = (1'h0);
  reg [(2'h2):(1'h0)] reg1009 = (1'h0);
  reg [(4'ha):(1'h0)] reg1008 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1007 = (1'h0);
  reg [(2'h2):(1'h0)] reg1006 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1005 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1003 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1002 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1001 = (1'h0);
  reg [(5'h14):(1'h0)] reg1000 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar996 = (1'h0);
  reg [(4'h8):(1'h0)] reg994 = (1'h0);
  reg [(3'h4):(1'h0)] reg992 = (1'h0);
  reg [(5'h15):(1'h0)] reg991 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg987 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg986 = (1'h0);
  reg [(4'h9):(1'h0)] reg984 = (1'h0);
  reg [(3'h7):(1'h0)] forvar983 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg982 = (1'h0);
  reg signed [(4'he):(1'h0)] reg981 = (1'h0);
  reg [(4'h8):(1'h0)] reg979 = (1'h0);
  reg [(2'h3):(1'h0)] reg975 = (1'h0);
  reg [(4'h9):(1'h0)] reg974 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg973 = (1'h0);
  reg [(5'h11):(1'h0)] reg972 = (1'h0);
  reg [(5'h19):(1'h0)] reg969 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg967 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg966 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg965 = (1'h0);
  reg [(5'h15):(1'h0)] reg964 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg962 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg961 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg959 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg958 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar955 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg954 = (1'h0);
  reg [(4'he):(1'h0)] reg953 = (1'h0);
  reg [(5'h1d):(1'h0)] reg952 = (1'h0);
  reg [(5'h12):(1'h0)] reg948 = (1'h0);
  reg [(5'h14):(1'h0)] reg947 = (1'h0);
  reg [(5'h12):(1'h0)] reg946 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg944 = (1'h0);
  reg [(4'hb):(1'h0)] reg943 = (1'h0);
  reg [(5'h12):(1'h0)] reg940 = (1'h0);
  reg [(4'hd):(1'h0)] reg939 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg938 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar937 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg936 = (1'h0);
  reg [(5'h1d):(1'h0)] reg935 = (1'h0);
  reg [(4'ha):(1'h0)] reg934 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg933 = (1'h0);
  reg [(5'h16):(1'h0)] reg931 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg930 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg928 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg927 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg925 = (1'h0);
  reg [(3'h6):(1'h0)] reg924 = (1'h0);
  reg [(3'h6):(1'h0)] reg923 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg922 = (1'h0);
  reg [(4'hf):(1'h0)] reg921 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg920 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar918 = (1'h0);
  reg [(5'h14):(1'h0)] reg917 = (1'h0);
  reg [(5'h1a):(1'h0)] reg915 = (1'h0);
  reg [(5'h19):(1'h0)] reg914 = (1'h0);
  reg [(3'h6):(1'h0)] reg913 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg912 = (1'h0);
  reg [(5'h18):(1'h0)] forvar911 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg908 = (1'h0);
  reg [(3'h6):(1'h0)] reg906 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg904 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar903 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg901 = (1'h0);
  reg [(5'h1f):(1'h0)] reg899 = (1'h0);
  reg [(5'h13):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg893 = (1'h0);
  reg [(4'hc):(1'h0)] reg892 = (1'h0);
  reg [(4'hf):(1'h0)] reg890 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg886 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg882 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg881 = (1'h0);
  reg [(5'h1e):(1'h0)] reg880 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg879 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar875 = (1'h0);
  reg [(4'hd):(1'h0)] reg874 = (1'h0);
  reg [(5'h1b):(1'h0)] reg873 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg871 = (1'h0);
  reg [(5'h13):(1'h0)] forvar869 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar865 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar862 = (1'h0);
  reg [(5'h19):(1'h0)] reg859 = (1'h0);
  reg [(5'h16):(1'h0)] forvar841 = (1'h0);
  reg [(4'he):(1'h0)] reg858 = (1'h0);
  reg [(5'h1a):(1'h0)] reg855 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg853 = (1'h0);
  reg [(4'hd):(1'h0)] reg852 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg851 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar847 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg844 = (1'h0);
  reg [(4'hf):(1'h0)] reg540 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg539 = (1'h0);
  reg [(5'h11):(1'h0)] reg538 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg535 = (1'h0);
  reg [(5'h1b):(1'h0)] reg534 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg531 = (1'h0);
  reg [(4'he):(1'h0)] forvar527 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg525 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg522 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg519 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg518 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg513 = (1'h0);
  reg [(5'h1e):(1'h0)] reg512 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg508 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar507 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg506 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg481 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg501 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg500 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg497 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg496 = (1'h0);
  reg [(4'hd):(1'h0)] reg494 = (1'h0);
  reg [(5'h1c):(1'h0)] reg493 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar490 = (1'h0);
  reg [(4'hf):(1'h0)] reg488 = (1'h0);
  reg [(5'h1c):(1'h0)] reg486 = (1'h0);
  reg [(5'h1f):(1'h0)] reg483 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar481 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg475 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg474 = (1'h0);
  reg [(5'h10):(1'h0)] reg472 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg462 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg460 = (1'h0);
  reg [(4'ha):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar458 = (1'h0);
  reg signed [(4'he):(1'h0)] reg455 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg454 = (1'h0);
  reg [(5'h16):(1'h0)] reg451 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg450 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg447 = (1'h0);
  reg [(3'h6):(1'h0)] forvar445 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar440 = (1'h0);
  assign y = {wire1993,
                 wire1992,
                 wire1990,
                 wire1478,
                 wire1247,
                 wire1246,
                 wire1244,
                 wire1059,
                 wire860,
                 wire838,
                 wire542,
                 reg1994,
                 reg1386,
                 reg1381,
                 reg1380,
                 reg1353,
                 reg1378,
                 reg1377,
                 reg1374,
                 reg1372,
                 reg1369,
                 reg1368,
                 reg1366,
                 reg1362,
                 reg1361,
                 reg1360,
                 reg1356,
                 reg1355,
                 reg1354,
                 reg1352,
                 reg1350,
                 reg1346,
                 reg1345,
                 reg1344,
                 reg1341,
                 reg1339,
                 reg1337,
                 reg1335,
                 reg1334,
                 reg1331,
                 reg1330,
                 reg1327,
                 reg1323,
                 reg1322,
                 reg1320,
                 reg1319,
                 reg1317,
                 reg1313,
                 reg1312,
                 reg1310,
                 reg1308,
                 reg1307,
                 reg1306,
                 reg1302,
                 reg1301,
                 reg1299,
                 reg1295,
                 reg1294,
                 reg1292,
                 reg1290,
                 reg1285,
                 reg1283,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1274,
                 reg1272,
                 reg1271,
                 reg1264,
                 reg1262,
                 reg1260,
                 reg1258,
                 reg1257,
                 reg1255,
                 reg1254,
                 reg1252,
                 reg1251,
                 reg1058,
                 reg1055,
                 reg1051,
                 reg1049,
                 reg1047,
                 reg1046,
                 reg1041,
                 reg1040,
                 reg1011,
                 reg1037,
                 reg1036,
                 reg1033,
                 reg1031,
                 reg1030,
                 reg1027,
                 reg1022,
                 reg1021,
                 reg1020,
                 reg1017,
                 reg1016,
                 reg1004,
                 reg999,
                 reg998,
                 reg997,
                 reg996,
                 reg995,
                 reg993,
                 reg990,
                 reg989,
                 reg988,
                 reg985,
                 reg980,
                 reg978,
                 reg977,
                 reg976,
                 reg971,
                 reg970,
                 reg968,
                 reg963,
                 reg960,
                 reg957,
                 reg956,
                 reg951,
                 reg950,
                 reg949,
                 reg945,
                 reg942,
                 reg941,
                 reg932,
                 reg929,
                 reg926,
                 reg919,
                 reg916,
                 reg910,
                 reg909,
                 reg907,
                 reg905,
                 reg902,
                 reg900,
                 reg898,
                 reg897,
                 reg895,
                 reg894,
                 reg891,
                 reg889,
                 reg888,
                 reg887,
                 reg885,
                 reg884,
                 reg883,
                 reg878,
                 reg877,
                 reg876,
                 reg872,
                 reg870,
                 reg868,
                 reg867,
                 reg866,
                 reg864,
                 reg863,
                 reg861,
                 reg847,
                 reg857,
                 reg856,
                 reg854,
                 reg850,
                 reg849,
                 reg848,
                 reg845,
                 reg843,
                 reg842,
                 reg841,
                 reg840,
                 reg541,
                 reg537,
                 reg536,
                 reg533,
                 reg532,
                 reg530,
                 reg529,
                 reg528,
                 reg524,
                 reg523,
                 reg507,
                 reg521,
                 reg520,
                 reg517,
                 reg516,
                 reg514,
                 reg511,
                 reg510,
                 reg509,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg498,
                 reg495,
                 reg492,
                 reg491,
                 reg489,
                 reg487,
                 reg485,
                 reg484,
                 reg482,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 reg473,
                 reg471,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg461,
                 reg457,
                 reg456,
                 reg453,
                 reg452,
                 reg449,
                 reg448,
                 reg446,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 reg1385,
                 forvar1384,
                 reg1383,
                 reg1382,
                 reg1371,
                 reg1363,
                 reg1358,
                 reg1379,
                 reg1376,
                 reg1375,
                 reg1373,
                 forvar1371,
                 reg1370,
                 reg1367,
                 reg1365,
                 reg1364,
                 forvar1363,
                 reg1359,
                 forvar1358,
                 reg1357,
                 forvar1353,
                 reg1351,
                 reg1349,
                 reg1348,
                 reg1347,
                 forvar1343,
                 reg1342,
                 reg1340,
                 reg1338,
                 forvar1336,
                 reg1333,
                 reg1332,
                 reg1329,
                 forvar1328,
                 reg1328,
                 reg1326,
                 reg1325,
                 reg1324,
                 forvar1321,
                 reg1318,
                 reg1316,
                 reg1315,
                 reg1314,
                 forvar1311,
                 reg1309,
                 forvar1305,
                 reg1304,
                 reg1303,
                 reg1300,
                 reg1298,
                 reg1297,
                 reg1296,
                 reg1293,
                 reg1291,
                 reg1289,
                 reg1288,
                 forvar1287,
                 reg1286,
                 reg1284,
                 reg1282,
                 reg1281,
                 reg1280,
                 forvar1275,
                 reg1273,
                 reg1270,
                 forvar1269,
                 reg1268,
                 forvar1267,
                 reg1266,
                 reg1265,
                 reg1263,
                 reg1261,
                 reg1259,
                 reg1256,
                 reg1253,
                 forvar1250,
                 forvar1249,
                 reg1248,
                 reg1057,
                 reg1056,
                 reg1054,
                 reg1053,
                 reg1052,
                 reg1050,
                 reg1048,
                 reg1045,
                 reg1044,
                 reg1043,
                 forvar1039,
                 reg1042,
                 reg1039,
                 reg1038,
                 forvar1010,
                 forvar1035,
                 reg1034,
                 reg1032,
                 reg1029,
                 reg1028,
                 reg1026,
                 reg1025,
                 reg1024,
                 reg1023,
                 reg1019,
                 forvar1018,
                 reg1015,
                 reg1014,
                 reg1013,
                 reg1012,
                 forvar1011,
                 reg1010,
                 reg1009,
                 reg1008,
                 reg1007,
                 reg1006,
                 reg1005,
                 reg1003,
                 reg1002,
                 forvar1001,
                 reg1000,
                 forvar996,
                 reg994,
                 reg992,
                 reg991,
                 reg987,
                 reg986,
                 reg984,
                 forvar983,
                 reg982,
                 reg981,
                 reg979,
                 reg975,
                 reg974,
                 reg973,
                 reg972,
                 reg969,
                 reg967,
                 reg966,
                 reg965,
                 reg964,
                 reg962,
                 reg961,
                 reg959,
                 reg958,
                 forvar955,
                 reg954,
                 reg953,
                 reg952,
                 reg948,
                 reg947,
                 reg946,
                 reg944,
                 reg943,
                 reg940,
                 reg939,
                 reg938,
                 forvar937,
                 reg936,
                 reg935,
                 reg934,
                 reg933,
                 reg931,
                 reg930,
                 reg928,
                 reg927,
                 reg925,
                 reg924,
                 reg923,
                 reg922,
                 reg921,
                 reg920,
                 forvar918,
                 reg917,
                 reg915,
                 reg914,
                 reg913,
                 reg912,
                 forvar911,
                 reg908,
                 reg906,
                 reg904,
                 forvar903,
                 reg901,
                 reg899,
                 reg896,
                 reg893,
                 reg892,
                 reg890,
                 reg886,
                 reg882,
                 reg881,
                 reg880,
                 reg879,
                 forvar875,
                 reg874,
                 reg873,
                 reg871,
                 forvar869,
                 forvar865,
                 forvar862,
                 reg859,
                 forvar841,
                 reg858,
                 reg855,
                 reg853,
                 reg852,
                 reg851,
                 forvar847,
                 reg846,
                 reg844,
                 reg540,
                 reg539,
                 reg538,
                 reg535,
                 reg534,
                 reg531,
                 forvar527,
                 reg526,
                 reg525,
                 reg522,
                 reg519,
                 reg518,
                 reg515,
                 reg513,
                 reg512,
                 reg508,
                 forvar507,
                 reg506,
                 reg481,
                 reg501,
                 reg500,
                 reg499,
                 reg497,
                 reg496,
                 reg494,
                 reg493,
                 forvar490,
                 reg488,
                 reg486,
                 reg483,
                 forvar481,
                 reg475,
                 reg474,
                 reg472,
                 reg462,
                 reg460,
                 reg459,
                 forvar458,
                 reg455,
                 reg454,
                 reg451,
                 reg450,
                 reg447,
                 forvar445,
                 forvar440,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar440 = (1'h0); (forvar440 < (3'h4)); forvar440 = (forvar440 + (1'h1)))
        begin
          if ((8'hb7))
            begin
              reg441 <= wire436;
              reg442 <= $unsigned((wire439[(2'h3):(1'h1)] ?
                  $signed((&(wire435 ?
                      wire436 : (7'h56)))) : {(reg441[(4'hb):(4'h9)] >>> (^wire436)),
                      reg441[(4'ha):(1'h1)]}));
              reg443 <= forvar440[(5'h13):(4'he)];
              reg444 <= $unsigned(((($signed(wire439) ?
                      wire437[(3'h5):(2'h2)] : reg442) != $signed(wire437[(5'h13):(3'h7)])) ?
                  $unsigned((^reg442)) : {(reg442 * $signed(wire435))}));
            end
          else
            begin
              reg441 <= {reg442[(3'h7):(3'h7)], $unsigned((7'h4a))};
              reg442 <= (~$signed(wire437));
            end
          for (forvar445 = (1'h0); (forvar445 < (2'h3)); forvar445 = (forvar445 + (1'h1)))
            begin
              reg446 <= (~&$signed((!$signed($unsigned(wire438)))));
              reg447 = (7'h45);
              reg448 <= ($unsigned((-(forvar445 != reg447))) || $unsigned($signed(wire436[(3'h7):(3'h7)])));
              reg449 <= $signed($signed({((reg448 == (8'ha6)) > (wire436 < wire437)),
                  (~|(~reg447))}));
              reg450 = (((|($signed((7'h47)) ?
                          reg441 : reg441[(1'h0):(1'h0)])) ?
                      (|{(reg448 ? reg448 : reg448),
                          (~|reg441),
                          (reg443 ? wire438 : wire437)}) : forvar445) ?
                  ($unsigned({{reg443, reg441},
                          $unsigned(reg443),
                          $signed(wire435)}) ?
                      reg449[(4'hc):(3'h5)] : ((+((7'h41) + reg444)) ?
                          (forvar440[(4'h8):(2'h3)] ?
                              ((7'h4b) >>> reg441) : wire439[(4'hd):(3'h4)]) : reg443)) : $signed(({(reg443 ~^ reg442),
                      {wire439}} != (reg443 ?
                      (reg447 ? wire437 : reg449) : $unsigned(reg449)))));
              reg451 = reg442;
            end
          if (({(+(&$signed(forvar440))), wire439} ? (^wire438) : (+reg446)))
            begin
              reg452 <= $signed(reg444[(1'h0):(1'h0)]);
            end
          else
            begin
              reg452 <= $signed(reg442);
              reg453 <= {$unsigned(reg444[(3'h4):(1'h1)]),
                  {{$unsigned(reg448[(4'he):(4'hb)]),
                          $signed((reg448 ? reg443 : wire438)),
                          $signed((forvar440 ? reg441 : reg441))}},
                  ($signed(((+forvar440) ?
                      (wire435 ?
                          forvar445 : wire435) : $signed(reg448))) << reg444[(1'h0):(1'h0)])};
              reg454 = $signed((8'hb5));
              reg455 = $signed($signed((((reg444 < (7'h52)) ?
                  reg443[(4'h8):(2'h2)] : $unsigned(reg441)) > ((reg443 ?
                      (7'h4a) : reg447) ?
                  (8'h9d) : wire438[(3'h4):(2'h2)]))));
              reg456 <= $signed($unsigned((^~{$unsigned(reg452), reg444})));
              reg457 <= $signed($unsigned({reg442[(5'h1a):(2'h2)],
                  reg451,
                  ($unsigned(reg448) || $unsigned(reg450))}));
            end
          for (forvar458 = (1'h0); (forvar458 < (2'h2)); forvar458 = (forvar458 + (1'h1)))
            begin
              reg459 = (wire438 ?
                  $unsigned($unsigned($unsigned({reg449,
                      reg441,
                      (7'h4b)}))) : ((~^wire436) >> reg454[(1'h1):(1'h1)]));
              reg460 = (~^$signed(reg450));
              reg461 <= ($signed(($signed(wire439[(4'he):(4'hc)]) ~^ $signed(reg447))) ?
                  reg443 : {forvar445, $signed({(reg446 ? (8'ha4) : reg444)})});
              reg462 = ($unsigned((wire438[(4'hf):(4'hc)] ?
                  ((~^reg446) ?
                      $signed(reg447) : (reg449 ?
                          reg443 : reg447)) : (~^$signed((8'hb8))))) <<< forvar458);
              reg463 <= reg444;
              reg464 <= (wire439[(4'he):(3'h6)] ?
                  (~^$signed((reg443[(3'h7):(2'h3)] ?
                      ((8'hbd) ?
                          reg448 : reg460) : (!reg451)))) : wire436[(2'h2):(2'h2)]);
            end
          reg465 <= wire439[(3'h4):(2'h2)];
          if (((reg464[(5'h17):(4'hf)] ?
              {$signed(reg452),
                  (reg463[(5'h1d):(3'h7)] ?
                      reg454 : (reg450 ?
                          reg459 : reg452))} : $unsigned(reg464)) * $signed((((reg447 ?
                      (8'ha3) : reg463) ?
                  reg459[(4'ha):(3'h4)] : (reg464 ? reg447 : reg453)) ?
              $unsigned(reg459) : ($unsigned(reg457) == reg444)))))
            begin
              reg466 <= ($signed((reg442 ?
                      {reg459} : (reg446[(1'h1):(1'h0)] >= (reg460 == reg456)))) ?
                  $unsigned($unsigned($signed((reg443 ?
                      reg459 : reg462)))) : {reg451,
                      ((reg454 >= (forvar458 ? (7'h52) : (8'hb6))) ?
                          {reg449} : reg462[(4'ha):(4'h8)])});
              reg467 <= ((^($signed(reg453[(5'h15):(5'h14)]) ?
                  reg456 : {(&(8'hbe))})) >>> reg461);
              reg468 <= ($unsigned($unsigned({reg455[(3'h7):(3'h5)],
                      reg449[(3'h5):(2'h2)]})) ?
                  ($signed((&(reg441 <= wire439))) ?
                      $unsigned($unsigned($signed(reg457))) : reg462) : (-($unsigned($signed((8'hba))) ?
                      (reg447 ?
                          reg464[(4'hd):(3'h6)] : $unsigned(reg448)) : {((8'ha8) ~^ (7'h40)),
                          $unsigned(reg464),
                          reg447})));
              reg469 <= ((-$signed((^~((8'hbd) && (7'h4d))))) ?
                  (&reg462) : $signed((reg456 && $signed((~&(8'hb7))))));
              reg470 <= ($unsigned({$unsigned((~&reg441)),
                  ((reg450 ? (8'hb6) : (7'h41)) || {reg450}),
                  reg457[(4'h9):(4'h8)]}) + {$unsigned(((reg441 >>> (7'h52)) ^~ $signed(reg448)))});
              reg471 <= (({reg444} && {reg450[(2'h3):(2'h2)]}) && (~(|((8'h9e) & reg470))));
              reg472 = (&$unsigned((~|wire439)));
            end
          else
            begin
              reg472 = ((8'hb1) ?
                  (reg456[(3'h7):(2'h2)] << (((reg451 && reg455) + $signed(wire438)) | (wire438 >>> reg459[(3'h7):(3'h4)]))) : (((+((8'ha9) ?
                      reg452 : wire436)) || (8'ha1)) == $signed($unsigned((reg468 ?
                      (8'ha4) : reg451)))));
              reg473 <= reg447[(1'h1):(1'h0)];
              reg474 = {reg466};
              reg475 = {reg469};
              reg476 <= $unsigned($unsigned((8'hb9)));
              reg477 <= (&$unsigned(($signed((~^reg465)) ?
                  {(wire435 ? (7'h46) : reg449)} : ($signed(reg463) >= (reg450 ?
                      reg456 : reg441)))));
            end
        end
      reg478 <= reg456[(4'ha):(2'h3)];
      reg479 <= (wire435[(1'h1):(1'h1)] ?
          reg456[(5'h10):(3'h4)] : (~^reg465[(1'h0):(1'h0)]));
      if ($signed((!$signed(((reg443 == reg460) ?
          wire438[(4'hc):(4'h9)] : (reg478 ? reg464 : (7'h44)))))))
        begin
          reg480 <= $unsigned(($signed(wire436) != ((~^$unsigned(reg452)) ?
              (+wire439) : forvar445[(3'h6):(2'h3)])));
          for (forvar481 = (1'h0); (forvar481 < (3'h6)); forvar481 = (forvar481 + (1'h1)))
            begin
              reg482 <= (+{forvar445});
            end
          if ({($unsigned(reg453) && (+reg457[(1'h1):(1'h1)])),
              $signed({reg478})})
            begin
              reg483 = reg456;
              reg484 <= $signed($unsigned((wire436[(3'h5):(3'h5)] ?
                  reg472 : reg469)));
              reg485 <= (-$unsigned({((!reg451) <<< (~|reg471)),
                  {reg470[(3'h6):(2'h2)], reg459, $signed(reg469)},
                  $signed((^reg451))}));
              reg486 = (reg467[(1'h0):(1'h0)] >> (($signed(reg456[(2'h3):(2'h2)]) ?
                  (+{reg457}) : ($unsigned(reg468) ?
                      (reg482 > reg473) : (reg474 ?
                          reg479 : reg449))) > $signed((^~((8'hb9) ~^ (8'haf))))));
              reg487 <= ($signed(reg469[(1'h1):(1'h0)]) > wire435);
            end
          else
            begin
              reg483 = {$signed(wire436[(3'h4):(1'h1)])};
              reg484 <= reg468;
            end
          reg488 = ($unsigned($unsigned((~|reg462))) == (|$signed((~$unsigned(reg452)))));
          reg489 <= (~($unsigned($signed(reg442[(5'h1b):(3'h5)])) == (reg450 | ((reg474 ?
              reg443 : reg446) & $unsigned(reg453)))));
          for (forvar490 = (1'h0); (forvar490 < (1'h0)); forvar490 = (forvar490 + (1'h1)))
            begin
              reg491 <= $unsigned(($unsigned($signed({(8'ha9)})) < forvar481));
              reg492 <= $unsigned((~&{(reg491 ~^ (-reg444)),
                  reg476[(3'h6):(2'h2)],
                  reg446}));
              reg493 = (~^$signed(($signed($unsigned(reg483)) != (!(8'ha6)))));
              reg494 = forvar445;
              reg495 <= reg466[(1'h1):(1'h0)];
              reg496 = (~reg451);
            end
          if (reg470[(3'h7):(3'h7)])
            begin
              reg497 = ({$signed((^~reg465[(1'h0):(1'h0)]))} ?
                  ({(~|(reg448 | reg453)),
                      $signed((reg443 ? reg463 : reg450)),
                      ($signed(reg484) ?
                          (reg495 || (8'ha9)) : (8'hbd))} <<< $unsigned($unsigned((~&(7'h56))))) : ((reg444[(1'h0):(1'h0)] > (&((8'ha9) ~^ wire435))) ?
                      $signed(((reg468 ?
                          reg461 : reg447) == $unsigned(reg441))) : reg471));
            end
          else
            begin
              reg498 <= reg495;
              reg499 = (({reg455,
                      ($signed((8'hbf)) ?
                          (reg492 ?
                              reg474 : reg444) : (forvar481 >> (7'h49)))} ?
                  {reg450,
                      $signed((reg484 ? (8'hab) : wire436)),
                      (~|(8'hb4))} : {$signed((~^reg469)),
                      ($signed(reg483) ?
                          (|reg482) : (reg469 ?
                              reg457 : (7'h4f)))}) | (reg492[(3'h4):(2'h3)] < reg482));
              reg500 = (~reg441);
              reg501 = (&(({$signed((8'hbb)),
                      (reg467 ? reg488 : (8'hb3)),
                      reg455[(2'h3):(1'h0)]} ?
                  ($signed((7'h4f)) ?
                      (7'h4b) : $signed((7'h46))) : $unsigned($unsigned(reg469))) >> reg456[(4'h8):(1'h1)]));
              reg502 <= ((~&{$unsigned((reg501 ? reg498 : reg482))}) & reg480);
              reg503 <= ($signed({$unsigned($unsigned(reg465))}) | (wire435[(1'h1):(1'h0)] ~^ $signed($unsigned(reg480))));
            end
        end
      else
        begin
          reg481 = ($signed({(^~(!forvar440)),
              ((reg482 ^~ reg476) ? (^~reg468) : (8'hb4)),
              {reg476[(3'h6):(3'h5)],
                  {reg477, reg464}}}) | (&$unsigned(reg444)));
        end
      reg504 <= reg488;
      reg505 <= $signed({($unsigned($unsigned(reg472)) ^ $unsigned((reg489 >= reg455)))});
    end
  always
    @(posedge clk) begin
      reg506 = reg471;
      if (((7'h4c) != ((!reg482) ?
          $unsigned({(~^reg487),
              {reg456,
                  wire437,
                  reg467}}) : $signed(((reg466 == reg467) >> (!reg479))))))
        begin
          for (forvar507 = (1'h0); (forvar507 < (3'h5)); forvar507 = (forvar507 + (1'h1)))
            begin
              reg508 = ((reg470[(4'h8):(3'h6)] ?
                      $signed($unsigned($signed(reg442))) : (-$unsigned(reg441))) ?
                  wire437[(3'h5):(1'h1)] : $signed((~^($unsigned(reg465) > reg473[(4'he):(4'h8)]))));
              reg509 <= {$unsigned((!reg470)),
                  reg503,
                  ({$unsigned($unsigned(wire437))} ^ reg480)};
              reg510 <= $signed($signed((8'hbd)));
              reg511 <= ((wire435 ?
                      $signed($unsigned(reg498[(1'h1):(1'h1)])) : ((!reg466) ^~ reg480)) ?
                  $signed($unsigned(($unsigned(reg477) ?
                      $unsigned(reg444) : reg456))) : reg504[(4'hb):(1'h1)]);
              reg512 = ($unsigned((($signed(reg508) != (reg469 == reg446)) || ($unsigned(reg502) ?
                      {reg489, reg511} : {reg484, wire438, wire436}))) ?
                  $unsigned($signed((reg484[(3'h5):(3'h5)] != reg468[(3'h4):(1'h1)]))) : ((~&{(wire435 ^~ reg466),
                      $unsigned(reg446)}) + ((~&$signed((8'hab))) ^ {$signed(reg446),
                      (-reg495)})));
              reg513 = (|reg489);
              reg514 <= {(reg492[(2'h3):(2'h3)] == (reg471 < reg491[(4'he):(1'h0)])),
                  (reg446[(4'he):(1'h1)] ?
                      (-(&{reg449,
                          reg505,
                          reg452})) : $signed(reg477[(3'h7):(1'h1)]))};
            end
          if ((^reg456))
            begin
              reg515 = $signed({(forvar507 ?
                      {wire439,
                          reg487[(4'hf):(1'h1)],
                          $unsigned((7'h53))} : (|((7'h41) >>> reg457))),
                  $signed((reg476[(3'h6):(3'h6)] & (reg509 ?
                      (7'h54) : reg489))),
                  reg461[(5'h11):(2'h2)]});
              reg516 <= reg464;
              reg517 <= forvar507;
              reg518 = $unsigned(reg487[(4'hf):(1'h0)]);
              reg519 = ((reg471[(1'h1):(1'h1)] >>> $unsigned((^(reg477 * reg461)))) * $unsigned($unsigned(({reg470} ?
                  (&reg495) : {reg514, reg473, reg468}))));
            end
          else
            begin
              reg515 = (+reg515[(4'hb):(2'h3)]);
            end
          reg520 <= {$unsigned({((7'h4d) ?
                      $unsigned(reg480) : (wire438 ? wire435 : (8'hb7)))})};
          reg521 <= $signed({(+(reg518 ? (reg515 >> (7'h49)) : {wire436})),
              $unsigned({(^~reg508)})});
          reg522 = $signed((~|$unsigned(((^~wire437) ^ $unsigned(reg495)))));
        end
      else
        begin
          reg507 <= $unsigned($unsigned($signed($unsigned(reg449[(4'hb):(4'hb)]))));
        end
      reg523 <= $signed((&$signed((7'h4f))));
      reg524 <= ((reg446 ? (7'h4f) : (~$unsigned(reg463[(5'h1d):(5'h1d)]))) ?
          (+(^~(reg442 >>> (&reg515)))) : $signed($signed(reg479)));
      if ({reg471[(3'h4):(3'h4)],
          ((((reg495 >= reg495) ? reg470 : ((7'h49) > wire435)) == (((8'haa) ?
                  reg442 : reg487) ?
              (!reg480) : (reg478 ?
                  reg469 : reg476))) ~^ $unsigned(((~^reg504) && $signed(reg478))))})
        begin
          reg525 = (reg448[(4'h8):(2'h3)] ~^ $signed($signed((8'hbe))));
        end
      else
        begin
          reg525 = reg506;
          reg526 = reg461[(1'h0):(1'h0)];
          for (forvar527 = (1'h0); (forvar527 < (2'h3)); forvar527 = (forvar527 + (1'h1)))
            begin
              reg528 <= reg463;
              reg529 <= $unsigned((reg492[(2'h3):(2'h2)] || (+reg498[(4'h9):(4'h9)])));
              reg530 <= reg467[(1'h1):(1'h1)];
              reg531 = $signed((|reg463));
              reg532 <= reg506[(3'h4):(1'h1)];
              reg533 <= reg446[(4'hd):(4'hc)];
              reg534 = reg531;
            end
          reg535 = $signed(($unsigned(({reg516,
              (8'hb6),
              reg487} * reg495)) | (reg514 ?
              $signed($unsigned((7'h4e))) : (+(reg468 == reg525)))));
          reg536 <= {$signed(reg470)};
        end
      if (reg489[(2'h3):(1'h1)])
        begin
          if ({reg456})
            begin
              reg537 <= $signed((-(~|(!(reg452 && reg513)))));
              reg538 = (wire437[(5'h10):(3'h4)] ?
                  reg471 : $unsigned((reg467 * $unsigned((reg452 * reg489)))));
            end
          else
            begin
              reg538 = reg482[(1'h1):(1'h0)];
              reg539 = ({({reg498[(3'h5):(1'h1)]} <<< $signed($unsigned(reg509))),
                      (|reg514[(2'h2):(1'h0)])} ?
                  $unsigned(reg506) : reg538);
              reg540 = reg528[(1'h0):(1'h0)];
            end
          reg541 <= (reg478 ?
              reg519 : $signed($unsigned($unsigned((~reg480)))));
        end
      else
        begin
          reg538 = (reg540 ?
              reg464[(5'h13):(4'hb)] : (^~$signed($unsigned((reg477 ?
                  (8'hb6) : reg524)))));
        end
    end
  assign wire542 = ((reg536[(4'h9):(3'h6)] ?
                       (|{(~|reg468),
                           (reg480 ? reg529 : reg452)}) : $signed(((reg477 ?
                           reg491 : reg477) < (reg530 | reg468)))) <<< (~^reg479[(3'h4):(1'h0)]));
  module543 #() modinst839 (wire838, clk, reg485, reg442, reg498, reg479);
  always
    @(posedge clk) begin
      reg840 <= $signed(wire542[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      if ({(({reg485[(3'h7):(3'h5)],
                  reg514,
                  $signed(reg482)} && reg524[(1'h0):(1'h0)]) ?
              ($unsigned(reg498[(3'h5):(3'h4)]) >> $unsigned($signed((8'hb7)))) : ($signed(((8'hac) ?
                  reg476 : reg529)) <= ($signed(reg478) != (reg528 ?
                  reg446 : reg510)))),
          reg523,
          (reg517 <= $unsigned(reg469[(2'h3):(1'h1)]))})
        begin
          if ($signed($unsigned((~&({reg479, reg533} <<< $signed(reg524))))))
            begin
              reg841 <= $unsigned({((&((7'h49) * reg491)) > $unsigned((~^reg469))),
                  (+$unsigned($unsigned(reg491))),
                  (($signed(reg480) ?
                      $unsigned(reg463) : $unsigned(reg484)) >> $unsigned((|reg840)))});
              reg842 <= $unsigned((reg476[(2'h3):(2'h2)] ?
                  {{$signed(reg523),
                          $signed(reg491)}} : wire435[(1'h1):(1'h0)]));
              reg843 <= (reg491[(3'h4):(3'h4)] > (reg461[(4'h8):(2'h3)] - (^~reg489[(5'h13):(3'h7)])));
              reg844 = (^(reg484[(3'h6):(1'h1)] ?
                  ((|$signed(reg448)) ?
                      (reg523[(4'he):(1'h1)] ?
                          $signed(reg537) : $signed((7'h55))) : (&(~|wire435))) : (-$unsigned($unsigned(reg502)))));
              reg845 <= ($signed(reg502) || ($signed(wire438) ?
                  $unsigned(($signed(reg479) ?
                      $unsigned(reg449) : (~^reg484))) : $signed(reg470[(4'h8):(1'h0)])));
              reg846 = (+(reg461 >> (^~$signed((~|reg502)))));
            end
          else
            begin
              reg841 <= {reg533[(5'h14):(2'h3)],
                  $signed(reg492[(2'h2):(2'h2)])};
              reg842 <= ({$unsigned((~(reg465 ?
                      reg530 : reg845)))} & ((~(reg478 & $signed(reg530))) > reg495));
            end
          for (forvar847 = (1'h0); (forvar847 < (2'h3)); forvar847 = (forvar847 + (1'h1)))
            begin
              reg848 <= wire438;
              reg849 <= ((|reg524) ?
                  (~&((wire437[(5'h14):(5'h12)] >>> reg537) ?
                      (reg840 ^~ reg470) : (reg524 ?
                          {reg484,
                              reg444} : reg482))) : $unsigned($signed((~|reg449[(3'h5):(2'h2)]))));
            end
          if (reg502)
            begin
              reg850 <= $signed(reg485[(3'h7):(1'h1)]);
              reg851 = (~|reg840);
              reg852 = (^~$signed((7'h42)));
            end
          else
            begin
              reg851 = reg468;
              reg852 = {$unsigned($unsigned(({reg467} ?
                      (reg479 ? (7'h51) : (8'hb2)) : $signed((8'hb9)))))};
              reg853 = reg846[(5'h19):(5'h15)];
            end
          if ((7'h43))
            begin
              reg854 <= ((reg502[(3'h7):(3'h5)] && ($signed($unsigned(reg502)) ^~ (reg452 ?
                      $signed(reg504) : {reg507}))) ?
                  ($signed(((~&reg504) ?
                      $unsigned(reg843) : reg840)) + (~^((reg514 ^~ reg480) ?
                      reg463 : $signed(reg845)))) : $signed((^~wire435)));
              reg855 = reg529;
              reg856 <= reg464;
            end
          else
            begin
              reg854 <= ($signed($signed((reg510 ^~ $signed(reg473)))) && reg444[(1'h1):(1'h0)]);
              reg856 <= $signed($unsigned((($signed(reg533) << $signed(reg478)) ?
                  $unsigned((wire438 ? reg840 : reg509)) : (reg503 ?
                      reg530[(5'h12):(3'h4)] : (reg529 ? reg446 : reg489)))));
              reg857 <= (-$unsigned((7'h47)));
            end
          reg858 = $signed(((((reg441 | wire438) ?
              (reg841 ?
                  (7'h4a) : reg851) : $unsigned(wire542)) >>> reg491[(4'he):(1'h1)]) || $unsigned((&reg449[(2'h3):(1'h1)]))));
        end
      else
        begin
          for (forvar841 = (1'h0); (forvar841 < (1'h0)); forvar841 = (forvar841 + (1'h1)))
            begin
              reg842 <= reg516;
              reg844 = reg457[(3'h4):(2'h3)];
              reg846 = (~$signed((reg479 - $signed((reg441 ?
                  reg840 : reg468)))));
            end
          reg847 <= (^~(~&$signed(reg441[(4'he):(1'h1)])));
          reg848 <= $signed($signed(({(^~reg842)} > (reg521 >> reg532[(5'h18):(5'h11)]))));
        end
      reg859 = (reg532 ?
          {(wire436[(4'h9):(3'h6)] ?
                  {wire435[(2'h3):(2'h2)]} : ((!reg855) ?
                      $signed(reg448) : wire435))} : reg473[(1'h0):(1'h0)]);
    end
  assign wire860 = $signed(((8'haa) ?
                       reg854 : $signed((!(wire438 >= reg476)))));
  always
    @(posedge clk) begin
      reg861 <= {wire439};
      for (forvar862 = (1'h0); (forvar862 < (1'h0)); forvar862 = (forvar862 + (1'h1)))
        begin
          reg863 <= ($unsigned((8'ha6)) ?
              $unsigned(reg457) : reg457[(2'h2):(2'h2)]);
          reg864 <= $signed($unsigned(reg511[(2'h2):(2'h2)]));
          for (forvar865 = (1'h0); (forvar865 < (3'h5)); forvar865 = (forvar865 + (1'h1)))
            begin
              reg866 <= reg505;
              reg867 <= {({(|reg520),
                          $unsigned((+reg441)),
                          reg465[(4'ha):(3'h6)]} ?
                      (^~$unsigned((^reg863))) : (reg866[(4'ha):(3'h7)] ?
                          $signed((reg856 * reg502)) : {(^reg524)}))};
            end
          reg868 <= (^(((~forvar862) ?
                  ($unsigned(reg533) ?
                      $unsigned((8'hae)) : {reg511,
                          (8'hbb),
                          reg467}) : ((reg843 ? reg523 : (8'h9c)) ?
                      $unsigned(wire860) : ((7'h42) ? reg470 : reg453))) ?
              {(8'hac), (~&$signed(reg476))} : reg867));
          for (forvar869 = (1'h0); (forvar869 < (3'h5)); forvar869 = (forvar869 + (1'h1)))
            begin
              reg870 <= $signed(reg456[(2'h2):(1'h1)]);
              reg871 = $signed({$signed($signed({reg541, reg485, reg448})),
                  {($unsigned(reg449) ? {(7'h57), reg868} : $signed(reg511)),
                      ($signed(reg466) * (forvar862 || reg487)),
                      $signed((reg480 < reg478))},
                  (($unsigned(reg870) ?
                      wire838[(3'h6):(3'h4)] : (reg476 ?
                          reg536 : reg521)) == ($unsigned((7'h46)) & reg463[(2'h3):(2'h2)]))});
              reg872 <= $signed(reg485[(3'h6):(2'h2)]);
              reg873 = ((&(!((-reg505) == reg511[(4'h9):(3'h5)]))) == reg861);
              reg874 = ($unsigned($unsigned($signed(((8'hac) ?
                  reg469 : reg482)))) | reg848[(1'h0):(1'h0)]);
            end
          for (forvar875 = (1'h0); (forvar875 < (2'h3)); forvar875 = (forvar875 + (1'h1)))
            begin
              reg876 <= reg532[(5'h10):(3'h5)];
              reg877 <= wire838[(4'hb):(1'h1)];
              reg878 <= reg441[(4'hf):(3'h5)];
              reg879 = (((((&reg444) | ((8'haf) == (8'hbc))) ?
                      reg842[(1'h1):(1'h0)] : ((forvar862 == reg850) ?
                          (reg504 ? reg470 : reg489) : (reg509 ?
                              reg842 : reg541))) || (^($unsigned(reg840) - $signed(reg466)))) ?
                  $signed(forvar862[(3'h4):(1'h1)]) : ($unsigned($signed(reg507[(3'h5):(2'h2)])) ?
                      $unsigned($signed(reg448[(1'h1):(1'h0)])) : $unsigned((reg504[(4'hc):(1'h1)] ?
                          (|(7'h40)) : $signed(reg854)))));
            end
        end
      reg880 = reg863[(5'h10):(1'h1)];
    end
  always
    @(posedge clk) begin
      if (({$signed((^{reg850})),
              ({reg845[(4'hd):(4'hb)]} ?
                  ($unsigned((7'h4f)) ? {(8'had)} : (!reg850)) : (7'h44))} ?
          $signed(reg456) : (^((7'h49) && reg843[(3'h4):(2'h2)]))))
        begin
          reg881 = ($unsigned((+reg840)) ?
              $unsigned(reg478[(2'h2):(2'h2)]) : $unsigned((({reg452,
                      wire439} || $signed(reg876)) ?
                  $signed((!reg480)) : reg466[(4'hb):(3'h7)])));
          reg882 = reg453[(3'h4):(1'h0)];
          if ((+reg876))
            begin
              reg883 <= reg509;
              reg884 <= $signed(reg457[(2'h3):(1'h0)]);
              reg885 <= {$signed($unsigned(($unsigned((7'h4f)) ?
                      (7'h40) : $signed(reg449))))};
              reg886 = $unsigned((8'h9e));
              reg887 <= ($unsigned((7'h43)) ?
                  {{($unsigned(reg505) ? $unsigned(reg867) : (7'h41)),
                          $signed((reg842 <<< reg528)),
                          reg530[(5'h14):(4'h8)]},
                      ($unsigned($unsigned(wire542)) > reg446[(4'hc):(2'h2)]),
                      $signed($unsigned($unsigned(reg536)))} : (^~$signed(reg464[(3'h4):(2'h3)])));
              reg888 <= {$signed(reg536[(5'h18):(5'h18)]),
                  $unsigned(($unsigned($unsigned(reg491)) == $unsigned(reg503[(3'h7):(3'h4)]))),
                  reg848};
              reg889 <= reg478[(3'h6):(3'h6)];
            end
          else
            begin
              reg883 <= (wire439 <= reg503[(4'ha):(4'h8)]);
              reg886 = (7'h47);
              reg890 = wire860;
              reg891 <= $signed(($unsigned((-$signed(reg843))) ?
                  $unsigned((reg864[(5'h13):(2'h3)] ?
                      ((8'hbf) ~^ reg510) : (reg857 ?
                          reg888 : reg877))) : ({reg889} ?
                      wire435[(3'h4):(3'h4)] : {$unsigned(reg523),
                          reg466,
                          (~&reg842)})));
              reg892 = ($unsigned($signed({(7'h4f), (8'hb4)})) ?
                  {{$signed((!reg449)), (reg504 >= reg524[(1'h0):(1'h0)])},
                      reg491[(5'h17):(4'ha)]} : reg864);
              reg893 = $signed(reg467[(4'h9):(3'h5)]);
              reg894 <= (!(reg878 >> ({$signed(reg856),
                  (reg452 == reg864)} >>> {$signed((8'ha8))})));
            end
          if (reg466[(2'h3):(1'h1)])
            begin
              reg895 <= ({reg845[(4'hc):(3'h7)], reg870} ?
                  $unsigned((($signed(reg463) ^ (~^reg537)) - $signed((reg509 ?
                      wire438 : wire436)))) : $signed((&$signed(reg520))));
            end
          else
            begin
              reg896 = ($signed($signed(($unsigned(reg495) | (8'ha6)))) ?
                  ($unsigned(reg872[(1'h1):(1'h1)]) | ({((8'ha3) ?
                              reg523 : reg885)} ?
                      (&reg533) : ($unsigned(reg889) ?
                          reg895[(4'h9):(3'h7)] : (~|reg443)))) : {reg882,
                      $signed(((~&reg887) || reg883[(4'hd):(4'h8)])),
                      (-((^~reg453) <<< $signed(reg444)))});
              reg897 <= $signed($unsigned(($unsigned({reg530, (8'ha8)}) ?
                  $signed($signed(reg502)) : ($signed(reg464) >> $unsigned((7'h4d))))));
              reg898 <= {(!reg886[(2'h3):(1'h0)])};
              reg899 = $unsigned($unsigned($signed((reg532 ?
                  (reg480 ? reg453 : reg868) : ((8'ha2) ? reg870 : reg898)))));
              reg900 <= ($signed(((|reg536[(5'h17):(3'h6)]) >>> {reg470,
                      (reg466 | (8'hb0)),
                      {reg895, (7'h52), reg530}})) ?
                  ($unsigned(reg467) ?
                      $unsigned($signed($signed(wire436))) : (~|$signed(reg845[(4'hb):(1'h0)]))) : (reg491 ^~ $unsigned(((!reg892) ?
                      {reg503} : $unsigned((8'hb5))))));
              reg901 = $unsigned(($signed($unsigned((reg466 ^ reg511))) && $unsigned(reg894[(3'h7):(2'h3)])));
              reg902 <= (^~(reg854 ? (7'h49) : reg864[(2'h2):(1'h0)]));
            end
          for (forvar903 = (1'h0); (forvar903 < (2'h3)); forvar903 = (forvar903 + (1'h1)))
            begin
              reg904 = (reg842 != (!(&(reg498 + (reg491 ^~ reg864)))));
              reg905 <= ($signed(($unsigned((|(8'hb6))) ?
                      ($signed(reg464) >>> reg444[(1'h1):(1'h1)]) : $signed($signed(reg893)))) ?
                  ($unsigned((reg841 + (reg523 ?
                      wire438 : reg848))) || ($signed((+reg536)) ^~ $unsigned((wire435 ?
                      reg902 : reg517)))) : (8'hb0));
              reg906 = {(~|($unsigned($signed(reg876)) | (forvar903[(3'h4):(1'h0)] ?
                      ((8'hb5) - reg883) : (reg882 ^~ reg901))))};
              reg907 <= reg890[(3'h4):(2'h2)];
              reg908 = (~|reg492);
              reg909 <= $unsigned(reg452);
              reg910 <= {reg444[(2'h2):(1'h0)],
                  (($unsigned($signed((7'h58))) ?
                          reg502 : ($signed((8'h9d)) ?
                              reg906[(3'h5):(3'h4)] : (+(7'h4a)))) ?
                      ($unsigned((reg456 + reg896)) ?
                          ({reg850, wire542, reg487} ?
                              reg482 : {reg896}) : ((~reg444) >> ((7'h48) << reg520))) : (~&({reg479} ?
                          reg864 : {wire439, reg480, reg901}))),
                  reg464[(4'hc):(3'h6)]};
            end
        end
      else
        begin
          reg881 = ((+reg892[(2'h3):(2'h2)]) || $signed(($unsigned(reg890[(3'h4):(3'h4)]) + reg883)));
          reg882 = $unsigned($signed((reg884 ~^ (~^$signed(reg446)))));
        end
      for (forvar911 = (1'h0); (forvar911 < (3'h6)); forvar911 = (forvar911 + (1'h1)))
        begin
          reg912 = {$unsigned((reg517 ?
                  reg876 : ((~reg889) ^~ $unsigned(reg899)))),
              reg877[(5'h17):(1'h0)]};
          if ((!{wire439,
              (((^~reg910) ?
                  {reg521, (7'h56), reg847} : reg892) >= ($signed(reg503) ?
                  (|reg905) : (reg883 >> (8'ha1)))),
              ((~^reg894[(4'hf):(4'hb)]) ?
                  $signed({reg441, reg502}) : ((!reg854) ?
                      ((7'h44) <<< reg476) : (&reg892)))}))
            begin
              reg913 = $signed($signed((($signed(reg489) ^~ reg910) ?
                  $unsigned((reg909 ^~ reg850)) : (reg520[(3'h4):(2'h2)] * reg487))));
              reg914 = reg443;
              reg915 = reg861;
              reg916 <= (~|reg498);
            end
          else
            begin
              reg913 = $signed(reg847[(2'h2):(1'h1)]);
              reg914 = (reg886 ?
                  (~^$signed(reg491[(5'h16):(1'h0)])) : $signed((~^($signed(reg467) ?
                      reg516[(4'h8):(2'h2)] : reg479))));
              reg916 <= ((-reg883) <<< {$unsigned($unsigned({reg442}))});
              reg917 = reg477;
            end
          for (forvar918 = (1'h0); (forvar918 < (3'h6)); forvar918 = (forvar918 + (1'h1)))
            begin
              reg919 <= reg881[(2'h3):(1'h1)];
              reg920 = ((&reg487[(5'h12):(4'ha)]) + (&reg886));
              reg921 = {{($signed(wire437) ? (~^(~|(7'h42))) : (8'hac))}};
              reg922 = (~|($unsigned(reg504) | {(+(reg441 - reg444)),
                  (~^reg882[(2'h3):(1'h1)])}));
              reg923 = $signed(((~((|reg442) ?
                  $signed(reg882) : (reg491 ?
                      (7'h4b) : reg470))) >= $signed($signed((reg896 ?
                  reg867 : reg850)))));
              reg924 = $unsigned((~$signed((^~reg856[(3'h6):(1'h0)]))));
            end
          reg925 = (|$unsigned({((reg897 != reg480) ?
                  (reg876 ? reg923 : reg441) : (reg889 != (8'hb7))),
              (&{reg882, reg890, reg536}),
              ({reg841} ? {reg900, (8'hbf), (8'hb6)} : $signed(reg919))}));
          reg926 <= (^({({reg877,
                  (7'h43),
                  reg876} > (~(7'h4c)))} >> (~&((reg856 - reg453) ?
              $signed(reg847) : (+reg476)))));
          if (($signed((((reg883 >>> (7'h40)) & $unsigned(reg470)) ^~ reg886)) ?
              (-(({reg485} & (~^reg907)) ?
                  $signed(((8'hb3) >= reg925)) : reg537[(1'h0):(1'h0)])) : (&{$signed((reg509 ?
                      reg467 : wire542)),
                  reg892[(4'h9):(2'h3)]})))
            begin
              reg927 = reg491[(5'h15):(4'h9)];
              reg928 = $unsigned($signed((reg881[(1'h0):(1'h0)] & reg464)));
            end
          else
            begin
              reg929 <= reg849;
              reg930 = ((+$signed($signed((reg922 ? reg902 : reg894)))) ?
                  $signed(wire437) : (+reg913));
              reg931 = (reg909[(2'h2):(1'h0)] >> (^(~|$signed($unsigned(reg505)))));
            end
          if ((8'ha1))
            begin
              reg932 <= reg491[(1'h0):(1'h0)];
            end
          else
            begin
              reg933 = (-reg884);
              reg934 = reg453;
              reg935 = reg900[(3'h7):(3'h6)];
              reg936 = (^~(-$unsigned(wire860)));
            end
        end
      for (forvar937 = (1'h0); (forvar937 < (1'h1)); forvar937 = (forvar937 + (1'h1)))
        begin
          reg938 = {forvar937[(1'h0):(1'h0)],
              (~(reg906 <= (^~(-reg470)))),
              (^reg884)};
          reg939 = reg505;
          if ((({$unsigned((!reg841)),
                  ($unsigned(reg913) >>> reg881[(4'hd):(4'hc)]),
                  $unsigned((|reg847))} & (|((reg471 >>> reg864) ?
                  (reg533 ? reg892 : reg938) : wire437))) ?
              {reg461,
                  $signed(forvar903[(3'h5):(3'h5)])} : (((8'ha2) ~^ (~&(^~wire542))) == (reg480[(1'h0):(1'h0)] ?
                  (&$signed(reg896)) : (^~(reg902 ? reg448 : reg932))))))
            begin
              reg940 = ($unsigned(($unsigned($signed(reg929)) >> (reg926 ?
                  (reg938 ?
                      reg916 : reg897) : $signed(reg533)))) & reg901[(2'h2):(1'h0)]);
              reg941 <= reg881;
              reg942 <= reg889[(5'h16):(4'hc)];
              reg943 = (reg485 ?
                  $unsigned(forvar911[(5'h18):(1'h1)]) : (^~(~reg521)));
              reg944 = reg476;
              reg945 <= (8'hab);
              reg946 = $signed((8'hb6));
            end
          else
            begin
              reg941 <= ((^~$unsigned(((reg484 << reg533) << reg489))) ?
                  ($unsigned($signed((8'hb1))) | $signed($unsigned((+reg478)))) : $signed(reg894[(5'h11):(5'h10)]));
              reg943 = reg504[(4'hf):(4'he)];
              reg944 = (reg930 <= $unsigned((($signed(reg902) ?
                  ((8'hac) <= forvar903) : $unsigned(reg914)) <<< reg915[(5'h16):(5'h14)])));
              reg945 <= (reg449 ?
                  $signed((({reg872} ?
                      (reg884 ? wire438 : reg478) : (reg442 ?
                          reg532 : reg931)) == ($unsigned(reg883) ?
                      reg528[(2'h2):(1'h1)] : reg944))) : $signed(({reg870,
                      {reg463, (7'h42)},
                      $signed(reg446)} || (reg514[(1'h0):(1'h0)] ?
                      (reg894 != reg935) : reg877[(4'hb):(2'h2)]))));
              reg946 = reg465;
              reg947 = $unsigned($unsigned($signed($unsigned(((7'h40) >> (8'hb9))))));
            end
          reg948 = {(8'ha6), (&$unsigned($signed($unsigned(reg463))))};
          if (($signed((8'hb5)) * ($unsigned((^~$signed(reg842))) ?
              ((~$unsigned(reg904)) ^~ ((^~reg936) ?
                  $signed(reg466) : $unsigned(reg926))) : (+$unsigned($unsigned((7'h52)))))))
            begin
              reg949 <= $signed((7'h44));
            end
          else
            begin
              reg949 <= $signed({{$unsigned((8'hbd)),
                      $signed(reg924[(2'h3):(1'h1)])}});
              reg950 <= reg938;
              reg951 <= (reg863[(3'h4):(1'h1)] == (~^$signed($signed((reg925 ?
                  (8'hb4) : reg934)))));
            end
          if (wire437)
            begin
              reg952 = $unsigned($unsigned(reg928));
            end
          else
            begin
              reg952 = ((({$signed(reg927), (reg951 ? reg441 : (8'ha3))} ?
                      reg520[(2'h2):(1'h1)] : $signed(((8'h9c) >>> reg936))) ?
                  (~|reg917[(4'hf):(2'h2)]) : $signed((~^forvar903[(1'h1):(1'h0)]))) <= {$signed($signed({reg484,
                      (8'hbf)})),
                  ($unsigned((&reg883)) ?
                      $unsigned((&reg947)) : (|reg931[(1'h1):(1'h1)])),
                  wire542});
              reg953 = (reg507 ? reg456[(4'hb):(3'h4)] : reg882[(1'h1):(1'h1)]);
              reg954 = reg477;
            end
        end
      for (forvar955 = (1'h0); (forvar955 < (3'h6)); forvar955 = (forvar955 + (1'h1)))
        begin
          if ($signed((wire838[(5'h13):(2'h3)] ~^ $signed(reg885))))
            begin
              reg956 <= reg894[(5'h1e):(5'h19)];
              reg957 <= ($signed(($unsigned($unsigned((7'h49))) | (reg896 + $unsigned(reg456)))) ?
                  reg848 : reg482);
            end
          else
            begin
              reg958 = $unsigned($unsigned(reg882));
              reg959 = (reg930 << (^~(^(|$signed(reg882)))));
            end
          if (reg507[(2'h3):(1'h0)])
            begin
              reg960 <= ({reg463[(5'h1a):(5'h19)],
                      $unsigned($signed(reg532)),
                      $signed(({wire437} << reg505))} ?
                  reg959[(4'hc):(4'h9)] : $signed($unsigned(reg941)));
              reg961 = ($signed((-({reg901, reg478, reg951} >= reg861))) ?
                  reg441 : (reg476[(3'h4):(3'h4)] ^~ reg887));
              reg962 = reg881;
            end
          else
            begin
              reg960 <= $unsigned({(reg864[(4'hc):(4'ha)] >> ((reg962 <= reg866) ?
                      reg895 : $signed(reg948))),
                  ({(8'hab)} <= ($unsigned(reg467) ?
                      (reg919 ? reg514 : reg864) : reg456[(4'h8):(1'h0)]))});
              reg963 <= (8'h9c);
              reg964 = reg489;
            end
          reg965 = reg523;
          reg966 = (~|$unsigned(reg866[(1'h1):(1'h0)]));
        end
      reg967 = reg840;
    end
  always
    @(posedge clk) begin
      reg968 <= ($unsigned((&(^reg524[(3'h6):(1'h0)]))) ?
          $unsigned((((reg536 && reg464) >>> reg482) >> wire439)) : reg950);
      reg969 = {(reg465 <= reg902[(4'h8):(4'h8)]), reg888[(4'h8):(4'h8)]};
    end
  always
    @(posedge clk) begin
      if ((~$unsigned((8'h9f))))
        begin
          reg970 <= (|$signed((reg951 ?
              $signed(reg867) : $signed((reg876 ~^ reg473)))));
          if (({(((reg461 ? (8'hbe) : (7'h43)) ?
                  reg487[(4'hc):(4'h8)] : (reg504 | wire436)) << reg968[(2'h3):(2'h2)]),
              $signed(reg461),
              (~&reg509[(4'h9):(3'h5)])} ~^ {reg841[(4'hc):(4'h9)],
              reg514[(1'h1):(1'h0)],
              ((|$unsigned(reg452)) >> ($unsigned(reg505) > $unsigned(reg456)))}))
            begin
              reg971 <= (~^wire838);
              reg972 = reg950;
              reg973 = (-$signed($unsigned((!(reg867 ? reg480 : reg884)))));
              reg974 = reg864;
              reg975 = $signed(reg452[(4'h8):(3'h7)]);
              reg976 <= ($signed($unsigned({(-reg888),
                      (reg867 ? reg975 : reg950),
                      (^wire437)})) ?
                  (~&$unsigned(((wire838 >>> (7'h53)) < $unsigned(reg524)))) : (^~(($unsigned(reg945) * (+reg446)) + reg489)));
              reg977 <= reg895;
            end
          else
            begin
              reg971 <= reg523;
              reg976 <= (reg895 >> (~&reg476[(2'h3):(2'h2)]));
              reg977 <= (-((reg949[(3'h6):(1'h1)] && ((7'h54) ?
                      ((8'haa) || (8'hb9)) : (reg461 ? reg963 : reg521))) ?
                  $unsigned((reg452[(3'h6):(3'h4)] <= $signed((8'ha1)))) : reg866[(1'h0):(1'h0)]));
              reg978 <= reg977;
              reg979 = reg536;
            end
          reg980 <= $unsigned((~^(|(reg532 - (reg877 << reg885)))));
          reg981 = reg897[(5'h10):(4'hf)];
          reg982 = reg541[(2'h3):(2'h2)];
          for (forvar983 = (1'h0); (forvar983 < (3'h4)); forvar983 = (forvar983 + (1'h1)))
            begin
              reg984 = (~&(~&((reg876 ?
                  ((8'hbb) ?
                      (8'hb3) : reg963) : {reg511}) <<< ((~reg448) ^ (reg476 <<< reg464)))));
              reg985 <= reg520[(5'h14):(4'he)];
              reg986 = reg446;
              reg987 = {$unsigned(reg464)};
              reg988 <= {reg528[(1'h0):(1'h0)]};
              reg989 <= (({reg905,
                      ($unsigned(reg511) ? $signed(wire438) : $signed(reg443)),
                      reg466[(3'h4):(1'h1)]} ?
                  $unsigned({(reg471 ?
                          reg480 : reg533)}) : (reg477 <<< reg974[(1'h1):(1'h1)])) >= reg883);
              reg990 <= $unsigned((reg856[(4'hd):(3'h7)] < reg986[(5'h10):(3'h4)]));
            end
        end
      else
        begin
          reg970 <= reg872;
        end
      if ($unsigned(reg849))
        begin
          if (reg861)
            begin
              reg991 = ((reg528[(3'h5):(3'h5)] ?
                      reg471[(2'h3):(1'h0)] : $unsigned(reg972[(5'h11):(4'h9)])) ?
                  {({reg988[(1'h1):(1'h1)], $unsigned(reg910), (^~reg471)} ?
                          (wire435 - {reg537, reg469, (8'hb9)}) : (~((7'h49) ?
                              reg536 : reg479)))} : (8'haa));
              reg992 = (reg476 <<< reg979[(3'h7):(3'h4)]);
              reg993 <= (reg987[(3'h7):(1'h0)] ?
                  $signed($unsigned((reg504[(5'h10):(4'h9)] ?
                      (&reg919) : $unsigned(reg990)))) : (|$signed(reg980[(2'h2):(2'h2)])));
              reg994 = reg876[(3'h6):(2'h3)];
            end
          else
            begin
              reg993 <= (^~forvar983[(2'h2):(1'h1)]);
              reg995 <= $unsigned((~{((reg932 ? reg477 : reg524) ?
                      reg900[(3'h4):(3'h4)] : (!reg847)),
                  reg510,
                  reg885[(4'hc):(3'h7)]}));
              reg996 <= $unsigned($signed($unsigned(((&reg929) ?
                  $signed(reg970) : (+forvar983)))));
            end
        end
      else
        begin
          reg993 <= ((^~reg971) ^~ (~(reg457 ^ reg979)));
          reg995 <= $signed(((^~$signed((reg516 && reg482))) ^~ (reg456 ?
              reg989[(5'h16):(4'he)] : reg521[(4'ha):(4'h8)])));
          for (forvar996 = (1'h0); (forvar996 < (1'h1)); forvar996 = (forvar996 + (1'h1)))
            begin
              reg997 <= (reg885 ?
                  $unsigned($unsigned($unsigned($signed(reg505)))) : $signed($signed((reg891[(3'h6):(2'h2)] > $unsigned(reg517)))));
              reg998 <= (&(reg847 <<< $unsigned($signed((wire439 ?
                  reg978 : reg850)))));
              reg999 <= $signed($signed((~|$signed(reg891))));
              reg1000 = (($signed(((reg465 <<< reg471) ~^ reg949)) ^ ($unsigned(reg868[(3'h7):(3'h7)]) ?
                      reg977 : (reg516[(5'h13):(4'hd)] <<< reg528[(1'h0):(1'h0)]))) ?
                  ((reg979 * (7'h54)) >> ((^$unsigned(reg990)) ?
                      reg849[(1'h1):(1'h1)] : $signed((reg888 ^ reg504)))) : $signed(reg850));
            end
          for (forvar1001 = (1'h0); (forvar1001 < (2'h3)); forvar1001 = (forvar1001 + (1'h1)))
            begin
              reg1002 = (~^reg510);
              reg1003 = $unsigned($unsigned(({(reg504 ^ reg484),
                      (reg872 | forvar996)} ?
                  reg509[(3'h5):(3'h5)] : ($signed(reg932) ?
                      (wire437 ? (7'h56) : (8'hb6)) : (reg963 ?
                          reg894 : reg854)))));
              reg1004 <= (reg889[(3'h6):(1'h1)] || reg894);
              reg1005 = $unsigned($signed($signed({reg968[(4'hc):(2'h2)],
                  (wire439 ? reg479 : forvar996)})));
              reg1006 = (reg465[(3'h5):(2'h2)] ?
                  {$unsigned(($unsigned(reg971) ?
                          (reg467 ?
                              reg471 : reg847) : reg484[(3'h6):(1'h1)]))} : (wire437 ?
                      (reg878 ?
                          ((^reg973) - $unsigned((7'h54))) : (8'ha2)) : wire438));
            end
        end
      reg1007 = reg956;
      reg1008 = reg950[(5'h10):(4'hd)];
    end
  always
    @(posedge clk) begin
      reg1009 = ($unsigned($signed((8'h9d))) ? (^reg884) : reg469);
      if (reg441)
        begin
          reg1010 = $unsigned(($unsigned(((~^reg509) <= reg907[(1'h1):(1'h0)])) <<< $signed(reg856)));
          for (forvar1011 = (1'h0); (forvar1011 < (1'h1)); forvar1011 = (forvar1011 + (1'h1)))
            begin
              reg1012 = (-({reg456[(5'h13):(4'h8)]} - (~&{(+reg870)})));
              reg1013 = (7'h4e);
              reg1014 = reg466;
              reg1015 = ($unsigned((($unsigned((8'hbf)) ?
                          (~&reg505) : {wire438}) ?
                      (~^$unsigned(reg861)) : $unsigned((reg1012 | reg960)))) ?
                  {$signed((+(reg872 ? reg533 : (8'ha6))))} : {$signed(reg941),
                      $signed($signed($unsigned(reg861)))});
              reg1016 <= $unsigned(wire860[(5'h1f):(3'h4)]);
              reg1017 <= ($signed(reg848) ?
                  reg905 : (~^(reg894 >> (reg876 ?
                      wire542[(2'h3):(1'h0)] : (reg446 == reg498)))));
            end
          for (forvar1018 = (1'h0); (forvar1018 < (2'h2)); forvar1018 = (forvar1018 + (1'h1)))
            begin
              reg1019 = $signed((reg877 ?
                  {$unsigned((&wire435)),
                      $unsigned({reg976}),
                      reg541[(3'h5):(1'h1)]} : {($signed(reg988) ?
                          {reg491, reg523} : $signed(reg1017))}));
              reg1020 <= (^reg884);
              reg1021 <= {(~&$unsigned($signed($signed(wire860))))};
              reg1022 <= {$signed(reg1021[(5'h13):(4'hb)])};
              reg1023 = (&(($signed((reg848 ? (8'ha9) : reg963)) ?
                      ((reg467 ? (7'h4a) : reg520) ?
                          reg898[(1'h0):(1'h0)] : $unsigned(reg910)) : (reg840 ?
                          $signed(reg443) : (!reg988))) ?
                  $signed((reg1021[(2'h3):(1'h0)] ?
                      (~reg848) : $signed(reg463))) : $signed((reg480 ?
                      {reg895} : (8'hbf)))));
            end
          if ((!wire437[(3'h4):(3'h4)]))
            begin
              reg1024 = ((reg487 << ($signed($unsigned(reg868)) ?
                  reg996[(4'ha):(2'h2)] : reg530[(4'hb):(4'ha)])) - ((~^$signed(reg990)) ?
                  reg951 : (-(reg997 ? $unsigned(reg1017) : reg1012))));
              reg1025 = $unsigned($unsigned($unsigned(((^reg854) ?
                  $signed(reg998) : (reg537 ? reg467 : reg524)))));
              reg1026 = $signed((~&reg479[(2'h3):(1'h1)]));
            end
          else
            begin
              reg1027 <= reg902;
              reg1028 = (7'h58);
              reg1029 = $unsigned($signed(reg480));
              reg1030 <= ((((|(~&reg470)) | (~(|reg514))) ?
                  reg1004 : reg502[(3'h4):(3'h4)]) & ((-(7'h40)) << (reg850 ?
                  $unsigned(reg1029) : ($unsigned(reg1021) - $signed(reg1024)))));
              reg1031 <= ($signed((&reg466[(1'h0):(1'h0)])) ?
                  $unsigned(reg1012[(4'ha):(1'h1)]) : (~($signed(((7'h4f) << reg529)) ?
                      (reg504[(5'h11):(5'h10)] ?
                          $signed(reg856) : reg866[(1'h0):(1'h0)]) : $signed(reg498))));
              reg1032 = (|reg861[(4'he):(2'h2)]);
              reg1033 <= reg902;
            end
          reg1034 = (reg877 ? reg457 : $unsigned(reg446));
          for (forvar1035 = (1'h0); (forvar1035 < (3'h4)); forvar1035 = (forvar1035 + (1'h1)))
            begin
              reg1036 <= (^~(8'hb7));
              reg1037 <= ($unsigned(($unsigned(reg840) == $signed(reg872[(3'h7):(1'h0)]))) ?
                  {{((reg530 ^ reg883) && (reg878 ?
                              reg480 : reg463))}} : (~|($unsigned((reg866 ?
                      (7'h43) : reg842)) || $signed((8'hb8)))));
            end
        end
      else
        begin
          for (forvar1010 = (1'h0); (forvar1010 < (2'h2)); forvar1010 = (forvar1010 + (1'h1)))
            begin
              reg1011 <= (reg849 | $signed(($signed({reg476,
                  reg495,
                  reg467}) != ((reg850 * forvar1011) ? {reg1034} : reg905))));
            end
          reg1016 <= (8'hb9);
        end
      reg1038 = {reg956[(1'h1):(1'h1)],
          ($unsigned(reg466[(2'h2):(1'h1)]) ?
              $signed((reg465 ?
                  (reg897 ?
                      (7'h4a) : reg988) : (|reg857))) : $signed((reg484 * reg854)))};
      if ((((reg910[(1'h1):(1'h1)] ?
              ({reg1024, reg963, (7'h56)} > (reg870 ?
                  forvar1018 : reg945)) : ((^reg1029) << reg1031)) >>> (8'hb9)) ?
          (~($signed($signed(reg847)) == $unsigned((reg495 ?
              reg1021 : reg845)))) : $signed($signed(reg461[(4'he):(4'ha)]))))
        begin
          reg1039 = {((+reg471[(3'h5):(3'h4)]) ?
                  reg932 : $unsigned($signed(reg444[(2'h2):(2'h2)]))),
              ((~((|reg872) ? $signed(reg877) : ((8'ha4) ~^ reg505))) ?
                  (reg1021 && reg951[(2'h2):(1'h1)]) : $signed(((~^reg878) ?
                      $unsigned((8'ha6)) : reg1015)))};
          reg1040 <= {reg520[(4'hb):(2'h2)]};
          reg1041 <= ({((~|$signed(reg995)) * reg849[(2'h2):(1'h1)]),
              (~^reg877[(2'h2):(1'h1)]),
              $signed((reg1037[(4'hc):(2'h2)] + reg877))} || $signed($unsigned(($signed(reg847) * $unsigned(reg510)))));
          if ($signed(((reg442 >= {$unsigned(reg530)}) <= $signed(($unsigned(reg1014) ?
              $unsigned(wire439) : $unsigned(forvar1035))))))
            begin
              reg1042 = $signed($signed(reg968));
            end
          else
            begin
              reg1042 = (^($signed((|(reg492 ?
                  wire436 : (8'hbd)))) ^~ {($signed(reg884) ?
                      {reg988, reg498} : (wire438 ? reg895 : forvar1035)),
                  reg840,
                  ({reg463, reg466, wire436} | (reg863 << reg1022))}));
            end
        end
      else
        begin
          for (forvar1039 = (1'h0); (forvar1039 < (1'h0)); forvar1039 = (forvar1039 + (1'h1)))
            begin
              reg1040 <= $signed($unsigned((+$signed($signed(reg1021)))));
              reg1042 = reg997[(4'hf):(2'h3)];
              reg1043 = {$unsigned({wire838[(4'ha):(4'h8)], (8'hb0), reg960}),
                  (|$signed({$signed((7'h56)),
                      reg970[(4'h8):(2'h2)],
                      $unsigned(forvar1010)})),
                  (&((reg1004[(2'h3):(1'h1)] ?
                      reg995[(5'h12):(4'hb)] : (~^reg446)) & reg457))};
              reg1044 = {$signed((reg523[(4'hf):(4'h9)] ?
                      $signed(reg999) : (^(reg942 ? reg502 : reg1014))))};
              reg1045 = $unsigned(reg468);
              reg1046 <= $signed($signed((|reg1014)));
            end
          if ((+$unsigned(reg863[(4'hc):(3'h4)])))
            begin
              reg1047 <= $signed(reg847);
              reg1048 = (^~reg476);
            end
          else
            begin
              reg1047 <= reg995[(3'h5):(3'h5)];
            end
          if (reg465[(4'h8):(2'h2)])
            begin
              reg1049 <= {{((reg916[(4'h8):(1'h0)] ^~ (+(7'h47))) ?
                          {$unsigned(reg980), $unsigned(reg857)} : (8'hb8)),
                      $unsigned(reg1010)},
                  ({(((8'ha1) >= wire838) > $unsigned(reg452)),
                      (^~reg503),
                      $signed((8'hbd))} != $signed(reg495)),
                  {reg471, (~reg532), $unsigned($unsigned(reg900))}};
              reg1050 = ($unsigned((~((^reg1033) == reg950))) ?
                  $signed($signed(reg511[(3'h5):(2'h2)])) : {{(((8'hb8) ?
                              (8'hbf) : reg491) || $unsigned(reg902)),
                          reg849[(2'h2):(1'h1)]},
                      ({(~|reg485), (reg985 <= reg446)} ?
                          ({(7'h58),
                              reg492} + $unsigned(reg505)) : $unsigned(reg883))});
              reg1051 <= {((8'ha3) >= ((|$signed(reg929)) <= $signed(reg889))),
                  $unsigned((8'ha1)),
                  ($unsigned(reg1041) >>> (~^((reg843 >>> forvar1039) ?
                      (reg471 ? reg1034 : reg885) : {reg1039,
                          reg1044,
                          reg998})))};
              reg1052 = (&$signed((reg842 ^~ $unsigned({reg988}))));
              reg1053 = ((^~(((reg1051 >= reg883) ?
                      reg495[(3'h4):(2'h3)] : (reg1052 ? reg530 : (7'h57))) ?
                  (wire437 ?
                      (reg524 ?
                          reg1010 : reg970) : (~|(8'hab))) : ($unsigned(forvar1010) ~^ (reg988 ?
                      reg469 : reg471)))) ^ (reg998 ?
                  (+$unsigned({reg536})) : (reg1017[(3'h4):(1'h0)] ?
                      reg529[(1'h1):(1'h1)] : reg1033)));
              reg1054 = reg887;
              reg1055 <= ((reg1022 >>> reg492) + reg482);
            end
          else
            begin
              reg1050 = {(|reg457[(4'hd):(4'ha)])};
              reg1051 <= $signed(($signed({(reg857 == reg1012)}) ?
                  (~$unsigned((reg929 && (8'hb6)))) : {($unsigned((8'hb6)) == reg998)}));
              reg1052 = (~&reg1012[(3'h6):(1'h1)]);
              reg1055 <= (+$signed((|(reg478 ^ $unsigned(reg897)))));
              reg1056 = reg495[(3'h5):(1'h1)];
              reg1057 = (8'hbb);
            end
          reg1058 <= reg997[(3'h4):(1'h1)];
        end
    end
  assign wire1059 = (8'hb1);
  module1060 #() modinst1245 (.y(wire1244), .clk(clk), .wire1066(reg902), .wire1061(reg867), .wire1065(reg457), .wire1064(reg857), .wire1062(reg521), .wire1063(reg888));
  assign wire1246 = (($unsigned((reg932 ?
                            $unsigned(wire542) : (reg1047 ?
                                reg1051 : reg509))) ?
                        $unsigned(wire439[(1'h0):(1'h0)]) : (8'hb6)) >>> ((((reg950 << (7'h42)) > (reg1004 ?
                            reg885 : wire838)) <<< reg847) ?
                        ($unsigned({reg842}) >>> $unsigned(reg1058[(1'h1):(1'h1)])) : $unsigned(reg898)));
  assign wire1247 = reg941;
  always
    @(posedge clk) begin
      reg1248 = reg443[(5'h10):(2'h3)];
      for (forvar1249 = (1'h0); (forvar1249 < (1'h1)); forvar1249 = (forvar1249 + (1'h1)))
        begin
          for (forvar1250 = (1'h0); (forvar1250 < (2'h3)); forvar1250 = (forvar1250 + (1'h1)))
            begin
              reg1251 <= $unsigned(($signed(wire542) ^ ({$unsigned(reg978)} - $unsigned(reg1040))));
              reg1252 <= ((+$unsigned({(7'h4a)})) && $signed($unsigned(((reg517 ?
                  reg1031 : (7'h54)) >> reg1011))));
              reg1253 = reg541[(2'h2):(1'h1)];
              reg1254 <= reg985[(2'h2):(1'h0)];
              reg1255 <= $unsigned((((~^(reg963 <= wire1244)) ~^ $signed(wire1246[(1'h0):(1'h0)])) > {$signed($unsigned((8'hbc))),
                  reg841,
                  ($signed(reg995) >= reg1033)}));
              reg1256 = wire838;
            end
          reg1257 <= $signed(reg988[(3'h5):(3'h5)]);
          reg1258 <= ((^~(+$signed(reg517))) ?
              $unsigned({wire1247[(3'h4):(2'h2)],
                  (~$unsigned(reg957)),
                  (reg511 >> (!(7'h4a)))}) : reg849);
          if ((reg1037 ?
              ($signed({reg990[(2'h2):(1'h0)]}) ?
                  $signed((~&reg504[(4'hf):(3'h7)])) : reg502[(4'h9):(2'h3)]) : reg878[(4'h8):(2'h3)]))
            begin
              reg1259 = reg529[(3'h4):(2'h2)];
              reg1260 <= (-(7'h45));
            end
          else
            begin
              reg1260 <= $unsigned((^~(8'hb9)));
              reg1261 = reg887[(5'h11):(4'h9)];
              reg1262 <= (reg1022[(5'h10):(4'h8)] ~^ ($signed($unsigned(wire437)) ?
                  {$unsigned($unsigned((7'h54)))} : $unsigned($signed(reg457))));
              reg1263 = $signed($signed({(reg1046 ? forvar1249 : (+reg996))}));
              reg1264 <= (^~((~$signed($signed(reg482))) || reg495));
            end
          reg1265 = reg480[(2'h2):(1'h0)];
          reg1266 = reg960[(1'h0):(1'h0)];
        end
      for (forvar1267 = (1'h0); (forvar1267 < (3'h4)); forvar1267 = (forvar1267 + (1'h1)))
        begin
          reg1268 = {$unsigned(reg1030[(3'h5):(2'h3)]),
              (^~reg877),
              reg963[(3'h5):(1'h1)]};
          for (forvar1269 = (1'h0); (forvar1269 < (3'h4)); forvar1269 = (forvar1269 + (1'h1)))
            begin
              reg1270 = (reg532 >= $signed(reg507[(4'h9):(3'h7)]));
              reg1271 <= ($unsigned(reg980[(4'hb):(1'h1)]) >> $unsigned((+$signed($signed(reg514)))));
              reg1272 <= reg894[(5'h17):(1'h0)];
            end
          reg1273 = reg997;
          reg1274 <= (~|(({(reg482 ? wire1059 : reg1251), (~|(7'h46))} ?
              (reg467[(4'h9):(2'h2)] ?
                  reg848 : reg900) : (+(reg487 > reg949))) >> reg530));
        end
      for (forvar1275 = (1'h0); (forvar1275 < (3'h5)); forvar1275 = (forvar1275 + (1'h1)))
        begin
          if ((reg521 < (((~&(&reg1259)) && $unsigned($signed(reg909))) ?
              reg1022[(1'h1):(1'h0)] : $unsigned(reg1262[(4'h9):(3'h6)]))))
            begin
              reg1276 <= $signed(reg478);
              reg1277 <= reg1058;
              reg1278 <= $unsigned({reg1271,
                  (!((8'hb3) >= $signed(reg999))),
                  $unsigned(((reg1248 ? reg1266 : reg1037) ?
                      $signed(reg857) : (reg1254 ? reg1264 : (8'h9e))))});
              reg1279 <= ($signed(reg1027) < ((wire437 & reg480) ?
                  (reg1040[(1'h0):(1'h0)] > {reg521,
                      (forvar1269 ^~ reg1253),
                      (reg529 && (7'h54))}) : $signed(((reg883 ?
                      reg509 : reg465) == (reg885 == reg949)))));
              reg1280 = ($unsigned($unsigned({{reg1274}})) ?
                  (reg1258 | $unsigned({(reg971 ?
                          reg520 : reg485)})) : (~&(&(~|{(7'h42),
                      reg864,
                      reg867}))));
              reg1281 = $signed(reg872[(3'h5):(2'h3)]);
              reg1282 = ($unsigned((forvar1267 && (^(reg1276 <<< reg1055)))) ?
                  {(~|reg850),
                      reg1261,
                      $unsigned($signed((reg971 < reg1271)))} : (reg1262 ?
                      {(|{reg1011, reg910, reg907}),
                          reg537,
                          ((reg482 ^ reg516) ?
                              {reg1252} : reg945)} : ((|$unsigned(reg465)) ?
                          (~reg993) : (~reg1253))));
            end
          else
            begin
              reg1276 <= (({reg877,
                  $unsigned({reg530}),
                  (~&$signed(reg1273))} == (&reg926)) ^ (~&reg876[(4'he):(4'ha)]));
              reg1280 = ($unsigned(wire1246) && (!reg473[(1'h0):(1'h0)]));
              reg1281 = reg470[(1'h0):(1'h0)];
              reg1282 = reg485;
              reg1283 <= ($unsigned(reg845[(4'hc):(4'hc)]) ? (7'h4c) : reg1281);
              reg1284 = (+reg867);
            end
          reg1285 <= $signed((7'h51));
          reg1286 = (&$unsigned({reg509[(4'h9):(2'h2)],
              $unsigned(((8'h9d) ? reg978 : reg1051)),
              {reg537[(2'h2):(2'h2)]}}));
          for (forvar1287 = (1'h0); (forvar1287 < (2'h2)); forvar1287 = (forvar1287 + (1'h1)))
            begin
              reg1288 = ((7'h54) ~^ ((8'ha9) ?
                  $signed(reg905) : (((reg970 > reg856) ?
                          $unsigned(reg464) : {reg971}) ?
                      $signed(((7'h4d) | reg900)) : (^reg840[(3'h7):(3'h4)]))));
              reg1289 = {{(reg919[(4'hd):(4'ha)] * $signed({reg476, reg471}))}};
              reg1290 <= $signed(($unsigned((reg464 <= reg849[(3'h4):(2'h3)])) << reg1049));
              reg1291 = ((((!reg985[(1'h0):(1'h0)]) > reg1274[(1'h1):(1'h0)]) ?
                  (7'h40) : $signed(reg884)) >>> (&{$signed(reg977)}));
              reg1292 <= {reg1046[(2'h2):(1'h1)],
                  (forvar1269 ?
                      $signed(reg999[(4'hd):(3'h6)]) : reg956[(2'h2):(1'h0)]),
                  (~&reg1254[(1'h1):(1'h1)])};
              reg1293 = {$unsigned(reg453),
                  (^~reg857[(5'h11):(1'h1)]),
                  reg1282};
            end
          if (reg883[(1'h1):(1'h0)])
            begin
              reg1294 <= reg1266[(2'h3):(2'h3)];
              reg1295 <= (reg1253[(4'he):(2'h3)] <<< $signed((7'h4b)));
            end
          else
            begin
              reg1294 <= $signed((|(8'hb5)));
              reg1296 = wire435;
            end
          if (($unsigned($signed($unsigned($signed(reg1252)))) ?
              (($signed(forvar1275[(2'h2):(1'h1)]) <<< (~&(reg1040 ?
                  (7'h43) : reg1017))) || reg895[(3'h7):(3'h6)]) : $unsigned(reg1268)))
            begin
              reg1297 = $signed(((-($signed(reg1283) ~^ ((8'ha0) ?
                  reg1285 : reg1257))) ^~ (&reg842[(2'h2):(1'h0)])));
              reg1298 = $signed(reg464[(5'h16):(5'h14)]);
              reg1299 <= reg877;
              reg1300 = reg489;
              reg1301 <= reg1263[(4'hc):(1'h0)];
              reg1302 <= (wire435 ?
                  reg1037 : (reg866[(3'h6):(1'h1)] ?
                      {reg489} : reg1262[(1'h0):(1'h0)]));
            end
          else
            begin
              reg1297 = reg448[(3'h5):(1'h0)];
              reg1298 = reg884;
              reg1300 = $signed($signed(reg977));
              reg1303 = $unsigned((8'hba));
            end
        end
      reg1304 = wire1244;
      for (forvar1305 = (1'h0); (forvar1305 < (3'h4)); forvar1305 = (forvar1305 + (1'h1)))
        begin
          reg1306 <= (~|$unsigned($unsigned(((reg452 ?
              reg1031 : reg950) & reg945[(4'he):(2'h3)]))));
          reg1307 <= {(reg872[(4'hf):(4'h8)] + (reg883 ?
                  ((~|wire435) >>> $unsigned(wire860)) : reg856[(5'h10):(3'h6)])),
              $unsigned($unsigned(((reg1301 >= reg905) == reg996)))};
          reg1308 <= $signed((($unsigned($unsigned(reg950)) ?
              (reg950 ^ {reg854,
                  reg847,
                  reg517}) : (~$signed(reg968))) >>> {$unsigned($signed(reg457))}));
          if (reg537)
            begin
              reg1309 = ((reg1017[(4'ha):(3'h7)] ?
                  reg900[(3'h6):(2'h2)] : ((~^(7'h4d)) + reg900)) || ((!reg504[(4'hf):(3'h4)]) & reg970[(1'h0):(1'h0)]));
              reg1310 <= $unsigned(reg1031);
            end
          else
            begin
              reg1309 = (reg1254[(3'h5):(3'h4)] ?
                  {((~&reg1284[(4'h8):(2'h2)]) ?
                          $unsigned(((8'ha3) | reg1049)) : reg1307[(5'h11):(2'h2)]),
                      {((-reg989) ?
                              (reg467 ? reg1268 : reg898) : {reg469,
                                  reg1031})}} : reg976[(5'h17):(5'h15)]);
            end
        end
      for (forvar1311 = (1'h0); (forvar1311 < (3'h4)); forvar1311 = (forvar1311 + (1'h1)))
        begin
          if ((reg523[(4'he):(4'h9)] * reg1282[(4'h9):(2'h2)]))
            begin
              reg1312 <= reg1271[(1'h0):(1'h0)];
              reg1313 <= ((($unsigned(reg1301[(4'h8):(1'h1)]) << reg891[(3'h5):(2'h3)]) ?
                  $signed(reg441[(4'hf):(3'h7)]) : ({$unsigned(reg1263),
                      $unsigned(reg533)} <= (&(reg1296 ?
                      (8'hae) : reg950)))) != (|reg861));
              reg1314 = reg465;
              reg1315 = reg985;
              reg1316 = reg1058;
              reg1317 <= reg1296[(3'h4):(2'h2)];
              reg1318 = ((reg1284 ^~ (&reg900)) & ($signed((reg478[(4'hb):(3'h6)] <<< $unsigned(reg1016))) && $unsigned((|{wire860,
                  (8'ha8)}))));
            end
          else
            begin
              reg1312 <= (-{$unsigned(forvar1287),
                  (^~$unsigned(reg471[(2'h3):(1'h1)]))});
              reg1313 <= (reg1317 ?
                  {reg848[(1'h0):(1'h0)],
                      $signed(reg521),
                      $unsigned({{reg509, reg541},
                          ((7'h4b) ?
                              reg997 : (8'ha1))})} : $signed(reg442[(5'h1a):(4'hf)]));
            end
          reg1319 <= reg467[(1'h0):(1'h0)];
          reg1320 <= $signed($unsigned(((8'hab) ^ reg446)));
          for (forvar1321 = (1'h0); (forvar1321 < (1'h1)); forvar1321 = (forvar1321 + (1'h1)))
            begin
              reg1322 <= (reg1021[(5'h18):(5'h14)] ?
                  $unsigned((|(!wire437[(5'h11):(4'hc)]))) : {($signed($signed((7'h54))) <<< (|reg894)),
                      $signed(($signed(reg1268) >> (|reg469))),
                      {{$unsigned(wire436), wire435, reg541}, reg1255}});
              reg1323 <= ((^$signed((reg1258 & (reg473 ? reg1027 : reg867)))) ?
                  (($unsigned(reg1292[(2'h3):(2'h2)]) ?
                      $unsigned(reg1021[(5'h10):(5'h10)]) : reg883) < (~reg878[(1'h1):(1'h0)])) : {$signed((reg885[(1'h1):(1'h0)] ?
                          $unsigned(reg444) : reg492[(3'h4):(1'h1)]))});
              reg1324 = $signed((!$unsigned($signed((~reg449)))));
            end
          reg1325 = $unsigned((((reg895 ~^ reg1314[(5'h15):(1'h1)]) - reg1259) ?
              $signed($unsigned((^~reg850))) : $unsigned((((8'had) ?
                  reg504 : reg1292) ~^ reg910[(1'h1):(1'h0)]))));
        end
    end
  always
    @(posedge clk) begin
      reg1326 = {reg905[(2'h3):(2'h3)]};
      reg1327 <= $signed({reg478, $unsigned($signed(reg883[(4'hd):(3'h7)]))});
      if ((reg848[(1'h1):(1'h1)] >>> $signed(reg529[(3'h6):(3'h4)])))
        begin
          reg1328 = reg457;
        end
      else
        begin
          for (forvar1328 = (1'h0); (forvar1328 < (2'h2)); forvar1328 = (forvar1328 + (1'h1)))
            begin
              reg1329 = ((~&(wire435[(1'h1):(1'h1)] & (!$signed(reg1290)))) <= ((reg843[(5'h18):(3'h4)] ?
                  ($signed(reg510) ? $signed(reg541) : reg1041) : (^~(reg1260 ?
                      reg503 : reg484))) ^ {$unsigned(reg850)}));
              reg1330 <= reg1279;
              reg1331 <= (reg1302[(4'h9):(4'h8)] ?
                  $unsigned((7'h40)) : (~(^~(&reg910))));
              reg1332 = $signed((reg980[(4'he):(3'h4)] ?
                  $unsigned($unsigned(((8'haf) ?
                      reg467 : reg889))) : $unsigned((^{(8'haa), reg870}))));
              reg1333 = {reg999[(4'hc):(4'ha)],
                  $signed(($unsigned(reg1046[(4'hf):(4'hd)]) ?
                      reg449[(2'h2):(1'h1)] : reg999[(2'h3):(2'h3)]))};
              reg1334 <= ((8'had) ?
                  (reg456 * ($unsigned((&reg452)) ?
                      (!$unsigned(reg537)) : (reg491[(1'h0):(1'h0)] ?
                          (reg487 ?
                              wire838 : (7'h4c)) : $signed(reg449)))) : $unsigned((+($signed(reg919) ?
                      (!(8'hb7)) : (reg461 == reg996)))));
              reg1335 <= ((reg850[(3'h4):(3'h4)] & (reg476 | (^reg1033[(4'h8):(3'h7)]))) ?
                  reg907[(1'h1):(1'h1)] : reg441);
            end
          for (forvar1336 = (1'h0); (forvar1336 < (1'h1)); forvar1336 = (forvar1336 + (1'h1)))
            begin
              reg1337 <= $signed(reg861);
              reg1338 = wire437[(4'h9):(3'h6)];
              reg1339 <= $signed(((reg1332[(4'h8):(3'h6)] <<< (~|(reg469 != reg1022))) ?
                  $signed((|reg1016[(2'h2):(1'h1)])) : {reg449[(1'h1):(1'h1)],
                      (7'h56)}));
              reg1340 = $unsigned($unsigned($signed($unsigned($unsigned(reg510)))));
            end
          reg1341 <= $unsigned({(($signed(reg495) ~^ $signed(reg897)) >= (|reg976[(4'h9):(2'h2)]))});
          reg1342 = ($unsigned((7'h44)) ^ (reg528[(1'h0):(1'h0)] >> reg945[(4'h9):(1'h0)]));
          for (forvar1343 = (1'h0); (forvar1343 < (2'h2)); forvar1343 = (forvar1343 + (1'h1)))
            begin
              reg1344 <= {((!reg1027[(1'h1):(1'h1)]) ?
                      (reg1258[(5'h13):(3'h5)] && ((reg841 ?
                              (8'h9e) : reg1271) ?
                          ((7'h42) >= reg521) : (^~reg470))) : $unsigned($unsigned($unsigned(wire1247)))),
                  (((!reg870) <= (~|$unsigned((8'hbc)))) ?
                      reg529[(2'h2):(2'h2)] : reg841)};
              reg1345 <= (^((7'h4c) || $unsigned(($unsigned((8'ha0)) ~^ $unsigned(reg894)))));
              reg1346 <= reg524;
              reg1347 = reg1294;
            end
          reg1348 = reg487;
        end
      reg1349 = ({$unsigned(($unsigned(reg498) ^~ $unsigned((8'hbd)))),
          (reg470[(3'h4):(2'h3)] ?
              $signed((reg1258 ?
                  reg877 : reg889)) : reg894[(4'hf):(4'h9)])} << (reg861[(3'h7):(1'h1)] ?
          reg469[(1'h0):(1'h0)] : $unsigned($unsigned($unsigned(reg1338)))));
      if ((8'hb1))
        begin
          reg1350 <= (~|(reg516[(5'h16):(4'hd)] << reg466[(3'h4):(2'h2)]));
        end
      else
        begin
          reg1351 = reg446;
          reg1352 <= $unsigned(((((reg898 | reg989) ?
                  $signed((7'h55)) : (&reg971)) ?
              (reg1350 ?
                  $signed(reg1348) : (reg469 ~^ reg536)) : ((^~reg498) * reg1331)) >= (((!wire438) ^~ reg524[(2'h3):(2'h3)]) ?
              reg968 : ((reg897 ? reg444 : reg514) ^ reg453[(3'h6):(1'h0)]))));
        end
      if ($unsigned($signed(reg1299)))
        begin
          for (forvar1353 = (1'h0); (forvar1353 < (1'h1)); forvar1353 = (forvar1353 + (1'h1)))
            begin
              reg1354 <= $unsigned(reg487[(2'h2):(1'h0)]);
              reg1355 <= (-$signed({(|$signed(reg1020)),
                  $signed((forvar1353 ? (7'h4c) : reg941))}));
              reg1356 <= ($unsigned((8'ha5)) * reg502);
            end
          reg1357 = reg1033;
          for (forvar1358 = (1'h0); (forvar1358 < (3'h5)); forvar1358 = (forvar1358 + (1'h1)))
            begin
              reg1359 = $unsigned(({((reg464 <= reg465) ^~ reg521[(1'h0):(1'h0)])} ?
                  ($unsigned($signed((7'h54))) ?
                      {reg891[(3'h5):(3'h4)],
                          reg511} : $unsigned($unsigned(reg990))) : $unsigned($unsigned(reg956))));
              reg1360 <= (!reg484[(4'h9):(2'h3)]);
              reg1361 <= wire437;
              reg1362 <= {{reg510[(5'h1c):(5'h11)], (^~$unsigned({reg1254}))}};
            end
          for (forvar1363 = (1'h0); (forvar1363 < (2'h2)); forvar1363 = (forvar1363 + (1'h1)))
            begin
              reg1364 = (((~^reg998[(4'h9):(3'h7)]) ?
                  wire860[(4'ha):(4'h9)] : (~&(reg514[(1'h1):(1'h1)] ?
                      reg444[(1'h1):(1'h0)] : reg868))) ^~ (~^reg521[(3'h6):(3'h5)]));
              reg1365 = reg1037[(3'h5):(3'h5)];
              reg1366 <= (((((forvar1328 - wire438) | reg1301[(3'h7):(3'h7)]) ?
                          reg503 : reg951) ?
                      reg524 : {$signed($unsigned((7'h54))),
                          $signed($unsigned(wire435))}) ?
                  (!(({reg867, (8'hba), reg1308} ?
                          $unsigned(reg878) : (^~reg1357)) ?
                      reg1264[(5'h17):(4'ha)] : (|(&reg484)))) : $signed($unsigned((reg894 ?
                      $signed((7'h52)) : (+reg523)))));
              reg1367 = {(~|reg847[(3'h7):(3'h7)]),
                  (!{reg1299,
                      $unsigned((reg509 ^~ reg877)),
                      forvar1343[(5'h15):(5'h10)]})};
              reg1368 <= (reg470[(2'h3):(1'h1)] ?
                  reg1290 : (~&$signed(reg897)));
              reg1369 <= {(&reg998[(4'h9):(3'h5)]),
                  $signed((wire1247[(3'h4):(2'h2)] ?
                      reg510[(2'h2):(1'h0)] : {(&reg1355),
                          $unsigned(reg1290),
                          reg1332})),
                  ($signed({$signed(reg1031),
                      (~|reg453),
                      reg916}) >> $signed(($unsigned(reg1328) >= reg1058[(1'h0):(1'h0)])))};
              reg1370 = ($signed($unsigned(reg1257[(1'h0):(1'h0)])) ?
                  (~$unsigned((reg1342[(1'h0):(1'h0)] ?
                      $signed(reg492) : {reg1360,
                          reg452,
                          reg489}))) : wire1059);
            end
          for (forvar1371 = (1'h0); (forvar1371 < (2'h2)); forvar1371 = (forvar1371 + (1'h1)))
            begin
              reg1372 <= $signed({(~reg1033)});
              reg1373 = (~reg929[(3'h5):(2'h3)]);
              reg1374 <= ($signed((reg465 ?
                  ($unsigned(reg1365) ?
                      $unsigned(reg473) : (reg997 >= reg870)) : {$unsigned(reg1342),
                      reg1299[(1'h0):(1'h0)],
                      reg517[(4'hc):(4'ha)]})) >> (&(reg452[(5'h12):(4'h9)] <<< reg1033)));
              reg1375 = $unsigned($signed(($signed(reg520[(5'h1a):(5'h14)]) && reg926)));
              reg1376 = reg507;
              reg1377 <= {($signed((reg1020[(3'h7):(1'h1)] ?
                      reg1292 : (reg465 && (8'hbd)))) > $unsigned(reg495)),
                  {(reg894 & $unsigned(((7'h44) ? (8'haf) : forvar1328)))},
                  (^({$unsigned(reg1352), (wire1247 ~^ reg1058)} != (|(reg507 ?
                      reg507 : (8'hb8)))))};
              reg1378 <= reg530;
            end
          reg1379 = $unsigned((8'hbb));
        end
      else
        begin
          if ((reg1338 ?
              reg1341 : (+{($unsigned(reg467) ? reg1372 : $signed(reg468))})))
            begin
              reg1353 <= (((&(~|reg970)) | (~^reg867[(5'h12):(1'h1)])) ?
                  reg1276[(3'h4):(2'h2)] : reg845[(3'h4):(2'h3)]);
              reg1354 <= (($signed($unsigned((8'hbc))) ?
                  $signed(((~&reg1379) && (reg870 ?
                      reg863 : (7'h46)))) : reg891) ~^ ({{{(8'ha9),
                              (8'ha0),
                              (8'haa)},
                          (8'hbc)}} ?
                  {reg1378, reg1307} : reg1278));
              reg1357 = $unsigned(reg1274);
              reg1358 = $unsigned(((^~(~^(reg1370 != reg907))) * (!reg1334[(3'h7):(3'h6)])));
              reg1360 <= $signed(($unsigned($signed($unsigned(reg537))) < reg840));
              reg1361 <= ($signed(reg1338) > {($signed($unsigned(reg443)) ?
                      $signed((~|reg520)) : ($unsigned(reg1306) ?
                          reg866[(4'ha):(4'h8)] : forvar1371)),
                  $unsigned(($signed(reg960) != (~|reg960)))});
              reg1362 <= $unsigned(reg1354[(3'h6):(3'h5)]);
            end
          else
            begin
              reg1357 = $unsigned({reg442});
              reg1358 = $signed((reg988[(4'h8):(1'h0)] ?
                  $signed(reg884[(2'h3):(1'h1)]) : ((forvar1358[(2'h3):(1'h0)] ?
                      reg864 : (reg1341 ?
                          reg1320 : reg1332)) && $signed(reg1370[(1'h0):(1'h0)]))));
              reg1360 <= $unsigned($signed((reg1370 - {{reg864,
                      reg1323,
                      reg891},
                  $unsigned(reg1264)})));
              reg1363 = reg1262[(5'h15):(4'hb)];
              reg1366 <= (~&$signed($unsigned((+$unsigned(reg909)))));
              reg1367 = ($signed(($signed($signed(reg461)) ?
                      $signed((reg1055 ? reg870 : reg1350)) : wire437)) ?
                  ($signed(((^~wire1246) <<< reg1310[(5'h1c):(5'h12)])) ?
                      (reg989[(5'h11):(3'h4)] == ((reg521 > reg951) ~^ $unsigned(reg1332))) : reg866) : $unsigned(reg1264));
            end
          reg1368 <= ($signed($signed(((reg1317 + reg532) - $signed(reg444)))) < $unsigned((7'h54)));
          reg1369 <= {{$unsigned(((^~(7'h50)) ?
                      $signed(reg537) : reg1359[(1'h1):(1'h0)])),
                  ((~|$unsigned(reg1260)) ?
                      {reg452} : $unsigned($signed((8'hac)))),
                  {((reg951 ~^ reg1051) >> (&reg941))}}};
          if ({$unsigned(reg489),
              ($signed((~&$unsigned(reg453))) >= (&$unsigned(reg480)))})
            begin
              reg1370 = ($signed($signed(((reg926 ? reg1022 : reg1329) ?
                  reg1313 : $signed(reg1340)))) | $signed((reg1379[(4'ha):(4'ha)] ^ {(reg951 ?
                      reg988 : reg1271),
                  ((8'h9e) | reg1375)})));
              reg1371 = reg1364;
              reg1373 = reg884[(4'h8):(3'h4)];
              reg1375 = (!(~&(-reg1295[(3'h5):(1'h1)])));
              reg1377 <= (reg1264 ?
                  $signed((~|(7'h46))) : reg1328[(5'h16):(5'h12)]);
            end
          else
            begin
              reg1372 <= (~reg919[(4'h9):(4'h9)]);
            end
          if ((|((8'hbf) ?
              (reg1363 ? reg1308 : ($unsigned(forvar1353) < reg476)) : reg845)))
            begin
              reg1378 <= (((!{(reg1352 << wire838),
                  (reg1031 == reg1278)}) >= ({(~|reg988),
                      ((8'hbc) <<< wire542),
                      $signed(reg1040)} ?
                  (reg995 != reg843) : (reg1330[(1'h1):(1'h0)] ?
                      {(7'h49), reg864} : (reg1049 ?
                          reg503 : reg1307)))) >>> $unsigned($signed(($unsigned(reg1051) ?
                  reg1378[(1'h0):(1'h0)] : reg509))));
              reg1379 = (7'h55);
            end
          else
            begin
              reg1379 = reg848[(1'h1):(1'h1)];
              reg1380 <= ({wire860} ?
                  reg1356[(4'h8):(2'h2)] : ((reg479 || {(+reg1033)}) ?
                      {(reg949[(2'h2):(1'h0)] >> $unsigned(reg1017)),
                          reg1335,
                          reg1055} : reg1355[(2'h2):(1'h0)]));
              reg1381 <= ({(^~$unsigned($signed(reg1328))),
                  ((~&reg1285) | ({reg926, reg511} ?
                      wire1247[(2'h3):(1'h0)] : $signed(reg1358)))} * $signed(({(&reg1332),
                  $signed(reg1283),
                  (reg1368 ? wire542 : reg1020)} >>> ($unsigned(reg916) ?
                  {(7'h52), (7'h51)} : ((7'h50) >>> reg1352)))));
              reg1382 = {reg1328, (!$signed($unsigned((reg1058 ~^ reg1294))))};
            end
          reg1383 = reg1017;
        end
      for (forvar1384 = (1'h0); (forvar1384 < (3'h5)); forvar1384 = (forvar1384 + (1'h1)))
        begin
          reg1385 = wire1247[(2'h3):(1'h0)];
          reg1386 <= (($signed($unsigned((7'h50))) ^~ reg1348) ?
              $signed((+reg1252[(4'hc):(4'hc)])) : (~&$signed($unsigned((forvar1371 < reg1041)))));
        end
    end
  module1387 #() modinst1479 (.clk(clk), .wire1390(reg533), .wire1391(reg1352), .wire1388(reg850), .wire1389(reg1257), .y(wire1478));
  module1480 #() modinst1991 (wire1990, clk, reg887, reg1283, reg883, reg1369);
  assign wire1992 = reg895;
  assign wire1993 = reg929;
  always
    @(posedge clk) begin
      reg1994 <= {($unsigned(reg514[(1'h0):(1'h0)]) ?
              (reg1319[(4'hb):(2'h3)] ?
                  reg850[(2'h3):(2'h3)] : reg487[(4'he):(4'hb)]) : wire438[(5'h12):(4'hb)])};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1480  (y, clk, wire1484, wire1483, wire1482, wire1481);
  output wire [(32'h20a6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire1484;
  input wire signed [(5'h1a):(1'h0)] wire1483;
  input wire [(5'h1b):(1'h0)] wire1482;
  input wire signed [(3'h4):(1'h0)] wire1481;
  wire [(3'h4):(1'h0)] wire1989;
  wire [(5'h11):(1'h0)] wire1988;
  wire [(5'h1f):(1'h0)] wire1987;
  wire signed [(2'h3):(1'h0)] wire1986;
  wire signed [(4'h8):(1'h0)] wire1985;
  wire [(4'hd):(1'h0)] wire1936;
  wire signed [(5'h13):(1'h0)] wire1836;
  wire [(5'h1b):(1'h0)] wire1835;
  wire signed [(5'h19):(1'h0)] wire1834;
  wire signed [(5'h1a):(1'h0)] wire1813;
  wire [(5'h15):(1'h0)] wire1812;
  wire [(2'h2):(1'h0)] wire1770;
  wire [(5'h12):(1'h0)] wire1769;
  wire signed [(5'h13):(1'h0)] wire1652;
  wire signed [(5'h1d):(1'h0)] wire1563;
  wire [(5'h1a):(1'h0)] wire1562;
  wire [(5'h1a):(1'h0)] wire1485;
  reg signed [(5'h11):(1'h0)] reg1984 = (1'h0);
  reg [(4'h8):(1'h0)] reg1983 = (1'h0);
  reg [(4'hb):(1'h0)] reg1980 = (1'h0);
  reg [(4'h9):(1'h0)] reg1979 = (1'h0);
  reg [(5'h15):(1'h0)] reg1978 = (1'h0);
  reg [(5'h19):(1'h0)] reg1977 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1976 = (1'h0);
  reg [(4'he):(1'h0)] reg1974 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1972 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1971 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1967 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1965 = (1'h0);
  reg [(5'h18):(1'h0)] reg1964 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1963 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1962 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1948 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1954 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1953 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1952 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1949 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1938 = (1'h0);
  reg [(5'h18):(1'h0)] reg1935 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1934 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1933 = (1'h0);
  reg [(5'h12):(1'h0)] reg1932 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1931 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1929 = (1'h0);
  reg [(5'h13):(1'h0)] reg1925 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1924 = (1'h0);
  reg [(4'hb):(1'h0)] reg1922 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1920 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1919 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1917 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1916 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1915 = (1'h0);
  reg [(5'h15):(1'h0)] reg1913 = (1'h0);
  reg [(3'h5):(1'h0)] reg1912 = (1'h0);
  reg [(4'ha):(1'h0)] reg1911 = (1'h0);
  reg [(5'h18):(1'h0)] reg1907 = (1'h0);
  reg [(4'ha):(1'h0)] reg1905 = (1'h0);
  reg [(2'h3):(1'h0)] reg1903 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1902 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1900 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1899 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1897 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1896 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1894 = (1'h0);
  reg [(3'h4):(1'h0)] reg1893 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1891 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1885 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1875 = (1'h0);
  reg [(5'h19):(1'h0)] reg1872 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1870 = (1'h0);
  reg [(4'ha):(1'h0)] reg1867 = (1'h0);
  reg [(4'hd):(1'h0)] reg1866 = (1'h0);
  reg [(3'h6):(1'h0)] reg1865 = (1'h0);
  reg [(5'h17):(1'h0)] reg1864 = (1'h0);
  reg [(2'h3):(1'h0)] reg1863 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1862 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1858 = (1'h0);
  reg [(5'h18):(1'h0)] reg1857 = (1'h0);
  reg [(4'hd):(1'h0)] reg1855 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1850 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1847 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1846 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1845 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1844 = (1'h0);
  reg [(5'h16):(1'h0)] reg1841 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1839 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1833 = (1'h0);
  reg [(3'h6):(1'h0)] reg1832 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1831 = (1'h0);
  reg [(5'h15):(1'h0)] reg1829 = (1'h0);
  reg [(5'h16):(1'h0)] reg1827 = (1'h0);
  reg [(5'h10):(1'h0)] reg1826 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1822 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1820 = (1'h0);
  reg [(4'ha):(1'h0)] reg1814 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1807 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1805 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1803 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1800 = (1'h0);
  reg [(5'h15):(1'h0)] reg1796 = (1'h0);
  reg [(5'h17):(1'h0)] reg1794 = (1'h0);
  reg [(4'hc):(1'h0)] reg1793 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1792 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1789 = (1'h0);
  reg [(4'hf):(1'h0)] reg1787 = (1'h0);
  reg [(4'h9):(1'h0)] reg1782 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1781 = (1'h0);
  reg [(3'h6):(1'h0)] reg1780 = (1'h0);
  reg [(5'h10):(1'h0)] reg1778 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1777 = (1'h0);
  reg [(5'h15):(1'h0)] reg1773 = (1'h0);
  reg [(5'h17):(1'h0)] reg1772 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1768 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1767 = (1'h0);
  reg [(4'h9):(1'h0)] reg1762 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1760 = (1'h0);
  reg [(5'h12):(1'h0)] reg1758 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1756 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1753 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1752 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1751 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1750 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1748 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1746 = (1'h0);
  reg [(2'h3):(1'h0)] reg1742 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1740 = (1'h0);
  reg [(5'h17):(1'h0)] reg1739 = (1'h0);
  reg [(4'h8):(1'h0)] reg1737 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1736 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1726 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1731 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1727 = (1'h0);
  reg [(5'h11):(1'h0)] reg1723 = (1'h0);
  reg [(4'ha):(1'h0)] reg1721 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1719 = (1'h0);
  reg [(3'h6):(1'h0)] reg1718 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1716 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1715 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1713 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1712 = (1'h0);
  reg [(3'h6):(1'h0)] reg1711 = (1'h0);
  reg [(5'h12):(1'h0)] reg1709 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1707 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1706 = (1'h0);
  reg [(5'h13):(1'h0)] reg1705 = (1'h0);
  reg [(5'h11):(1'h0)] reg1703 = (1'h0);
  reg [(5'h12):(1'h0)] reg1702 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1700 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1698 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1694 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1683 = (1'h0);
  reg [(5'h12):(1'h0)] reg1691 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1690 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1688 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1687 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1686 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1684 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1678 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1676 = (1'h0);
  reg [(5'h18):(1'h0)] reg1673 = (1'h0);
  reg [(3'h7):(1'h0)] reg1671 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1669 = (1'h0);
  reg [(5'h19):(1'h0)] reg1665 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1664 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1662 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1657 = (1'h0);
  reg [(2'h3):(1'h0)] reg1651 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1650 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1649 = (1'h0);
  reg [(2'h3):(1'h0)] reg1645 = (1'h0);
  reg [(5'h16):(1'h0)] reg1643 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1642 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1637 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1632 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1631 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1627 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1626 = (1'h0);
  reg [(3'h4):(1'h0)] reg1625 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1621 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1618 = (1'h0);
  reg [(5'h19):(1'h0)] reg1617 = (1'h0);
  reg [(3'h5):(1'h0)] reg1615 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1612 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1610 = (1'h0);
  reg [(4'ha):(1'h0)] reg1609 = (1'h0);
  reg [(4'hf):(1'h0)] reg1608 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1605 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1600 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1599 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1597 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1596 = (1'h0);
  reg [(2'h3):(1'h0)] reg1595 = (1'h0);
  reg [(4'h9):(1'h0)] reg1593 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1578 = (1'h0);
  reg [(5'h11):(1'h0)] reg1591 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1588 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1587 = (1'h0);
  reg [(5'h18):(1'h0)] reg1586 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1585 = (1'h0);
  reg [(2'h2):(1'h0)] reg1582 = (1'h0);
  reg [(5'h15):(1'h0)] reg1581 = (1'h0);
  reg [(5'h18):(1'h0)] reg1580 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1576 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1574 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1572 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1571 = (1'h0);
  reg [(5'h19):(1'h0)] reg1570 = (1'h0);
  reg [(2'h2):(1'h0)] reg1561 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1560 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1556 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1555 = (1'h0);
  reg [(5'h12):(1'h0)] reg1553 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1552 = (1'h0);
  reg [(4'h9):(1'h0)] reg1550 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1549 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1543 = (1'h0);
  reg [(4'h9):(1'h0)] reg1542 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1540 = (1'h0);
  reg [(5'h11):(1'h0)] reg1538 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1536 = (1'h0);
  reg [(3'h6):(1'h0)] reg1533 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1525 = (1'h0);
  reg [(4'ha):(1'h0)] reg1524 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1523 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1521 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1519 = (1'h0);
  reg [(5'h11):(1'h0)] reg1518 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1517 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1515 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1514 = (1'h0);
  reg [(4'h9):(1'h0)] reg1512 = (1'h0);
  reg [(3'h6):(1'h0)] reg1511 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1508 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1507 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1506 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1505 = (1'h0);
  reg [(2'h2):(1'h0)] reg1503 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1502 = (1'h0);
  reg [(5'h10):(1'h0)] reg1498 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1496 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1494 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1493 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1492 = (1'h0);
  reg [(5'h16):(1'h0)] reg1491 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1489 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1982 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1981 = (1'h0);
  reg [(3'h5):(1'h0)] reg1975 = (1'h0);
  reg [(4'hf):(1'h0)] reg1968 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1973 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1970 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1969 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1968 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1966 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1961 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1960 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1959 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1958 = (1'h0);
  reg [(2'h3):(1'h0)] reg1957 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1956 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1955 = (1'h0);
  reg [(5'h10):(1'h0)] reg1951 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1950 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1948 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1947 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1946 = (1'h0);
  reg [(2'h3):(1'h0)] reg1945 = (1'h0);
  reg [(4'hc):(1'h0)] reg1944 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1943 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1942 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1941 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1940 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1939 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1937 = (1'h0);
  reg [(5'h18):(1'h0)] reg1930 = (1'h0);
  reg [(4'h9):(1'h0)] reg1928 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1927 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1926 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1923 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1921 = (1'h0);
  reg [(3'h4):(1'h0)] reg1918 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1914 = (1'h0);
  reg [(5'h19):(1'h0)] reg1910 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1909 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1908 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1906 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1904 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1901 = (1'h0);
  reg [(3'h5):(1'h0)] reg1898 = (1'h0);
  reg [(3'h5):(1'h0)] reg1895 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1892 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1890 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1889 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1888 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1887 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1886 = (1'h0);
  reg [(2'h2):(1'h0)] reg1884 = (1'h0);
  reg [(5'h17):(1'h0)] reg1883 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1882 = (1'h0);
  reg [(3'h6):(1'h0)] reg1881 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1880 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar1879 = (1'h0);
  reg [(5'h15):(1'h0)] reg1878 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1877 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1876 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1874 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1873 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1859 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1871 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1869 = (1'h0);
  reg [(3'h6):(1'h0)] reg1868 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1861 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1860 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1859 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1856 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1854 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1853 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1852 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1851 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1849 = (1'h0);
  reg [(5'h13):(1'h0)] reg1848 = (1'h0);
  reg [(5'h17):(1'h0)] reg1843 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1842 = (1'h0);
  reg [(5'h15):(1'h0)] reg1840 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1838 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1837 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar1816 = (1'h0);
  reg [(4'hb):(1'h0)] reg1830 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1828 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1825 = (1'h0);
  reg [(3'h5):(1'h0)] reg1824 = (1'h0);
  reg [(3'h4):(1'h0)] reg1823 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1821 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1819 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1818 = (1'h0);
  reg [(5'h15):(1'h0)] reg1817 = (1'h0);
  reg [(5'h14):(1'h0)] reg1816 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1815 = (1'h0);
  reg [(5'h18):(1'h0)] reg1811 = (1'h0);
  reg [(5'h16):(1'h0)] reg1810 = (1'h0);
  reg [(5'h19):(1'h0)] reg1809 = (1'h0);
  reg [(5'h18):(1'h0)] reg1808 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1806 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1804 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1802 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1801 = (1'h0);
  reg [(2'h3):(1'h0)] reg1799 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1798 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1797 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1795 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1791 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar1790 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1788 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1786 = (1'h0);
  reg [(4'hc):(1'h0)] reg1785 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1784 = (1'h0);
  reg [(3'h4):(1'h0)] reg1783 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1779 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar1775 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1771 = (1'h0);
  reg [(4'he):(1'h0)] reg1779 = (1'h0);
  reg [(2'h2):(1'h0)] reg1776 = (1'h0);
  reg [(5'h11):(1'h0)] reg1775 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1774 = (1'h0);
  reg [(2'h2):(1'h0)] reg1771 = (1'h0);
  reg [(5'h15):(1'h0)] reg1766 = (1'h0);
  reg [(5'h11):(1'h0)] reg1765 = (1'h0);
  reg [(3'h7):(1'h0)] reg1764 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1763 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1760 = (1'h0);
  reg [(3'h6):(1'h0)] reg1761 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1759 = (1'h0);
  reg [(2'h2):(1'h0)] reg1757 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1755 = (1'h0);
  reg [(3'h4):(1'h0)] reg1754 = (1'h0);
  reg [(5'h13):(1'h0)] reg1749 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1747 = (1'h0);
  reg [(3'h4):(1'h0)] reg1745 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1744 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1743 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1741 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1738 = (1'h0);
  reg [(3'h4):(1'h0)] reg1735 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1734 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1733 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1721 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1732 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1730 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1729 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1728 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1726 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1725 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1724 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1722 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1720 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1717 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1714 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1710 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1708 = (1'h0);
  reg [(3'h6):(1'h0)] reg1704 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1701 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1699 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1697 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1696 = (1'h0);
  reg [(5'h14):(1'h0)] reg1695 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1693 = (1'h0);
  reg [(4'hc):(1'h0)] reg1692 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1689 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1685 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1683 = (1'h0);
  reg [(4'hf):(1'h0)] reg1682 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1681 = (1'h0);
  reg [(5'h17):(1'h0)] reg1680 = (1'h0);
  reg [(5'h16):(1'h0)] reg1679 = (1'h0);
  reg [(3'h4):(1'h0)] reg1677 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1675 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1674 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1672 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1670 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1668 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1667 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1666 = (1'h0);
  reg [(2'h2):(1'h0)] reg1663 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1661 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1660 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1659 = (1'h0);
  reg [(4'hf):(1'h0)] reg1658 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1656 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1655 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1654 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1653 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1648 = (1'h0);
  reg [(2'h3):(1'h0)] reg1647 = (1'h0);
  reg [(5'h13):(1'h0)] reg1646 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1643 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1644 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1641 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1640 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1639 = (1'h0);
  reg [(5'h12):(1'h0)] reg1638 = (1'h0);
  reg [(5'h11):(1'h0)] reg1636 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1635 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1634 = (1'h0);
  reg [(3'h4):(1'h0)] reg1633 = (1'h0);
  reg [(5'h12):(1'h0)] reg1630 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1629 = (1'h0);
  reg [(5'h19):(1'h0)] reg1628 = (1'h0);
  reg [(3'h7):(1'h0)] reg1624 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1623 = (1'h0);
  reg [(5'h11):(1'h0)] reg1622 = (1'h0);
  reg [(5'h10):(1'h0)] reg1620 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1619 = (1'h0);
  reg [(4'hf):(1'h0)] reg1616 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1614 = (1'h0);
  reg [(4'h8):(1'h0)] reg1613 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1611 = (1'h0);
  reg [(5'h19):(1'h0)] reg1607 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1606 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1604 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1603 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1602 = (1'h0);
  reg [(5'h19):(1'h0)] reg1601 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1598 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1594 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1592 = (1'h0);
  reg [(3'h5):(1'h0)] reg1590 = (1'h0);
  reg [(4'h9):(1'h0)] reg1589 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1584 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1583 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1579 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1578 = (1'h0);
  reg [(5'h14):(1'h0)] reg1577 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1575 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1573 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1569 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1568 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1567 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1566 = (1'h0);
  reg [(3'h5):(1'h0)] reg1565 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1564 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1559 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1558 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1557 = (1'h0);
  reg [(3'h5):(1'h0)] reg1554 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1551 = (1'h0);
  reg [(4'hf):(1'h0)] reg1548 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1547 = (1'h0);
  reg [(5'h13):(1'h0)] reg1546 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1545 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1544 = (1'h0);
  reg [(2'h2):(1'h0)] reg1541 = (1'h0);
  reg [(4'he):(1'h0)] forvar1539 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar1537 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1516 = (1'h0);
  reg [(5'h16):(1'h0)] reg1513 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1535 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1534 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1532 = (1'h0);
  reg [(2'h3):(1'h0)] reg1531 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1530 = (1'h0);
  reg [(5'h18):(1'h0)] reg1529 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1528 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1527 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1526 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1522 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1520 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1516 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1513 = (1'h0);
  reg [(3'h7):(1'h0)] reg1510 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1509 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1504 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1501 = (1'h0);
  reg [(5'h10):(1'h0)] reg1500 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1499 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1497 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1488 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1486 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1495 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1490 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1488 = (1'h0);
  reg [(2'h2):(1'h0)] reg1487 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1486 = (1'h0);
  assign y = {wire1989,
                 wire1988,
                 wire1987,
                 wire1986,
                 wire1985,
                 wire1936,
                 wire1836,
                 wire1835,
                 wire1834,
                 wire1813,
                 wire1812,
                 wire1770,
                 wire1769,
                 wire1652,
                 wire1563,
                 wire1562,
                 wire1485,
                 reg1984,
                 reg1983,
                 reg1980,
                 reg1979,
                 reg1978,
                 reg1977,
                 reg1976,
                 reg1974,
                 reg1972,
                 reg1971,
                 reg1967,
                 reg1965,
                 reg1964,
                 reg1963,
                 reg1962,
                 reg1948,
                 reg1954,
                 reg1953,
                 reg1952,
                 reg1949,
                 reg1938,
                 reg1935,
                 reg1934,
                 reg1933,
                 reg1932,
                 reg1931,
                 reg1929,
                 reg1925,
                 reg1924,
                 reg1922,
                 reg1920,
                 reg1919,
                 reg1917,
                 reg1916,
                 reg1915,
                 reg1913,
                 reg1912,
                 reg1911,
                 reg1907,
                 reg1905,
                 reg1903,
                 reg1902,
                 reg1900,
                 reg1899,
                 reg1897,
                 reg1896,
                 reg1894,
                 reg1893,
                 reg1891,
                 reg1885,
                 reg1875,
                 reg1872,
                 reg1870,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1864,
                 reg1863,
                 reg1862,
                 reg1858,
                 reg1857,
                 reg1855,
                 reg1850,
                 reg1847,
                 reg1846,
                 reg1845,
                 reg1844,
                 reg1841,
                 reg1839,
                 reg1833,
                 reg1832,
                 reg1831,
                 reg1829,
                 reg1827,
                 reg1826,
                 reg1822,
                 reg1820,
                 reg1814,
                 reg1807,
                 reg1805,
                 reg1803,
                 reg1800,
                 reg1796,
                 reg1794,
                 reg1793,
                 reg1792,
                 reg1789,
                 reg1787,
                 reg1782,
                 reg1781,
                 reg1780,
                 reg1778,
                 reg1777,
                 reg1773,
                 reg1772,
                 reg1768,
                 reg1767,
                 reg1762,
                 reg1760,
                 reg1758,
                 reg1756,
                 reg1753,
                 reg1752,
                 reg1751,
                 reg1750,
                 reg1748,
                 reg1746,
                 reg1742,
                 reg1740,
                 reg1739,
                 reg1737,
                 reg1736,
                 reg1726,
                 reg1731,
                 reg1727,
                 reg1723,
                 reg1721,
                 reg1719,
                 reg1718,
                 reg1716,
                 reg1715,
                 reg1713,
                 reg1712,
                 reg1711,
                 reg1709,
                 reg1707,
                 reg1706,
                 reg1705,
                 reg1703,
                 reg1702,
                 reg1700,
                 reg1698,
                 reg1694,
                 reg1683,
                 reg1691,
                 reg1690,
                 reg1688,
                 reg1687,
                 reg1686,
                 reg1684,
                 reg1678,
                 reg1676,
                 reg1673,
                 reg1671,
                 reg1669,
                 reg1665,
                 reg1664,
                 reg1662,
                 reg1657,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1645,
                 reg1643,
                 reg1642,
                 reg1637,
                 reg1632,
                 reg1631,
                 reg1627,
                 reg1626,
                 reg1625,
                 reg1621,
                 reg1618,
                 reg1617,
                 reg1615,
                 reg1612,
                 reg1610,
                 reg1609,
                 reg1608,
                 reg1605,
                 reg1600,
                 reg1599,
                 reg1597,
                 reg1596,
                 reg1595,
                 reg1593,
                 reg1578,
                 reg1591,
                 reg1588,
                 reg1587,
                 reg1586,
                 reg1585,
                 reg1582,
                 reg1581,
                 reg1580,
                 reg1576,
                 reg1574,
                 reg1572,
                 reg1571,
                 reg1570,
                 reg1561,
                 reg1560,
                 reg1556,
                 reg1555,
                 reg1553,
                 reg1552,
                 reg1550,
                 reg1549,
                 reg1543,
                 reg1542,
                 reg1540,
                 reg1538,
                 reg1536,
                 reg1533,
                 reg1525,
                 reg1524,
                 reg1523,
                 reg1521,
                 reg1519,
                 reg1518,
                 reg1517,
                 reg1515,
                 reg1514,
                 reg1512,
                 reg1511,
                 reg1508,
                 reg1507,
                 reg1506,
                 reg1505,
                 reg1503,
                 reg1502,
                 reg1498,
                 reg1496,
                 reg1494,
                 reg1493,
                 reg1492,
                 reg1491,
                 reg1489,
                 reg1982,
                 reg1981,
                 reg1975,
                 reg1968,
                 reg1973,
                 reg1970,
                 reg1969,
                 forvar1968,
                 reg1966,
                 forvar1961,
                 reg1960,
                 forvar1959,
                 forvar1958,
                 reg1957,
                 reg1956,
                 reg1955,
                 reg1951,
                 reg1950,
                 forvar1948,
                 reg1947,
                 reg1946,
                 reg1945,
                 reg1944,
                 reg1943,
                 reg1942,
                 reg1941,
                 forvar1940,
                 reg1939,
                 forvar1937,
                 reg1930,
                 reg1928,
                 forvar1927,
                 reg1926,
                 reg1923,
                 forvar1921,
                 reg1918,
                 reg1914,
                 reg1910,
                 reg1909,
                 reg1908,
                 reg1906,
                 reg1904,
                 forvar1901,
                 reg1898,
                 reg1895,
                 forvar1892,
                 forvar1890,
                 forvar1889,
                 reg1888,
                 reg1887,
                 reg1886,
                 reg1884,
                 reg1883,
                 reg1882,
                 reg1881,
                 forvar1880,
                 forvar1879,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1874,
                 reg1873,
                 forvar1859,
                 reg1871,
                 forvar1869,
                 reg1868,
                 reg1861,
                 reg1860,
                 reg1859,
                 reg1856,
                 reg1854,
                 reg1853,
                 reg1852,
                 forvar1851,
                 forvar1849,
                 reg1848,
                 reg1843,
                 reg1842,
                 reg1840,
                 reg1838,
                 forvar1837,
                 forvar1816,
                 reg1830,
                 reg1828,
                 forvar1825,
                 reg1824,
                 reg1823,
                 reg1821,
                 reg1819,
                 reg1818,
                 reg1817,
                 reg1816,
                 reg1815,
                 reg1811,
                 reg1810,
                 reg1809,
                 reg1808,
                 reg1806,
                 forvar1804,
                 reg1802,
                 reg1801,
                 reg1799,
                 reg1798,
                 reg1797,
                 reg1795,
                 forvar1791,
                 forvar1790,
                 reg1788,
                 reg1786,
                 reg1785,
                 reg1784,
                 reg1783,
                 forvar1779,
                 forvar1775,
                 forvar1771,
                 reg1779,
                 reg1776,
                 reg1775,
                 reg1774,
                 reg1771,
                 reg1766,
                 reg1765,
                 reg1764,
                 reg1763,
                 forvar1760,
                 reg1761,
                 reg1759,
                 reg1757,
                 reg1755,
                 reg1754,
                 reg1749,
                 reg1747,
                 reg1745,
                 reg1744,
                 reg1743,
                 reg1741,
                 reg1738,
                 reg1735,
                 reg1734,
                 forvar1733,
                 forvar1721,
                 reg1732,
                 forvar1730,
                 reg1729,
                 reg1728,
                 forvar1726,
                 reg1725,
                 reg1724,
                 reg1722,
                 reg1720,
                 reg1717,
                 reg1714,
                 reg1710,
                 reg1708,
                 reg1704,
                 reg1701,
                 forvar1699,
                 reg1697,
                 reg1696,
                 reg1695,
                 forvar1693,
                 reg1692,
                 reg1689,
                 reg1685,
                 forvar1683,
                 reg1682,
                 reg1681,
                 reg1680,
                 reg1679,
                 reg1677,
                 reg1675,
                 reg1674,
                 forvar1672,
                 reg1670,
                 reg1668,
                 reg1667,
                 reg1666,
                 reg1663,
                 reg1661,
                 forvar1660,
                 reg1659,
                 reg1658,
                 reg1656,
                 reg1655,
                 reg1654,
                 forvar1653,
                 reg1648,
                 reg1647,
                 reg1646,
                 forvar1643,
                 reg1644,
                 reg1641,
                 reg1640,
                 reg1639,
                 reg1638,
                 reg1636,
                 reg1635,
                 reg1634,
                 reg1633,
                 reg1630,
                 reg1629,
                 reg1628,
                 reg1624,
                 forvar1623,
                 reg1622,
                 reg1620,
                 reg1619,
                 reg1616,
                 reg1614,
                 reg1613,
                 reg1611,
                 reg1607,
                 reg1606,
                 reg1604,
                 forvar1603,
                 reg1602,
                 reg1601,
                 reg1598,
                 reg1594,
                 reg1592,
                 reg1590,
                 reg1589,
                 reg1584,
                 reg1583,
                 reg1579,
                 forvar1578,
                 reg1577,
                 reg1575,
                 reg1573,
                 reg1569,
                 forvar1568,
                 reg1567,
                 forvar1566,
                 reg1565,
                 forvar1564,
                 reg1559,
                 reg1558,
                 reg1557,
                 reg1554,
                 reg1551,
                 reg1548,
                 reg1547,
                 reg1546,
                 reg1545,
                 reg1544,
                 reg1541,
                 forvar1539,
                 forvar1537,
                 reg1516,
                 reg1513,
                 reg1535,
                 reg1534,
                 reg1532,
                 reg1531,
                 forvar1530,
                 reg1529,
                 reg1528,
                 reg1527,
                 reg1526,
                 reg1522,
                 reg1520,
                 forvar1516,
                 forvar1513,
                 reg1510,
                 reg1509,
                 reg1504,
                 reg1501,
                 reg1500,
                 forvar1499,
                 forvar1497,
                 reg1488,
                 forvar1486,
                 reg1495,
                 reg1490,
                 forvar1488,
                 reg1487,
                 reg1486,
                 (1'h0)};
  assign wire1485 = wire1483[(2'h3):(1'h1)];
  always
    @(posedge clk) begin
      if (($signed($unsigned($signed(wire1484))) & $signed((((wire1482 ?
                  (7'h43) : wire1484) ?
              $signed(wire1481) : $signed(wire1483)) ?
          (8'h9c) : (&wire1483)))))
        begin
          reg1486 = {$signed($signed({(+wire1485)}))};
          reg1487 = (($signed(((-wire1485) ^~ (wire1485 ?
                  wire1482 : wire1482))) | $signed($unsigned($unsigned(reg1486)))) ?
              wire1484 : ($unsigned($unsigned((wire1485 ? reg1486 : (7'h56)))) ?
                  (|(^~wire1481)) : ($unsigned((8'ha1)) || (-reg1486))));
          for (forvar1488 = (1'h0); (forvar1488 < (3'h4)); forvar1488 = (forvar1488 + (1'h1)))
            begin
              reg1489 <= $unsigned(wire1484);
              reg1490 = ((~&wire1484[(1'h0):(1'h0)]) ?
                  (7'h4e) : wire1482[(4'hd):(3'h7)]);
              reg1491 <= $unsigned(({(~&(wire1485 + reg1487)),
                  {(~|reg1489), $unsigned(reg1490), wire1482},
                  (~&(wire1485 ?
                      wire1485 : wire1481))} <<< {{((8'hac) != (8'ha2)),
                      $signed(wire1485)},
                  ($signed(reg1487) <<< (reg1486 ? wire1484 : reg1487)),
                  ((7'h45) || $signed(reg1487))}));
              reg1492 <= $signed(wire1483);
              reg1493 <= reg1487;
              reg1494 <= (&($unsigned(reg1491) ?
                  forvar1488 : (wire1485[(5'h19):(4'hd)] < reg1486)));
              reg1495 = reg1487;
            end
        end
      else
        begin
          for (forvar1486 = (1'h0); (forvar1486 < (2'h3)); forvar1486 = (forvar1486 + (1'h1)))
            begin
              reg1487 = $unsigned((-$unsigned($signed((~|forvar1488)))));
              reg1488 = $signed($unsigned({(wire1481[(2'h2):(1'h0)] ?
                      $unsigned(forvar1488) : $unsigned((8'h9e)))}));
              reg1489 <= ((wire1484[(1'h1):(1'h1)] ?
                      $unsigned({{wire1485, reg1493},
                          reg1489}) : ((^~$signed(wire1484)) ?
                          $unsigned((8'ha5)) : (forvar1488[(3'h7):(2'h2)] ^~ wire1484[(2'h2):(2'h2)]))) ?
                  (~^$unsigned({$signed((8'ha0))})) : $signed(($signed(reg1492[(3'h7):(2'h2)]) ?
                      $unsigned(reg1492) : reg1495[(2'h2):(2'h2)])));
              reg1491 <= (&(((7'h4c) >>> $signed((wire1482 ?
                      reg1487 : forvar1488))) ?
                  wire1483[(3'h4):(1'h0)] : wire1485[(4'hd):(1'h1)]));
            end
        end
      reg1496 <= wire1484[(2'h2):(2'h2)];
      for (forvar1497 = (1'h0); (forvar1497 < (1'h0)); forvar1497 = (forvar1497 + (1'h1)))
        begin
          reg1498 <= reg1492;
          for (forvar1499 = (1'h0); (forvar1499 < (1'h1)); forvar1499 = (forvar1499 + (1'h1)))
            begin
              reg1500 = ($unsigned(({wire1482,
                      $unsigned(reg1488)} && $signed($signed(forvar1499)))) ?
                  ({reg1489} ?
                      wire1485[(3'h4):(1'h0)] : forvar1486[(3'h7):(3'h5)]) : ((~&wire1481) ?
                      (^$signed((wire1484 ?
                          reg1498 : forvar1486))) : (!(^~(8'hab)))));
            end
          reg1501 = $signed({reg1487,
              (wire1485 ?
                  reg1491 : (forvar1499 ?
                      $unsigned(wire1483) : $signed((8'hb0))))});
          if ({$signed((($signed(forvar1499) ?
                  $unsigned(forvar1486) : reg1496[(4'h8):(3'h5)]) < ($unsigned(reg1488) ?
                  (forvar1499 < forvar1497) : (reg1490 ?
                      (8'h9e) : wire1483))))})
            begin
              reg1502 <= reg1496;
              reg1503 <= {forvar1497[(3'h5):(3'h4)],
                  (~&wire1485),
                  wire1484[(1'h0):(1'h0)]};
              reg1504 = (8'hb2);
              reg1505 <= (reg1489[(3'h4):(2'h3)] ?
                  wire1485[(1'h0):(1'h0)] : reg1493);
              reg1506 <= $unsigned({((~&(^forvar1499)) >> (~^(-reg1502))),
                  forvar1488[(3'h5):(1'h0)]});
            end
          else
            begin
              reg1502 <= $signed($unsigned($unsigned({$unsigned(reg1490),
                  $signed(wire1482)})));
              reg1503 <= wire1481;
              reg1504 = reg1492;
              reg1505 <= (forvar1488[(1'h0):(1'h0)] ^~ reg1494[(5'h14):(4'ha)]);
            end
          reg1507 <= $unsigned(($signed($unsigned($signed(reg1492))) <= {(forvar1486[(4'h9):(4'h8)] ?
                  (reg1504 ? reg1488 : reg1505) : {reg1493, reg1503}),
              $unsigned($signed(reg1505)),
              reg1493}));
          reg1508 <= reg1503;
          if (reg1491[(3'h4):(2'h2)])
            begin
              reg1509 = (-$unsigned(wire1485));
              reg1510 = reg1500;
            end
          else
            begin
              reg1511 <= $unsigned($unsigned((8'hab)));
              reg1512 <= (reg1498 - wire1481);
            end
        end
      if (reg1506[(5'h15):(4'ha)])
        begin
          for (forvar1513 = (1'h0); (forvar1513 < (3'h6)); forvar1513 = (forvar1513 + (1'h1)))
            begin
              reg1514 <= (&(forvar1499[(1'h1):(1'h0)] * (+(8'ha1))));
              reg1515 <= $unsigned({$unsigned((-reg1506[(4'ha):(2'h2)]))});
            end
          for (forvar1516 = (1'h0); (forvar1516 < (1'h1)); forvar1516 = (forvar1516 + (1'h1)))
            begin
              reg1517 <= reg1487[(2'h2):(2'h2)];
              reg1518 <= reg1498[(4'hf):(3'h6)];
              reg1519 <= (reg1498[(3'h7):(3'h6)] ?
                  reg1494 : $signed(({(&reg1500),
                          reg1514[(5'h1a):(5'h12)],
                          (reg1509 | reg1504)} ?
                      $signed($unsigned(reg1509)) : $unsigned((reg1518 ?
                          reg1507 : wire1484)))));
              reg1520 = (((~&(!(|reg1491))) ?
                      ($signed($unsigned(forvar1499)) << (8'hbf)) : {(|reg1509[(5'h12):(4'hd)]),
                          (~&(~wire1484))}) ?
                  {$signed((wire1484 >= (reg1488 ?
                          reg1496 : reg1514)))} : (~|((~((8'hb1) >> (8'ha8))) << reg1512[(2'h3):(1'h1)])));
              reg1521 <= (reg1491[(2'h2):(2'h2)] - {(reg1509 ?
                      reg1520[(2'h3):(2'h3)] : reg1515)});
              reg1522 = reg1506;
              reg1523 <= (!reg1491);
            end
          if ($signed(reg1495[(1'h0):(1'h0)]))
            begin
              reg1524 <= wire1484[(2'h2):(1'h1)];
              reg1525 <= {$unsigned(($signed($signed(reg1522)) ?
                      ((reg1511 & forvar1488) - (forvar1499 ?
                          (8'h9d) : reg1509)) : forvar1499[(1'h0):(1'h0)])),
                  (($unsigned((|reg1514)) == reg1523) < $signed(($unsigned(reg1508) ?
                      $unsigned(reg1507) : reg1500[(4'he):(3'h7)])))};
            end
          else
            begin
              reg1526 = reg1495[(4'hb):(1'h0)];
              reg1527 = (forvar1516 ?
                  forvar1499[(2'h3):(2'h3)] : (reg1493 && $unsigned(reg1511)));
              reg1528 = $signed(($signed($signed($unsigned(reg1490))) ?
                  reg1488[(4'h8):(3'h5)] : ((~^{reg1489, forvar1513}) ?
                      ((reg1493 ? reg1511 : wire1482) ~^ ((8'ha8) ?
                          reg1487 : reg1512)) : (&reg1517[(1'h0):(1'h0)]))));
            end
          reg1529 = {reg1508,
              (~^(wire1483 ?
                  ((forvar1513 ? wire1481 : reg1527) ?
                      reg1501[(4'h8):(3'h7)] : reg1490) : ((~&reg1510) ?
                      reg1491 : {reg1502, (8'hba), forvar1488})))};
          for (forvar1530 = (1'h0); (forvar1530 < (3'h5)); forvar1530 = (forvar1530 + (1'h1)))
            begin
              reg1531 = (&(((~&{reg1527}) ?
                      reg1488[(3'h5):(3'h5)] : {reg1498, $unsigned((7'h51))}) ?
                  {reg1490} : ((~^wire1481) ?
                      reg1496[(4'hb):(2'h2)] : ($unsigned(reg1490) ?
                          reg1522 : (forvar1488 ? reg1517 : reg1501)))));
              reg1532 = $unsigned(reg1506);
              reg1533 <= (~&(reg1493[(5'h12):(5'h11)] && (8'ha3)));
              reg1534 = ((&forvar1516) ?
                  $signed($unsigned($signed({reg1521,
                      reg1494}))) : $signed((~reg1509)));
              reg1535 = $unsigned((^$signed(wire1483)));
              reg1536 <= $unsigned({(reg1522 + reg1522), $unsigned((8'hb2))});
            end
        end
      else
        begin
          if ((reg1495 ?
              (($unsigned(wire1484) != reg1528[(3'h5):(3'h4)]) ^~ forvar1499) : (+reg1531[(1'h1):(1'h1)])))
            begin
              reg1513 = (~reg1524[(2'h2):(1'h0)]);
              reg1514 <= (((~&$unsigned($unsigned((7'h57)))) ?
                      {$unsigned(reg1534),
                          ((reg1512 & forvar1488) << ((8'ha8) ?
                              reg1531 : wire1482)),
                          ($signed(reg1524) ?
                              $signed(reg1527) : (~&forvar1497))} : forvar1488) ?
                  $unsigned((^~$unsigned($unsigned(reg1488)))) : forvar1488[(3'h4):(1'h0)]);
              reg1516 = (+$signed(reg1512[(4'h8):(2'h3)]));
              reg1520 = reg1536[(1'h0):(1'h0)];
              reg1522 = reg1520;
              reg1523 <= ((reg1486 ?
                      $signed((wire1483[(5'h19):(5'h12)] << reg1500[(3'h6):(3'h6)])) : reg1510[(3'h7):(3'h4)]) ?
                  reg1511[(1'h1):(1'h1)] : $unsigned((reg1534 <<< ({forvar1516,
                      reg1488,
                      (8'hbd)} + $signed(reg1535)))));
            end
          else
            begin
              reg1513 = reg1517;
              reg1516 = reg1518[(4'hf):(4'he)];
              reg1520 = (8'hbc);
            end
          reg1526 = reg1516;
        end
      for (forvar1537 = (1'h0); (forvar1537 < (1'h0)); forvar1537 = (forvar1537 + (1'h1)))
        begin
          reg1538 <= reg1510[(1'h0):(1'h0)];
          for (forvar1539 = (1'h0); (forvar1539 < (2'h3)); forvar1539 = (forvar1539 + (1'h1)))
            begin
              reg1540 <= $signed(((reg1510 ?
                      $signed((reg1508 || forvar1488)) : reg1538[(4'h9):(3'h4)]) ?
                  $signed(wire1483) : $signed(((+reg1509) ~^ $signed(reg1505)))));
              reg1541 = $unsigned(($signed((reg1517[(3'h5):(2'h2)] - (8'hac))) >> ($signed($signed(forvar1539)) * {$unsigned((8'had)),
                  forvar1497[(4'hd):(2'h2)]})));
              reg1542 <= $unsigned(($signed(((reg1536 >> reg1495) & $unsigned(reg1511))) << forvar1497[(4'hd):(4'hc)]));
              reg1543 <= (&$unsigned(({wire1485, reg1536, $signed(reg1506)} ?
                  ($signed((8'hbc)) || reg1524[(3'h5):(1'h0)]) : $signed($signed((8'hb3))))));
              reg1544 = reg1541[(1'h1):(1'h0)];
              reg1545 = $unsigned((7'h40));
              reg1546 = $unsigned(reg1534);
            end
          if (forvar1537)
            begin
              reg1547 = reg1519;
              reg1548 = {({$signed(reg1488[(3'h6):(2'h2)]), reg1543} ?
                      (reg1509 ?
                          $signed((reg1546 <<< reg1517)) : reg1531) : $unsigned(((reg1503 | reg1504) ?
                          (reg1498 ? forvar1513 : reg1547) : reg1540))),
                  reg1528};
              reg1549 <= reg1504[(4'hd):(1'h1)];
              reg1550 <= ((-($signed(reg1511[(3'h6):(3'h6)]) ?
                      wire1481[(2'h3):(1'h0)] : ((reg1549 ?
                          reg1549 : forvar1516) >= (-forvar1486)))) ?
                  ((-$unsigned({reg1487,
                      reg1540})) > (reg1538[(3'h5):(1'h0)] | reg1527[(3'h6):(3'h5)])) : (($unsigned($signed(reg1531)) ?
                          $signed({reg1491, wire1483}) : reg1536) ?
                      reg1509[(4'h9):(3'h7)] : reg1495[(1'h1):(1'h1)]));
            end
          else
            begin
              reg1549 <= ({reg1487[(1'h0):(1'h0)],
                      (forvar1516[(2'h3):(1'h0)] ^~ {$unsigned(reg1543)})} ?
                  $signed($unsigned((forvar1486 ?
                      reg1514[(1'h1):(1'h0)] : (reg1540 ?
                          reg1523 : reg1495)))) : ((((reg1502 ?
                              (8'hb9) : (7'h54)) ?
                          (reg1491 ? reg1487 : reg1512) : (reg1516 | reg1516)) ?
                      reg1486[(4'hd):(4'h8)] : {(reg1517 ? reg1506 : reg1488),
                          $unsigned(reg1526),
                          (&reg1542)}) || reg1534));
              reg1550 <= $unsigned($signed(forvar1539));
              reg1551 = ($signed($signed(reg1543[(4'hd):(2'h3)])) ?
                  reg1512 : reg1511);
              reg1552 <= $unsigned($unsigned(reg1541));
              reg1553 <= $signed((^{reg1543, (~^(^~wire1481))}));
              reg1554 = reg1550[(2'h3):(1'h1)];
              reg1555 <= forvar1486[(5'h17):(4'ha)];
            end
          if (reg1554[(3'h4):(1'h0)])
            begin
              reg1556 <= wire1483[(2'h2):(1'h0)];
              reg1557 = forvar1486[(4'h8):(3'h6)];
              reg1558 = (~{$unsigned(($signed(reg1504) ?
                      (-reg1525) : $unsigned(forvar1488)))});
              reg1559 = (reg1487 >> $unsigned(reg1511));
            end
          else
            begin
              reg1556 <= (reg1488[(1'h1):(1'h0)] ?
                  {(({(8'h9e)} ?
                          $signed(reg1496) : ((8'hb6) || reg1556)) >= reg1505)} : $unsigned(reg1534));
              reg1557 = (-(reg1526 ?
                  $unsigned((reg1534[(3'h6):(2'h3)] ?
                      (forvar1488 ?
                          reg1517 : reg1509) : reg1516)) : ($signed({wire1485}) < (wire1485 && $unsigned((8'ha6))))));
              reg1558 = reg1513[(5'h10):(4'he)];
              reg1559 = $unsigned((-((((8'hbf) ?
                  reg1551 : reg1504) ^~ (reg1513 >= reg1553)) >>> reg1559)));
              reg1560 <= {($signed($signed({wire1485, (8'ha7)})) ?
                      (+{(reg1543 > reg1526),
                          (reg1554 ? reg1489 : forvar1486),
                          (+wire1483)}) : ($signed((^~forvar1499)) ?
                          {{reg1492, reg1519, reg1486}} : reg1545))};
            end
          reg1561 <= $unsigned(reg1502);
        end
    end
  assign wire1562 = (&($unsigned(((reg1493 <<< reg1493) ?
                        $signed(reg1549) : $signed(reg1489))) && (((reg1515 ?
                            reg1538 : reg1512) == wire1485) ?
                        ({reg1519} >>> {reg1533,
                            (8'hb2),
                            reg1506}) : $signed(reg1533))));
  assign wire1563 = ($unsigned((&$signed(((8'hb0) & reg1506)))) ~^ reg1493);
  always
    @(posedge clk) begin
      for (forvar1564 = (1'h0); (forvar1564 < (1'h1)); forvar1564 = (forvar1564 + (1'h1)))
        begin
          reg1565 = $unsigned(reg1517[(1'h1):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar1566 = (1'h0); (forvar1566 < (3'h5)); forvar1566 = (forvar1566 + (1'h1)))
        begin
          reg1567 = (~|(reg1538 ?
              (~reg1514) : ({reg1521,
                  (reg1494 ? reg1552 : (7'h4c))} ~^ wire1562)));
          for (forvar1568 = (1'h0); (forvar1568 < (2'h3)); forvar1568 = (forvar1568 + (1'h1)))
            begin
              reg1569 = $signed({reg1512[(2'h2):(1'h0)],
                  reg1505[(5'h1a):(5'h10)]});
              reg1570 <= reg1519;
              reg1571 <= $unsigned((((-reg1553[(4'ha):(1'h0)]) * {{wire1481,
                          reg1549}}) ?
                  {reg1502[(4'he):(4'hc)],
                      reg1494,
                      ($unsigned((8'hac)) ~^ (!(8'h9f)))} : reg1525));
              reg1572 <= $unsigned((!$signed((reg1493 ?
                  (&reg1569) : (reg1550 * wire1481)))));
            end
          reg1573 = reg1570;
          reg1574 <= $unsigned(reg1502[(4'hc):(4'hc)]);
          reg1575 = $signed((reg1538 ?
              reg1519[(4'ha):(4'ha)] : $unsigned(($signed((8'hbe)) ?
                  (&reg1514) : reg1521[(3'h4):(3'h4)]))));
          reg1576 <= $unsigned((|((^~$signed(reg1560)) < reg1508[(5'h16):(4'he)])));
        end
      reg1577 = (&(^~$signed((reg1525 ?
          {reg1525, reg1524, wire1563} : $signed(reg1569)))));
      if (({reg1555,
              $signed($unsigned({reg1493, reg1561})),
              (($unsigned(reg1533) | $unsigned(wire1563)) <= $signed({reg1492,
                  (8'ha5),
                  reg1567}))} ?
          $unsigned((forvar1566[(3'h4):(2'h2)] >>> wire1562)) : (-((~$unsigned(reg1512)) ?
              $unsigned((reg1523 ? (8'hbc) : wire1482)) : $signed({wire1563,
                  reg1507,
                  reg1515})))))
        begin
          for (forvar1578 = (1'h0); (forvar1578 < (3'h4)); forvar1578 = (forvar1578 + (1'h1)))
            begin
              reg1579 = reg1536;
              reg1580 <= {(~&$signed((7'h52))),
                  $unsigned(reg1489),
                  (reg1493 ?
                      ($unsigned((&reg1540)) ?
                          (reg1493[(5'h13):(3'h6)] <<< (reg1540 ?
                              reg1553 : reg1538)) : {$signed(reg1571),
                              forvar1568,
                              reg1507[(1'h0):(1'h0)]}) : wire1481)};
              reg1581 <= (7'h54);
            end
          if ((reg1506 + $unsigned(forvar1568)))
            begin
              reg1582 <= ((~|$unsigned(reg1498[(2'h3):(2'h2)])) ?
                  $unsigned(((reg1579[(2'h3):(2'h3)] || forvar1578[(3'h4):(1'h1)]) != (~^reg1498[(2'h2):(1'h1)]))) : (&{$signed({reg1505,
                          wire1482})}));
            end
          else
            begin
              reg1583 = (~wire1484);
              reg1584 = $unsigned($unsigned(wire1484[(2'h2):(2'h2)]));
              reg1585 <= $unsigned((reg1582[(1'h0):(1'h0)] == (reg1508[(1'h0):(1'h0)] < (((8'hba) ?
                  wire1481 : reg1540) >> reg1491))));
            end
          reg1586 <= (({reg1584,
                      (reg1585[(4'ha):(3'h7)] > (reg1517 ? (8'hb6) : reg1493)),
                      (~^{reg1571})} ?
                  reg1571 : $unsigned({reg1560[(3'h5):(2'h3)],
                      ((8'ha7) || reg1521)})) ?
              reg1533[(2'h2):(2'h2)] : (7'h58));
          if ($signed($unsigned(((-(reg1560 ? reg1498 : reg1540)) ?
              ($unsigned(wire1562) ^ $unsigned((7'h56))) : (reg1511 ?
                  (~&reg1552) : $unsigned(reg1572))))))
            begin
              reg1587 <= ($unsigned((reg1525[(2'h2):(2'h2)] - wire1483[(5'h10):(2'h3)])) | (reg1579[(1'h0):(1'h0)] ?
                  reg1508[(5'h14):(1'h0)] : reg1518[(4'hf):(2'h2)]));
              reg1588 <= $unsigned((forvar1568[(3'h5):(1'h0)] ?
                  $unsigned((~(reg1494 ?
                      reg1508 : reg1549))) : (~(reg1555[(4'ha):(1'h1)] * (reg1543 ?
                      reg1582 : reg1508)))));
              reg1589 = reg1503[(1'h0):(1'h0)];
              reg1590 = {$unsigned(reg1502[(3'h5):(1'h1)])};
              reg1591 <= $unsigned(reg1577[(1'h0):(1'h0)]);
              reg1592 = {reg1573[(1'h1):(1'h0)],
                  ({wire1485[(3'h5):(2'h2)],
                      (reg1552[(1'h1):(1'h1)] ?
                          {reg1579, wire1482} : wire1483[(3'h4):(2'h3)]),
                      (7'h53)} * $unsigned({$unsigned(wire1485),
                      $unsigned((7'h40))}))};
            end
          else
            begin
              reg1589 = reg1521[(4'he):(4'ha)];
            end
        end
      else
        begin
          reg1578 <= $signed({(+$unsigned(((8'ha3) * reg1502))),
              (^~({reg1543} ? (reg1508 | (7'h4e)) : $signed(reg1580))),
              wire1482});
        end
      if ({reg1577[(4'h9):(2'h2)],
          reg1494,
          $unsigned(($unsigned((reg1553 ?
              reg1556 : reg1498)) ^ $signed(reg1507[(1'h0):(1'h0)])))})
        begin
          reg1593 <= (-$signed(reg1572));
          reg1594 = (~|(((((8'hbe) - reg1577) ?
                  $unsigned(reg1523) : (reg1517 <= (7'h4c))) <<< reg1491[(3'h6):(3'h5)]) ?
              (7'h44) : ($signed((~&(7'h51))) ?
                  (reg1560 & $signed(reg1533)) : $signed($unsigned(forvar1568)))));
        end
      else
        begin
          if (reg1570[(5'h13):(5'h11)])
            begin
              reg1594 = ($signed((8'had)) ? (^~{reg1549}) : reg1573);
              reg1595 <= $unsigned(wire1563[(4'h9):(3'h6)]);
              reg1596 <= (~|({(^((7'h53) ? (7'h4f) : reg1592))} ?
                  {$signed($unsigned(reg1523))} : (7'h54)));
              reg1597 <= {reg1505[(4'he):(3'h6)],
                  reg1588[(2'h2):(1'h0)],
                  $signed(($signed(wire1483[(5'h13):(4'hd)]) == ((reg1569 != reg1493) ?
                      (reg1578 ?
                          reg1505 : wire1563) : reg1498[(3'h7):(1'h0)])))};
              reg1598 = ({$unsigned($unsigned(reg1521))} ?
                  ((((~forvar1568) ? reg1577 : wire1483[(5'h17):(4'hf)]) ?
                          ((7'h53) ?
                              reg1536[(3'h4):(1'h1)] : {reg1515,
                                  (8'hae)}) : reg1583[(3'h4):(1'h0)]) ?
                      (7'h44) : $signed(((^(8'ha2)) ?
                          (&reg1572) : (reg1550 ?
                              reg1593 : reg1597)))) : (reg1489[(4'hf):(3'h6)] ?
                      (reg1549 ?
                          $signed({wire1485}) : ($unsigned(reg1592) ?
                              (reg1523 ?
                                  wire1485 : reg1536) : reg1578[(2'h3):(2'h3)])) : reg1569));
            end
          else
            begin
              reg1594 = $signed($unsigned(reg1494[(5'h1c):(5'h10)]));
              reg1598 = $signed(({reg1550[(3'h7):(3'h7)],
                  (^reg1519[(5'h19):(4'ha)]),
                  reg1580[(5'h13):(4'ha)]} > (reg1503[(1'h1):(1'h0)] ?
                  (reg1555[(1'h0):(1'h0)] >= wire1483) : $signed($unsigned(wire1485)))));
              reg1599 <= {reg1494[(4'ha):(1'h0)]};
              reg1600 <= (reg1511[(2'h2):(1'h0)] ?
                  $unsigned(forvar1566) : reg1519);
              reg1601 = {reg1587,
                  $signed((((~reg1586) <= reg1578[(5'h10):(3'h5)]) != (reg1594 ^ (reg1571 && wire1563))))};
              reg1602 = (~&$signed(reg1524));
            end
        end
      for (forvar1603 = (1'h0); (forvar1603 < (3'h4)); forvar1603 = (forvar1603 + (1'h1)))
        begin
          if ((&$unsigned($unsigned(($unsigned(wire1563) - $unsigned((8'hbd)))))))
            begin
              reg1604 = $unsigned(($signed({(wire1485 ? (8'had) : reg1575),
                  wire1481[(1'h1):(1'h0)],
                  reg1533}) ~^ {forvar1566}));
            end
          else
            begin
              reg1604 = $signed((wire1481 == $signed((reg1543 ?
                  (reg1567 | reg1523) : (reg1604 ? reg1584 : reg1506)))));
              reg1605 <= (reg1572[(2'h3):(1'h0)] ^ {reg1533[(1'h1):(1'h0)],
                  reg1525});
              reg1606 = ($unsigned((+(reg1581[(1'h0):(1'h0)] + {reg1601,
                      (8'had),
                      reg1538}))) ?
                  $unsigned((wire1563[(5'h18):(4'he)] ?
                      (8'ha6) : reg1503)) : (|$signed((+(reg1550 ^~ reg1514)))));
              reg1607 = reg1549;
              reg1608 <= (-(~^(~|{(!reg1581),
                  (^~reg1540),
                  (reg1523 <<< reg1578)})));
              reg1609 <= (reg1570[(5'h11):(4'ha)] > $unsigned(wire1484));
              reg1610 <= (^~reg1567[(5'h10):(1'h0)]);
            end
          reg1611 = $unsigned(reg1607[(4'hc):(4'h9)]);
          reg1612 <= reg1597;
          if ((+reg1612[(5'h10):(4'h8)]))
            begin
              reg1613 = reg1489;
              reg1614 = reg1583;
              reg1615 <= $signed(wire1482[(5'h17):(3'h5)]);
              reg1616 = ((~^reg1609[(2'h2):(1'h0)]) | reg1606[(3'h4):(1'h1)]);
            end
          else
            begin
              reg1615 <= reg1601;
              reg1616 = {{{$unsigned((reg1542 ? (7'h44) : reg1549)),
                          reg1598,
                          forvar1568},
                      reg1600,
                      $signed((reg1592[(2'h3):(1'h0)] < {reg1538}))}};
              reg1617 <= ((7'h47) ?
                  {(8'hb0),
                      ($unsigned((reg1493 ?
                          reg1610 : reg1494)) + (^~(+(8'hbf))))} : reg1498[(1'h0):(1'h0)]);
              reg1618 <= $signed($unsigned(reg1587[(5'h17):(5'h11)]));
              reg1619 = (8'hb5);
              reg1620 = (~&($unsigned(reg1570[(3'h7):(3'h7)]) >>> (reg1491 ?
                  (!wire1483[(5'h12):(4'ha)]) : reg1540)));
              reg1621 <= reg1543[(2'h2):(2'h2)];
            end
          reg1622 = $signed(((~^reg1605[(2'h2):(1'h0)]) >> reg1578));
          for (forvar1623 = (1'h0); (forvar1623 < (3'h5)); forvar1623 = (forvar1623 + (1'h1)))
            begin
              reg1624 = {(-$unsigned(((reg1605 ?
                      reg1508 : wire1562) - (|reg1581)))),
                  reg1524[(3'h4):(1'h0)]};
              reg1625 <= (^~(!(reg1617 ?
                  ((~^reg1555) ?
                      $unsigned(reg1588) : $unsigned(reg1514)) : $unsigned(reg1508[(5'h17):(3'h5)]))));
              reg1626 <= ((reg1494 ?
                  {reg1612,
                      reg1552[(1'h0):(1'h0)],
                      reg1567} : (|{$signed((8'h9d)),
                      $unsigned(reg1594)})) - (~^$signed(forvar1568)));
              reg1627 <= ((~^(8'ha3)) + (^~((reg1579 ?
                      $unsigned(reg1595) : reg1598) ?
                  (!$signed(reg1517)) : $signed(reg1624))));
              reg1628 = (reg1533[(1'h1):(1'h0)] ?
                  (8'hba) : ($signed(reg1606[(1'h0):(1'h0)]) ?
                      (reg1619 ?
                          reg1493[(5'h18):(4'ha)] : reg1616) : $unsigned($unsigned({reg1576}))));
            end
        end
      if (reg1503[(1'h0):(1'h0)])
        begin
          reg1629 = reg1542[(3'h6):(1'h0)];
          reg1630 = reg1624;
          if ({{(-reg1611[(1'h1):(1'h1)]),
                  ((|((8'ha3) ? reg1508 : reg1505)) ?
                      $signed((&reg1569)) : ($unsigned(wire1483) ?
                          {reg1589} : (|forvar1566))),
                  wire1481[(1'h0):(1'h0)]},
              $signed(forvar1623),
              reg1586})
            begin
              reg1631 <= (~^({$signed((~^reg1580)),
                      {$unsigned(reg1494),
                          (reg1569 ^ reg1512),
                          $signed(reg1592)}} ?
                  {$unsigned((~reg1597)),
                      ($signed((8'hbe)) && (~&reg1573)),
                      reg1549[(2'h2):(1'h0)]} : reg1517));
              reg1632 <= reg1585[(3'h4):(1'h0)];
              reg1633 = (8'hb5);
            end
          else
            begin
              reg1633 = reg1570;
              reg1634 = (($signed(((reg1625 ? reg1586 : wire1481) ?
                  (8'hb9) : reg1609)) & ((~^reg1573[(1'h1):(1'h1)]) ^ ($unsigned(reg1556) ?
                  wire1563 : reg1505))) | reg1627);
            end
          if ({(((~{reg1574,
                  reg1514,
                  reg1601}) << $signed(reg1597[(1'h0):(1'h0)])) >>> ((reg1519 < forvar1578[(2'h3):(2'h2)]) ?
                  $unsigned($signed(reg1505)) : reg1579)),
              $unsigned($unsigned($signed(((8'hb5) ? (8'h9d) : reg1605))))})
            begin
              reg1635 = $unsigned($signed((~^$unsigned($signed(reg1561)))));
              reg1636 = reg1524[(3'h4):(3'h4)];
              reg1637 <= forvar1566[(1'h1):(1'h0)];
              reg1638 = $unsigned(reg1626);
              reg1639 = (($signed(reg1605[(4'he):(4'h8)]) ~^ (reg1615[(2'h2):(1'h1)] ?
                      reg1560[(3'h6):(1'h1)] : {$signed(reg1514)})) ?
                  (reg1584 ?
                      reg1498[(3'h4):(1'h0)] : reg1614[(4'ha):(1'h0)]) : (+$signed(((-(7'h54)) < reg1533))));
              reg1640 = reg1621;
              reg1641 = reg1588[(1'h0):(1'h0)];
            end
          else
            begin
              reg1635 = {$unsigned(wire1563[(2'h3):(2'h2)]),
                  (+((~|$unsigned(reg1573)) * reg1579[(1'h0):(1'h0)]))};
              reg1637 <= reg1577[(5'h13):(4'h8)];
              reg1638 = (^~((^$unsigned($unsigned(reg1610))) ^ $signed((8'hbd))));
            end
          reg1642 <= $unsigned(reg1622);
          reg1643 <= ((|({(reg1491 - reg1521)} >>> ($unsigned(reg1624) ?
              $unsigned(reg1556) : (8'ha8)))) >>> ((7'h43) ~^ reg1582));
          reg1644 = ($unsigned(reg1594[(1'h1):(1'h0)]) ?
              reg1590 : (($unsigned($unsigned(reg1636)) ?
                      (|reg1618[(4'hb):(3'h5)]) : (reg1631[(1'h1):(1'h1)] ?
                          $signed(wire1563) : (reg1611 >>> (8'hb7)))) ?
                  $signed(reg1592) : $unsigned((8'hb4))));
        end
      else
        begin
          reg1631 <= reg1622[(5'h10):(5'h10)];
          if (((~^(~^(reg1552 ? $unsigned(reg1523) : {reg1543}))) ?
              reg1578[(4'ha):(1'h0)] : reg1579))
            begin
              reg1632 <= reg1593;
            end
          else
            begin
              reg1632 <= ((reg1612[(5'h15):(2'h2)] > $signed(reg1492)) ^ (7'h51));
              reg1637 <= (reg1493 ?
                  ((8'hb5) ?
                      ((~&(reg1494 - reg1574)) ?
                          {(wire1485 ? reg1616 : reg1582)} : (forvar1623 ?
                              reg1602[(4'h9):(4'h8)] : $signed(reg1614))) : ($signed((reg1585 <= wire1485)) ?
                          reg1594 : ((~&reg1619) ?
                              (reg1498 >>> reg1503) : (|(7'h46))))) : (((|reg1621[(3'h4):(2'h3)]) ?
                      (+(^reg1508)) : ($signed((8'hbb)) ?
                          reg1496[(5'h10):(4'hc)] : (reg1633 <<< reg1588))) & {reg1584}));
              reg1638 = $unsigned(((~|{(reg1538 | reg1615),
                  $unsigned((7'h4e))}) <<< reg1585[(2'h3):(1'h1)]));
            end
          reg1642 <= (!(~reg1602[(3'h6):(3'h5)]));
          for (forvar1643 = (1'h0); (forvar1643 < (3'h5)); forvar1643 = (forvar1643 + (1'h1)))
            begin
              reg1644 = wire1482[(2'h2):(1'h0)];
              reg1645 <= $unsigned($unsigned((reg1505 ?
                  ($signed(reg1540) ?
                      (reg1579 * reg1593) : reg1525) : $signed((reg1635 ?
                      (8'hab) : reg1644)))));
              reg1646 = (reg1506 == (-$unsigned(reg1489[(3'h7):(1'h0)])));
              reg1647 = ((~^($signed((reg1622 ^ reg1492)) ^ reg1635)) ^ $unsigned((&{(forvar1623 ?
                      reg1627 : reg1573),
                  $signed(reg1606),
                  $signed(reg1602)})));
              reg1648 = reg1614;
              reg1649 <= (|{$unsigned(((~^reg1540) | {reg1577,
                      reg1507,
                      reg1605})),
                  ((7'h56) + ($signed(reg1584) ?
                      (&(8'ha5)) : (reg1498 ? reg1515 : reg1612)))});
              reg1650 <= $signed((($signed($unsigned((8'h9d))) <<< $signed(reg1574[(4'hf):(4'hd)])) ~^ ($signed((reg1577 ^~ reg1610)) | (-((7'h55) ~^ forvar1568)))));
            end
          reg1651 <= (wire1483 ?
              reg1561[(2'h2):(1'h1)] : {(((reg1622 >> reg1591) >= (reg1576 ^~ reg1496)) ?
                      (8'hb2) : (wire1482[(4'hc):(3'h6)] < (reg1589 <= (7'h42)))),
                  (8'h9c)});
        end
    end
  assign wire1652 = {$unsigned((({reg1571,
                            reg1587,
                            reg1521} - $unsigned((7'h51))) & $signed((reg1631 ?
                            reg1608 : wire1484))))};
  always
    @(posedge clk) begin
      for (forvar1653 = (1'h0); (forvar1653 < (2'h2)); forvar1653 = (forvar1653 + (1'h1)))
        begin
          reg1654 = $unsigned($unsigned(reg1651));
          if ($signed({$signed(reg1524[(4'h8):(3'h5)]), reg1625}))
            begin
              reg1655 = $unsigned((~^(reg1650[(3'h6):(2'h3)] ?
                  (~|(8'h9f)) : (((8'hae) | reg1507) ?
                      {reg1538, reg1519, reg1651} : {reg1511, reg1494}))));
              reg1656 = $unsigned((8'ha4));
            end
          else
            begin
              reg1657 <= reg1543;
              reg1658 = reg1621;
              reg1659 = (~&((|(((8'haa) ?
                      wire1652 : wire1563) << reg1578[(5'h18):(1'h0)])) ?
                  ((|{(7'h45), wire1481}) < ((^~reg1538) ?
                      $signed(reg1578) : (reg1498 ?
                          reg1654 : reg1489))) : (^($unsigned(wire1483) ?
                      (reg1556 >>> reg1627) : reg1600))));
            end
          for (forvar1660 = (1'h0); (forvar1660 < (1'h0)); forvar1660 = (forvar1660 + (1'h1)))
            begin
              reg1661 = ((reg1650 > ($signed({(8'hb9),
                      reg1588}) ^ (((8'hb0) ~^ reg1596) ?
                      {reg1574, reg1621} : (reg1576 ? (8'ha7) : reg1519)))) ?
                  $unsigned((($signed((7'h41)) ? $signed(reg1625) : {reg1618}) ?
                      reg1571[(4'he):(3'h6)] : (reg1580[(5'h18):(5'h13)] ?
                          $signed(reg1599) : {reg1632,
                              reg1593,
                              reg1599}))) : (!$unsigned(reg1543[(5'h19):(3'h6)])));
              reg1662 <= reg1576[(1'h1):(1'h0)];
              reg1663 = ((~(reg1618[(4'ha):(3'h4)] ?
                  ($unsigned(wire1483) && $unsigned(reg1550)) : (7'h52))) >= $unsigned(reg1581[(1'h0):(1'h0)]));
              reg1664 <= $unsigned(($unsigned(reg1649) ?
                  $signed(reg1615[(2'h2):(2'h2)]) : (~&$unsigned({(8'hac)}))));
            end
          if ((~&reg1651[(1'h1):(1'h0)]))
            begin
              reg1665 <= {(reg1588[(2'h2):(1'h0)] ?
                      reg1503[(1'h1):(1'h0)] : reg1585[(3'h7):(1'h1)]),
                  ($unsigned((7'h53)) <= wire1485[(3'h4):(1'h1)]),
                  $signed(((reg1511[(1'h1):(1'h0)] ?
                          (reg1570 && wire1562) : (~^reg1553)) ?
                      reg1631 : $unsigned(reg1593[(1'h0):(1'h0)])))};
              reg1666 = (-(reg1491[(3'h5):(2'h2)] << (~&(&((8'hbf) ?
                  reg1588 : reg1549)))));
              reg1667 = $unsigned($unsigned(reg1498));
              reg1668 = reg1585;
              reg1669 <= $unsigned($unsigned((($unsigned((8'hbb)) > {reg1631}) ?
                  $unsigned(((8'hb3) ? reg1578 : reg1657)) : (8'ha9))));
              reg1670 = (+$signed({{(~&reg1654),
                      $unsigned(reg1645),
                      reg1595[(2'h3):(2'h2)]},
                  $signed(reg1664[(1'h0):(1'h0)])}));
              reg1671 <= ((reg1600[(3'h6):(1'h0)] | (({reg1549} << {(8'hae)}) <= {reg1662,
                      (&(8'ha1)),
                      {reg1617}})) ?
                  (reg1576[(1'h1):(1'h1)] ?
                      $signed(reg1643) : reg1595[(1'h0):(1'h0)]) : $signed((((reg1508 >= reg1491) ?
                      (reg1507 ? reg1489 : reg1511) : (reg1521 ?
                          reg1626 : reg1655)) * ($signed(reg1549) ?
                      reg1550[(4'h9):(2'h2)] : reg1505[(5'h16):(3'h4)]))));
            end
          else
            begin
              reg1666 = $signed(reg1612);
              reg1669 <= reg1580;
            end
          for (forvar1672 = (1'h0); (forvar1672 < (1'h0)); forvar1672 = (forvar1672 + (1'h1)))
            begin
              reg1673 <= $signed((wire1482[(4'h9):(4'h9)] + (|(reg1525 - (reg1665 > (8'h9e))))));
              reg1674 = reg1536[(2'h3):(2'h3)];
              reg1675 = ((-(((reg1637 >= reg1503) << $unsigned(reg1502)) ?
                  $signed($signed(wire1652)) : reg1549[(4'h8):(3'h7)])) & (~&reg1615[(2'h2):(1'h1)]));
            end
          reg1676 <= forvar1672[(1'h1):(1'h1)];
        end
      reg1677 = {$signed(reg1580),
          ($signed($signed(reg1670[(3'h4):(1'h1)])) != reg1492[(5'h16):(4'h9)])};
      if ((^((reg1580[(3'h5):(2'h2)] ?
              (-{(7'h54), reg1578}) : ((reg1512 ?
                  reg1615 : (8'ha2)) <= reg1512)) ?
          $signed(((8'hbf) * reg1593[(1'h1):(1'h0)])) : {$signed((^~wire1562))})))
        begin
          reg1678 <= reg1514;
          if ((({$signed($unsigned(reg1625))} ?
              (&$signed((!reg1612))) : (~|(~&$signed(reg1588)))) << $signed($signed($unsigned(reg1632)))))
            begin
              reg1679 = (reg1674 << $unsigned(((reg1678 ^ reg1588) ?
                  {(7'h45)} : $signed({reg1588, (8'ha6), reg1503}))));
              reg1680 = reg1612;
            end
          else
            begin
              reg1679 = $unsigned($unsigned(reg1591));
              reg1680 = ({$signed(reg1560[(4'h9):(1'h0)]),
                  (7'h41)} | (reg1627[(5'h10):(4'hd)] ?
                  $signed(($signed(reg1642) >>> {wire1484,
                      reg1561})) : reg1540));
              reg1681 = $signed((^~reg1663[(1'h0):(1'h0)]));
              reg1682 = $signed(reg1524[(4'ha):(3'h4)]);
            end
          for (forvar1683 = (1'h0); (forvar1683 < (2'h2)); forvar1683 = (forvar1683 + (1'h1)))
            begin
              reg1684 <= ($unsigned({reg1536, {wire1563}}) ?
                  {$unsigned(($unsigned(reg1667) ?
                          reg1553 : (wire1563 ? wire1485 : reg1582))),
                      (reg1662[(2'h3):(2'h3)] ~^ $signed(((8'hb0) & reg1586)))} : $unsigned(reg1585[(3'h7):(3'h6)]));
              reg1685 = $signed($signed($signed(reg1659[(5'h12):(1'h1)])));
              reg1686 <= (~($unsigned(((~reg1512) ?
                  $signed((8'hbf)) : $unsigned(reg1493))) | {(reg1668 || (reg1615 ?
                      wire1485 : reg1673)),
                  ((reg1681 - wire1483) < $unsigned(reg1605))}));
              reg1687 <= (+$signed($unsigned((~^{reg1669, reg1542}))));
              reg1688 <= $unsigned(reg1687[(4'hc):(2'h2)]);
              reg1689 = (((8'hab) + $signed(({reg1621} ?
                  {reg1684} : reg1542))) != ($signed((8'haa)) < (reg1665 & $signed($signed(reg1555)))));
              reg1690 <= reg1570;
            end
          reg1691 <= ((reg1599 == ($signed(reg1643) - {reg1582,
                  $signed((7'h45)),
                  ((8'hb1) - reg1665)})) ?
              ($unsigned({(~|reg1553), (-(7'h41)), (reg1685 != reg1519)}) ?
                  (7'h48) : reg1519) : ((|(~$signed(reg1650))) & reg1599[(4'hd):(4'h8)]));
        end
      else
        begin
          if ($signed((^(~&$signed(((7'h44) ^ reg1612))))))
            begin
              reg1678 <= (|(($unsigned($signed((7'h4f))) ?
                  $unsigned(reg1525[(5'h10):(1'h1)]) : (-{reg1690,
                      reg1543})) <= reg1626));
              reg1683 <= {$signed((~|((reg1552 ? reg1599 : (8'ha0)) ?
                      reg1512[(4'h8):(3'h5)] : (~^reg1572)))),
                  ($unsigned((((8'ha2) ?
                      forvar1683 : (7'h49)) & $unsigned(reg1556))) < ($unsigned((~reg1588)) ?
                      $signed((~^wire1562)) : $unsigned($signed(reg1595))))};
              reg1684 <= (~&(7'h49));
              reg1686 <= (-$signed((wire1484 ?
                  (((8'hbd) ? reg1687 : reg1550) ?
                      reg1514 : $unsigned(reg1506)) : $signed({reg1678,
                      reg1587,
                      (7'h49)}))));
              reg1689 = (~&$unsigned((((reg1587 ? wire1484 : reg1581) ?
                  $signed(reg1597) : reg1610[(4'hf):(3'h6)]) || $unsigned(reg1578[(4'he):(4'hd)]))));
              reg1692 = {reg1582[(2'h2):(1'h1)],
                  $unsigned((((8'hb9) >= (forvar1683 << reg1609)) <= ({reg1637,
                      reg1496} || $signed(reg1682))))};
            end
          else
            begin
              reg1679 = reg1655;
              reg1680 = $unsigned($unsigned(reg1645));
              reg1683 <= reg1585[(3'h6):(1'h0)];
              reg1684 <= $unsigned($signed($signed((&(7'h4d)))));
            end
          for (forvar1693 = (1'h0); (forvar1693 < (2'h2)); forvar1693 = (forvar1693 + (1'h1)))
            begin
              reg1694 <= $unsigned((!(((reg1682 >= reg1662) >>> wire1481[(2'h3):(2'h3)]) ?
                  (reg1668 < reg1680[(2'h3):(2'h3)]) : ($signed(reg1519) + reg1508))));
            end
          reg1695 = ({$signed(((reg1608 ? reg1576 : wire1652) ?
                      $signed(reg1553) : $unsigned(reg1521))),
                  reg1684} ?
              $unsigned($signed(reg1651)) : $signed($signed(wire1652[(1'h0):(1'h0)])));
          reg1696 = (($signed(reg1655) ? $signed($signed(reg1587)) : reg1521) ?
              $signed(reg1605[(3'h5):(1'h0)]) : reg1574);
          reg1697 = wire1483;
          reg1698 <= reg1676[(2'h2):(1'h0)];
          for (forvar1699 = (1'h0); (forvar1699 < (1'h1)); forvar1699 = (forvar1699 + (1'h1)))
            begin
              reg1700 <= reg1654[(3'h4):(3'h4)];
              reg1701 = {({$unsigned((&reg1700))} << reg1561[(1'h0):(1'h0)]),
                  $signed(forvar1683),
                  (-(reg1494 ?
                      (reg1605[(3'h4):(2'h3)] << (&reg1668)) : $signed($signed((8'ha9)))))};
              reg1702 <= reg1494;
              reg1703 <= (reg1688 ?
                  $signed($unsigned((reg1550[(4'h9):(3'h4)] ^ ((8'ha1) ?
                      reg1588 : reg1550)))) : reg1676[(2'h2):(1'h1)]);
              reg1704 = $signed((!$unsigned($unsigned(reg1656[(2'h2):(1'h1)]))));
            end
        end
      reg1705 <= reg1536;
      reg1706 <= (8'hb1);
      if (((reg1657 ? reg1702 : $signed({$unsigned(reg1618)})) ?
          {$signed(reg1560),
              (-reg1503)} : (~&((!(forvar1683 ^~ reg1591)) - $signed($unsigned(reg1610))))))
        begin
          reg1707 <= reg1605[(1'h0):(1'h0)];
        end
      else
        begin
          reg1708 = ($unsigned($signed(reg1651)) * ($unsigned(reg1503) || $unsigned(reg1696[(1'h1):(1'h0)])));
          reg1709 <= $unsigned(($signed($unsigned({reg1524})) + reg1645[(2'h3):(1'h1)]));
          if ($signed($signed($signed($unsigned((reg1679 < reg1685))))))
            begin
              reg1710 = (reg1655 >>> ((reg1533[(3'h5):(2'h3)] == $unsigned(forvar1699[(3'h7):(1'h0)])) ?
                  {((reg1492 ? reg1572 : reg1659) ?
                          $signed(reg1621) : (reg1618 <<< reg1709))} : {$signed(reg1625),
                      (&$signed(reg1608))}));
              reg1711 <= $signed((7'h49));
              reg1712 <= (^~$signed(reg1687[(4'he):(4'hd)]));
              reg1713 <= reg1553[(4'hc):(1'h1)];
            end
          else
            begin
              reg1711 <= $signed((-wire1485));
              reg1714 = (~$unsigned($signed($unsigned((reg1489 ?
                  reg1632 : reg1496)))));
            end
          reg1715 <= ((((7'h48) <= reg1714) > (^$signed(reg1680[(4'h9):(2'h2)]))) ?
              {(reg1657 ?
                      reg1578 : ($signed((8'hbd)) ?
                          (reg1517 ?
                              reg1680 : reg1591) : $signed(forvar1672)))} : (7'h47));
        end
    end
  always
    @(posedge clk) begin
      reg1716 <= (~&{reg1574});
    end
  always
    @(posedge clk) begin
      reg1717 = ($signed({reg1618, reg1703}) ?
          reg1496[(5'h11):(5'h11)] : (&((&reg1715[(3'h4):(3'h4)]) ?
              {(!reg1688), (-(8'ha7))} : reg1586)));
    end
  always
    @(posedge clk) begin
      reg1718 <= {$signed(wire1485)};
      if (wire1484[(1'h1):(1'h1)])
        begin
          reg1719 <= reg1596;
          if (((+reg1517[(1'h1):(1'h0)]) && $unsigned($signed($signed((+reg1678))))))
            begin
              reg1720 = (~&(~$signed(((reg1709 * (7'h44)) >= $signed(reg1540)))));
            end
          else
            begin
              reg1720 = wire1484[(1'h1):(1'h1)];
              reg1721 <= ($unsigned(((^~$unsigned(reg1519)) >>> (~^reg1694[(4'he):(1'h1)]))) && reg1709[(5'h11):(3'h4)]);
              reg1722 = $unsigned($signed(reg1618));
              reg1723 <= ((8'hb5) ?
                  (~$unsigned(reg1690[(4'hc):(4'hc)])) : {reg1694});
              reg1724 = ($signed($unsigned(reg1718[(2'h3):(1'h1)])) != reg1596[(2'h2):(1'h1)]);
              reg1725 = ($signed({((!reg1662) ?
                      $signed(reg1538) : ((8'ha1) ? (8'ha9) : (7'h44))),
                  {(reg1626 | (8'ha9)), reg1503},
                  {(reg1570 ? reg1621 : (8'ha0)),
                      reg1496[(5'h10):(4'hf)],
                      (&(8'hbf))}}) << $signed((~|(~&{reg1657, (7'h4f)}))));
            end
          for (forvar1726 = (1'h0); (forvar1726 < (2'h2)); forvar1726 = (forvar1726 + (1'h1)))
            begin
              reg1727 <= $unsigned((reg1657 + $unsigned($signed({(8'hbe),
                  reg1536,
                  wire1485}))));
              reg1728 = {(&wire1484),
                  (reg1706[(4'hc):(3'h7)] < $signed({reg1518[(4'hd):(1'h0)],
                      $unsigned(wire1482)})),
                  (reg1686 ?
                      $signed(($signed(reg1712) ?
                          (reg1524 - (7'h53)) : reg1676)) : (|$unsigned((~reg1493))))};
              reg1729 = $signed(reg1720);
            end
          for (forvar1730 = (1'h0); (forvar1730 < (2'h2)); forvar1730 = (forvar1730 + (1'h1)))
            begin
              reg1731 <= reg1725;
            end
          reg1732 = ((^~$signed($unsigned(reg1519))) ?
              reg1514 : {$signed((-{(7'h43)})),
                  (8'hbb),
                  (reg1555[(4'hc):(3'h7)] ?
                      ($signed(reg1642) ? (|reg1706) : reg1621) : (~^{reg1605,
                          reg1507}))});
        end
      else
        begin
          if (wire1482)
            begin
              reg1720 = reg1700;
            end
          else
            begin
              reg1719 <= (reg1498 ?
                  {$signed(reg1632[(3'h7):(2'h2)]),
                      $unsigned(($unsigned((8'ha2)) == (reg1578 * reg1580))),
                      $signed((reg1669 ^~ $unsigned((7'h46))))} : (8'h9e));
              reg1720 = reg1694;
            end
          for (forvar1721 = (1'h0); (forvar1721 < (1'h1)); forvar1721 = (forvar1721 + (1'h1)))
            begin
              reg1723 <= wire1562[(3'h5):(2'h2)];
              reg1726 <= $unsigned(({((^reg1561) + (^~reg1645)),
                      ((^reg1683) ? {reg1582} : (^~(8'hbf))),
                      $unsigned($unsigned(reg1665))} ?
                  (((~^(7'h4f)) >> (reg1571 ? reg1533 : reg1657)) ?
                      (^~(reg1662 * (7'h51))) : $signed((reg1625 ?
                          reg1694 : reg1627))) : reg1556[(4'hd):(4'hb)]));
              reg1727 <= ({(|$unsigned((reg1508 <<< wire1481))),
                      ((|$signed((8'hb6))) ?
                          (reg1561[(2'h2):(1'h0)] + (reg1511 ?
                              reg1627 : reg1637)) : ($signed((7'h44)) <<< (8'hb5)))} ?
                  {(|{(~^reg1698), reg1514[(5'h19):(5'h12)]}),
                      reg1489} : $unsigned((8'h9c)));
              reg1728 = $signed(({((!reg1664) ?
                          (reg1542 <= reg1631) : (-reg1706))} ?
                  reg1580 : forvar1726));
            end
        end
      for (forvar1733 = (1'h0); (forvar1733 < (2'h3)); forvar1733 = (forvar1733 + (1'h1)))
        begin
          reg1734 = reg1688;
          reg1735 = $unsigned(((reg1580[(5'h12):(4'h9)] ?
              {((8'hbd) == reg1560),
                  (reg1576 ?
                      reg1600 : (8'ha2))} : $unsigned({(8'haa)})) - reg1515));
          reg1736 <= $signed($unsigned(reg1503));
          if (($unsigned(($signed((reg1706 ? reg1736 : reg1588)) >>> reg1724)) ?
              wire1563 : $signed(forvar1730)))
            begin
              reg1737 <= reg1676;
              reg1738 = reg1657;
              reg1739 <= reg1723[(3'h5):(1'h1)];
              reg1740 <= $signed({reg1514, reg1553});
              reg1741 = {reg1678,
                  $signed((7'h42)),
                  ((|reg1595) - $signed($signed((reg1632 ?
                      reg1715 : reg1518))))};
              reg1742 <= ((reg1684 ?
                  $signed(reg1525[(4'h8):(3'h7)]) : (reg1702 ?
                      reg1673 : reg1739)) ~^ ($unsigned(wire1483) * reg1723));
            end
          else
            begin
              reg1738 = reg1694[(4'h8):(2'h3)];
            end
          if (reg1580)
            begin
              reg1743 = (~|($signed((|(reg1632 || reg1540))) >= (~$unsigned(reg1728[(1'h0):(1'h0)]))));
              reg1744 = (~reg1600);
              reg1745 = $unsigned(((($unsigned(reg1540) ?
                  ((8'hb5) <<< reg1684) : {reg1729, reg1494}) ^ ({reg1608,
                      reg1505,
                      (8'hb1)} ?
                  ((8'hb9) ?
                      reg1552 : reg1650) : $unsigned(reg1587))) < (+($unsigned(reg1643) >> reg1507[(1'h1):(1'h0)]))));
              reg1746 <= reg1578[(5'h14):(5'h14)];
              reg1747 = reg1745;
              reg1748 <= ($signed((+($unsigned((8'haa)) >= wire1652))) ?
                  ($unsigned(($unsigned(reg1709) >>> (reg1649 ?
                          reg1683 : reg1715))) ?
                      {$signed($signed(reg1691)),
                          reg1627,
                          ($signed(reg1687) ^~ $signed(reg1555))} : $signed(($unsigned(reg1561) ?
                          ((8'hb9) || reg1494) : (forvar1721 - reg1524)))) : reg1512);
              reg1749 = $signed(reg1555[(1'h1):(1'h0)]);
            end
          else
            begin
              reg1743 = (~|((+reg1560[(3'h7):(1'h0)]) ?
                  $unsigned($unsigned(reg1720[(3'h7):(1'h1)])) : ((reg1587[(5'h1a):(3'h6)] - reg1728[(5'h12):(3'h4)]) ?
                      ((8'hb4) ^~ {reg1637}) : {reg1599,
                          {(8'ha3), reg1716, reg1556}})));
              reg1744 = $signed((reg1671[(2'h3):(2'h3)] >= $unsigned($signed((reg1673 ?
                  (8'h9c) : reg1540)))));
              reg1746 <= {((^~$unsigned((reg1626 ?
                      (8'hab) : reg1538))) <<< reg1731),
                  ($unsigned(reg1574) ^~ (+reg1627[(4'hf):(4'h9)]))};
              reg1747 = (($signed((^$signed(reg1713))) ^~ forvar1730) ?
                  (~|$signed(((reg1489 ? (8'h9f) : wire1652) < (reg1726 ?
                      reg1600 : reg1734)))) : reg1649[(4'ha):(3'h4)]);
              reg1748 <= (8'ha3);
              reg1750 <= reg1684;
              reg1751 <= (((+(-$unsigned(reg1731))) && $signed($signed($unsigned(reg1581)))) && $signed(($unsigned(reg1718) ?
                  $signed($unsigned(wire1483)) : (reg1515[(3'h5):(3'h4)] ?
                      (reg1519 < reg1553) : ((8'hb2) << reg1506)))));
            end
          reg1752 <= reg1665[(4'he):(2'h2)];
        end
      reg1753 <= reg1518[(5'h10):(3'h6)];
      reg1754 = reg1538;
      reg1755 = {reg1627[(4'h9):(2'h2)]};
    end
  always
    @(posedge clk) begin
      if ((reg1508[(5'h1a):(3'h7)] ?
          $signed(reg1645[(1'h0):(1'h0)]) : ((reg1742[(2'h2):(2'h2)] ?
                  reg1662[(4'hd):(3'h5)] : (&reg1627)) ?
              (reg1705[(5'h13):(4'hb)] <<< $signed(reg1585[(1'h0):(1'h0)])) : reg1645[(2'h3):(1'h1)])))
        begin
          reg1756 <= reg1650[(2'h3):(2'h3)];
          reg1757 = reg1505[(3'h5):(3'h5)];
          reg1758 <= $signed(reg1691);
          if (((-(({reg1665, reg1715} ? (8'ha6) : $signed(reg1752)) ?
              reg1750 : $unsigned(reg1631[(4'h8):(3'h6)]))) > reg1736[(1'h0):(1'h0)]))
            begin
              reg1759 = reg1727;
              reg1760 <= (~|(reg1571[(1'h0):(1'h0)] << (|reg1711[(1'h1):(1'h0)])));
            end
          else
            begin
              reg1759 = reg1574;
              reg1761 = $signed(reg1517[(3'h7):(1'h0)]);
              reg1762 <= (reg1617 >>> reg1605);
            end
        end
      else
        begin
          if (((&(|$unsigned(reg1515[(5'h15):(5'h11)]))) ~^ reg1642[(5'h11):(3'h5)]))
            begin
              reg1757 = {($signed((reg1609[(4'h8):(4'h8)] >= reg1707)) << reg1752[(4'he):(4'h9)]),
                  (~^reg1494[(4'hd):(4'hb)])};
              reg1758 <= reg1556;
              reg1759 = $signed(((+{reg1705, reg1540}) ?
                  (~(reg1555 ?
                      reg1553 : reg1612[(5'h16):(4'ha)])) : $unsigned({$unsigned((8'hb6)),
                      $unsigned(reg1758),
                      (&reg1719)})));
            end
          else
            begin
              reg1756 <= ($unsigned(((!{reg1493,
                      reg1631,
                      wire1484}) * $unsigned({reg1612, (7'h49), reg1507}))) ?
                  reg1760[(4'hb):(1'h1)] : $unsigned($unsigned(((|wire1563) ?
                      {reg1626, reg1574} : reg1739))));
              reg1757 = reg1596[(4'h9):(3'h6)];
              reg1758 <= $signed(((7'h51) * ($signed(reg1627) ?
                  {(reg1600 <<< reg1690)} : (~reg1723))));
              reg1759 = {{({(~&reg1552), {(8'hae)}} & reg1698[(2'h3):(2'h2)])},
                  $unsigned({$unsigned((reg1512 ~^ (7'h51))),
                      reg1517[(4'h9):(2'h3)]})};
            end
          for (forvar1760 = (1'h0); (forvar1760 < (1'h0)); forvar1760 = (forvar1760 + (1'h1)))
            begin
              reg1761 = $unsigned((((~&$unsigned(reg1494)) > ((reg1665 * (8'hb7)) ?
                      $unsigned(reg1489) : (-reg1673))) ?
                  (^reg1662[(5'h15):(4'hd)]) : ((reg1739[(3'h5):(2'h3)] == reg1700) ?
                      ($signed(reg1711) >= reg1514[(4'hd):(3'h4)]) : reg1560[(1'h0):(1'h0)])));
              reg1763 = (reg1761[(3'h5):(3'h4)] ?
                  (reg1608 ?
                      $signed((reg1515 + ((7'h44) ?
                          wire1484 : (7'h44)))) : {(reg1713 ?
                              $unsigned(reg1698) : (~reg1637)),
                          $unsigned(reg1700[(1'h0):(1'h0)]),
                          $signed(reg1711[(3'h6):(3'h4)])}) : (($signed(reg1610[(5'h19):(5'h15)]) | ((~|reg1703) ^ $unsigned(reg1740))) && {{{reg1719,
                              reg1571,
                              reg1587}}}));
              reg1764 = ($unsigned(reg1506) <= $unsigned($unsigned(((-reg1610) ?
                  (reg1664 ? reg1700 : reg1605) : reg1742))));
              reg1765 = $signed(reg1494);
              reg1766 = (7'h41);
              reg1767 <= ((~^{reg1492,
                      ($signed(reg1542) * $unsigned((8'hb5))),
                      ({reg1610, (7'h48)} || $signed(reg1686))}) ?
                  (^(~|(reg1669 ? (reg1621 << reg1581) : reg1746))) : reg1726);
              reg1768 <= reg1540;
            end
        end
    end
  assign wire1769 = $unsigned({(~&{{reg1517, reg1574, (8'hb5)}, (~|reg1713)}),
                        $unsigned($unsigned((reg1571 ? (8'ha8) : reg1502)))});
  assign wire1770 = (reg1716 * (~^$signed(((wire1652 >= reg1750) ~^ $signed(reg1518)))));
  always
    @(posedge clk) begin
      if (reg1753[(4'hb):(2'h3)])
        begin
          reg1771 = (reg1758[(2'h2):(1'h0)] >= ($unsigned(reg1721[(3'h6):(3'h6)]) * $unsigned((^~reg1610))));
          reg1772 <= $signed($unsigned((~&$signed(reg1706))));
          reg1773 <= ((~|reg1715[(1'h1):(1'h1)]) ?
              $signed({(reg1505 ?
                      (reg1507 >>> reg1574) : (reg1493 ?
                          reg1687 : reg1615))}) : (reg1525[(3'h7):(2'h3)] >> (~(|(wire1563 ?
                  reg1585 : reg1737)))));
          if ($signed((&$signed($signed(reg1686)))))
            begin
              reg1774 = {reg1709[(5'h10):(3'h6)],
                  ($unsigned(reg1711) != reg1552[(1'h0):(1'h0)])};
              reg1775 = reg1560;
              reg1776 = {reg1570[(4'hc):(4'h9)],
                  ((((reg1665 != reg1748) ?
                              (reg1774 && reg1615) : $signed(reg1707)) ?
                          (^~((8'h9c) >>> reg1549)) : (&(wire1563 ?
                              wire1769 : reg1676))) ?
                      (reg1543[(1'h1):(1'h0)] * (+(reg1645 << reg1600))) : reg1687)};
              reg1777 <= ((8'ha4) ?
                  (7'h4d) : ((({reg1758, reg1493, (7'h41)} ?
                          wire1563[(5'h16):(4'h9)] : reg1683) ^~ {$unsigned(reg1737)}) ?
                      (reg1772[(3'h7):(3'h6)] >> reg1758[(1'h0):(1'h0)]) : ((^~reg1760) >>> $signed({reg1518,
                          reg1493}))));
              reg1778 <= ($signed((|$unsigned(reg1632))) ?
                  reg1711 : $unsigned((7'h58)));
              reg1779 = (+reg1651);
              reg1780 <= ({reg1760[(4'h9):(3'h5)],
                      (reg1521 - ($unsigned((8'ha5)) & $unsigned(reg1580)))} ?
                  {reg1515,
                      $unsigned($unsigned((7'h50)))} : $signed($unsigned((((8'h9d) * (8'h9c)) << (reg1669 > reg1649)))));
            end
          else
            begin
              reg1777 <= (($signed(reg1684[(1'h1):(1'h1)]) ?
                      $unsigned((+reg1698[(3'h6):(3'h6)])) : (reg1767[(3'h6):(3'h6)] == (((7'h4a) << reg1651) ?
                          $unsigned((8'ha5)) : $signed(reg1760)))) ?
                  $unsigned({((^reg1706) ?
                          (reg1684 || reg1742) : $unsigned(wire1770))}) : (~^(^reg1723[(1'h0):(1'h0)])));
              reg1778 <= ((~|{$signed(reg1780),
                  (reg1774 ? (reg1746 ? reg1615 : (8'haa)) : $signed(reg1571)),
                  $unsigned($unsigned(reg1610))}) ~^ ((~{$signed(reg1570),
                      reg1712,
                      $signed(reg1519)}) ?
                  $signed({$unsigned((7'h48))}) : $unsigned($unsigned((reg1772 ^~ reg1599)))));
            end
        end
      else
        begin
          for (forvar1771 = (1'h0); (forvar1771 < (3'h6)); forvar1771 = (forvar1771 + (1'h1)))
            begin
              reg1774 = $signed(((^~{(8'hbb)}) ?
                  (^~$signed(((8'hbf) ^ reg1626))) : ((~|$unsigned(reg1706)) ?
                      $signed((+reg1571)) : ((wire1769 ? reg1772 : reg1664) ?
                          (7'h49) : (-reg1760)))));
            end
          for (forvar1775 = (1'h0); (forvar1775 < (3'h4)); forvar1775 = (forvar1775 + (1'h1)))
            begin
              reg1777 <= $signed(((+reg1691[(1'h1):(1'h0)]) ?
                  ($signed($unsigned(reg1727)) <<< (~|reg1582[(1'h0):(1'h0)])) : reg1493[(5'h15):(5'h14)]));
              reg1778 <= reg1621[(3'h5):(2'h2)];
            end
          for (forvar1779 = (1'h0); (forvar1779 < (1'h1)); forvar1779 = (forvar1779 + (1'h1)))
            begin
              reg1780 <= $unsigned(reg1514);
              reg1781 <= (7'h42);
              reg1782 <= $signed((!{reg1676}));
            end
          reg1783 = {reg1683[(1'h1):(1'h1)],
              (reg1712 ~^ $unsigned(({reg1627} | (reg1645 + reg1649))))};
          if ($signed((reg1596[(2'h3):(1'h1)] != ($signed($unsigned(reg1712)) & ($signed((7'h42)) <= reg1727)))))
            begin
              reg1784 = $signed({{reg1555, (&reg1582[(1'h1):(1'h0)])},
                  forvar1771[(4'h9):(3'h6)],
                  reg1600[(3'h7):(2'h2)]});
              reg1785 = reg1496[(2'h3):(1'h1)];
              reg1786 = (!(!reg1587));
              reg1787 <= wire1484;
              reg1788 = reg1560[(2'h3):(1'h1)];
            end
          else
            begin
              reg1784 = ($signed((~$signed(reg1762))) - $unsigned((reg1618[(3'h4):(1'h1)] ^~ reg1767[(5'h10):(4'he)])));
              reg1785 = $unsigned((forvar1771 ?
                  (!{(|reg1489), reg1753[(4'hc):(3'h4)]}) : (7'h45)));
            end
        end
      reg1789 <= (wire1482 << reg1649);
      for (forvar1790 = (1'h0); (forvar1790 < (3'h6)); forvar1790 = (forvar1790 + (1'h1)))
        begin
          for (forvar1791 = (1'h0); (forvar1791 < (2'h2)); forvar1791 = (forvar1791 + (1'h1)))
            begin
              reg1792 <= $signed($signed((^~(~|(-(8'hb4))))));
              reg1793 <= {($signed(reg1586) | ({$unsigned(reg1574)} ^~ reg1713[(3'h4):(2'h2)])),
                  ({$unsigned((|reg1649)),
                          {(+(7'h44)),
                              $unsigned(reg1792),
                              forvar1771[(2'h2):(1'h0)]},
                          $signed(reg1498[(4'h9):(4'h9)])} ?
                      reg1691 : (+(8'h9e))),
                  (~^$unsigned(({reg1599, reg1649} ?
                      (reg1518 ?
                          reg1621 : reg1727) : reg1739[(4'hd):(4'hd)])))};
              reg1794 <= reg1756[(3'h5):(2'h3)];
              reg1795 = reg1684;
            end
          reg1796 <= {($unsigned((~&(8'h9d))) ?
                  ({(8'hb9),
                      (~|reg1795),
                      (reg1678 ?
                          reg1709 : reg1739)} ^ ($unsigned(reg1788) <= (~^reg1752))) : (reg1588[(1'h0):(1'h0)] ?
                      reg1712 : (reg1665 * reg1570[(4'ha):(4'h9)])))};
          if ((reg1678 <= reg1739))
            begin
              reg1797 = $signed(reg1576);
              reg1798 = $unsigned(($signed($signed(reg1795[(5'h10):(3'h5)])) ?
                  reg1525[(2'h3):(2'h2)] : reg1507));
              reg1799 = $signed(reg1676[(3'h4):(2'h3)]);
            end
          else
            begin
              reg1797 = reg1760;
              reg1800 <= $unsigned(({reg1543[(4'h9):(1'h0)],
                      reg1748,
                      ({reg1707, wire1483, (8'ha1)} & (reg1727 == reg1505))} ?
                  reg1751[(3'h5):(2'h2)] : ((reg1787 < reg1721) - reg1784[(5'h11):(4'hc)])));
              reg1801 = reg1712;
              reg1802 = reg1794;
            end
          reg1803 <= (reg1570[(4'hf):(4'hc)] ~^ $signed({reg1576[(1'h0):(1'h0)],
              (~{reg1570, reg1756, reg1585}),
              ((^~forvar1775) < (reg1492 ^~ reg1555))}));
          for (forvar1804 = (1'h0); (forvar1804 < (3'h5)); forvar1804 = (forvar1804 + (1'h1)))
            begin
              reg1805 <= $unsigned(((reg1707 >= reg1776) + (($unsigned(reg1731) ?
                      (~&reg1794) : reg1502[(5'h15):(5'h11)]) ?
                  {reg1502} : $unsigned((reg1794 <<< reg1760)))));
              reg1806 = reg1718;
              reg1807 <= $unsigned((reg1540[(2'h2):(2'h2)] ?
                  (^~$unsigned(reg1632)) : $unsigned((~(reg1801 ?
                      (8'h9f) : reg1508)))));
            end
          reg1808 = (((8'ha8) << ((reg1784[(5'h19):(5'h11)] ?
                  reg1771 : (reg1691 & reg1515)) ?
              reg1703 : ((reg1511 - reg1610) >> $unsigned(reg1802)))) ^ ($unsigned((&(+reg1684))) || (($signed(reg1519) ?
                  (reg1669 ? reg1556 : reg1793) : {reg1773, reg1605}) ?
              (+$unsigned(reg1605)) : ($signed(reg1496) * (~|reg1560)))));
          reg1809 = {(({$unsigned(reg1721)} > $unsigned((reg1801 && reg1719))) ?
                  $unsigned({reg1651[(2'h2):(1'h0)],
                      (reg1688 ^~ reg1673)}) : reg1777[(1'h0):(1'h0)]),
              $signed($unsigned(reg1774[(4'hc):(4'h9)])),
              reg1700};
        end
      reg1810 = $unsigned($signed((8'h9e)));
      reg1811 = reg1756;
    end
  assign wire1812 = (&(({(reg1514 >= reg1746),
                        {wire1482,
                            (7'h4e),
                            reg1536}} == ((^reg1758) <= ((8'h9d) ?
                        reg1626 : reg1684))) & ({reg1645,
                        wire1769} + reg1751)));
  assign wire1813 = $unsigned((($unsigned((reg1552 ~^ wire1485)) == (&(reg1742 ?
                        reg1637 : wire1485))) >> $unsigned($signed(reg1762))));
  always
    @(posedge clk) begin
      reg1814 <= (~|(&{(~|(reg1752 ? reg1787 : (8'hb4))),
          $signed((&reg1519))}));
      if ({(reg1780[(1'h1):(1'h1)] == ((reg1756 ?
              (reg1570 ?
                  (7'h53) : reg1617) : ((8'hba) ^~ reg1512)) + (|reg1767[(5'h1f):(4'hf)]))),
          reg1605[(5'h10):(4'he)]})
        begin
          if (reg1716[(2'h3):(2'h3)])
            begin
              reg1815 = wire1483[(4'hf):(4'he)];
              reg1816 = $unsigned((&($unsigned(reg1585) ?
                  (reg1721 ? wire1769 : reg1496) : $unsigned(reg1690))));
            end
          else
            begin
              reg1815 = reg1803;
            end
          if (reg1493[(5'h13):(3'h6)])
            begin
              reg1817 = reg1773;
              reg1818 = reg1574;
              reg1819 = $signed(reg1591);
            end
          else
            begin
              reg1820 <= ($unsigned(reg1515) + $signed(reg1711[(1'h0):(1'h0)]));
              reg1821 = $unsigned((^(8'hb8)));
            end
          reg1822 <= reg1706;
          reg1823 = reg1700;
          reg1824 = reg1503;
          for (forvar1825 = (1'h0); (forvar1825 < (1'h1)); forvar1825 = (forvar1825 + (1'h1)))
            begin
              reg1826 <= (~^{reg1605,
                  (reg1627 <= $signed((+reg1617))),
                  reg1505[(5'h10):(2'h2)]});
              reg1827 <= reg1768[(1'h1):(1'h0)];
              reg1828 = {(&$unsigned($signed($signed(reg1556)))),
                  (reg1792[(1'h0):(1'h0)] ?
                      (($unsigned(reg1794) ?
                              reg1506[(3'h4):(3'h4)] : (reg1796 - (7'h49))) ?
                          {reg1615[(2'h2):(2'h2)],
                              (reg1492 ?
                                  reg1517 : reg1678)} : {reg1703}) : (~|$unsigned((~|reg1489))))};
              reg1829 <= (+(7'h51));
              reg1830 = $unsigned(($signed(reg1508[(5'h19):(3'h4)]) > (((reg1703 + reg1750) * (~^reg1503)) ?
                  reg1694[(5'h1b):(5'h14)] : {$unsigned(reg1740),
                      reg1768,
                      (reg1507 ^ reg1829)})));
              reg1831 <= (($signed({reg1822, $unsigned((7'h54))}) ?
                  $unsigned($signed((~^reg1489))) : wire1482) ^~ reg1507[(1'h1):(1'h1)]);
              reg1832 <= $signed((&reg1823));
            end
        end
      else
        begin
          reg1815 = (reg1781 == (reg1561 > ($signed(reg1662) ?
              (^~(reg1828 ?
                  (8'ha7) : reg1781)) : $signed($unsigned((8'hbf))))));
          for (forvar1816 = (1'h0); (forvar1816 < (3'h5)); forvar1816 = (forvar1816 + (1'h1)))
            begin
              reg1820 <= reg1823[(2'h2):(1'h0)];
              reg1821 = $unsigned($signed({($unsigned(reg1574) && reg1550[(2'h2):(1'h1)]),
                  (~|{(7'h48), reg1508}),
                  (~|(reg1817 ? reg1686 : reg1610))}));
            end
        end
      reg1833 <= {(~^$signed(reg1726[(4'h8):(3'h4)])),
          $unsigned((((8'hb2) ?
              ((8'ha6) ? reg1506 : reg1816) : (reg1752 ?
                  reg1597 : (8'hb2))) || wire1484))};
    end
  assign wire1834 = $signed(reg1615);
  assign wire1835 = ($signed((8'h9d)) ?
                        ((!reg1517[(1'h1):(1'h1)]) == {((^~reg1700) ^~ {(8'haa),
                                reg1746,
                                (8'ha8)}),
                            (!((8'h9f) ?
                                reg1591 : reg1800))}) : reg1773[(3'h7):(1'h0)]);
  assign wire1836 = {$unsigned(($signed({reg1767,
                            reg1756,
                            (8'ha8)}) >= ((~^reg1665) >>> (reg1533 ?
                            reg1800 : reg1515)))),
                        reg1600[(5'h1c):(5'h18)]};
  always
    @(posedge clk) begin
      for (forvar1837 = (1'h0); (forvar1837 < (3'h4)); forvar1837 = (forvar1837 + (1'h1)))
        begin
          reg1838 = $unsigned({$signed(wire1562),
              reg1570[(5'h14):(4'h8)],
              (($signed(reg1773) >= wire1836[(2'h3):(2'h3)]) > ((reg1782 ^~ (8'hae)) != (!(8'ha0))))});
          reg1839 <= (~(reg1593 >>> reg1760));
          if ((~&(~^$unsigned((-$signed(reg1571))))))
            begin
              reg1840 = $signed($unsigned($unsigned(((reg1803 != (8'hb6)) ?
                  reg1632 : (reg1642 ~^ reg1593)))));
              reg1841 <= reg1642;
              reg1842 = $unsigned($unsigned(((7'h45) * ((8'hb0) ?
                  $unsigned(reg1665) : (reg1536 != (8'hab))))));
              reg1843 = $unsigned(reg1596);
            end
          else
            begin
              reg1841 <= $signed($signed($signed(reg1796)));
              reg1844 <= ($unsigned(((forvar1837 ?
                          (~reg1555) : $signed((7'h45))) ?
                      (~$unsigned(reg1657)) : (+$unsigned((7'h4c))))) ?
                  reg1723[(4'he):(4'ha)] : ({(((7'h40) ? (8'ha9) : reg1827) ?
                              reg1814 : $signed(reg1773)),
                          $unsigned($unsigned(reg1570))} ?
                      reg1580 : ((~&(~^reg1580)) ?
                          ($signed(wire1563) ?
                              (^~reg1687) : (reg1502 <<< reg1586)) : reg1691[(4'hf):(4'hc)])));
              reg1845 <= reg1507;
              reg1846 <= $unsigned(($unsigned($unsigned((~&reg1742))) + $unsigned(($signed((7'h51)) && (reg1793 | reg1578)))));
              reg1847 <= (reg1796 ^ (~^((|reg1608[(4'h9):(2'h3)]) && $signed((reg1842 ?
                  reg1683 : reg1615)))));
              reg1848 = $signed(reg1542[(3'h4):(1'h1)]);
            end
          for (forvar1849 = (1'h0); (forvar1849 < (3'h5)); forvar1849 = (forvar1849 + (1'h1)))
            begin
              reg1850 <= {reg1712[(5'h12):(4'he)]};
            end
          for (forvar1851 = (1'h0); (forvar1851 < (3'h4)); forvar1851 = (forvar1851 + (1'h1)))
            begin
              reg1852 = $unsigned($signed($unsigned((^(reg1669 ?
                  (8'hba) : reg1618)))));
              reg1853 = reg1599[(5'h1a):(4'hb)];
              reg1854 = {$signed($signed($unsigned(reg1740[(3'h7):(3'h7)]))),
                  reg1847[(3'h4):(1'h0)],
                  ($signed(reg1570[(4'hc):(2'h3)]) ?
                      (+((reg1787 <= reg1687) || $unsigned(reg1726))) : reg1702)};
              reg1855 <= (!(8'hb0));
              reg1856 = ({(~|({reg1782} <<< reg1768))} || $unsigned(wire1770[(1'h0):(1'h0)]));
              reg1857 <= (wire1835[(4'hc):(2'h2)] ?
                  reg1669[(5'h13):(3'h5)] : (!($signed((reg1707 >= reg1621)) >= $unsigned($signed(reg1572)))));
            end
        end
      reg1858 <= $signed(reg1687[(4'ha):(3'h5)]);
      if (($unsigned({reg1618[(3'h5):(3'h5)],
          (wire1834[(2'h3):(2'h2)] < {reg1593,
              wire1836,
              reg1665})}) ^ $unsigned(reg1524[(3'h6):(3'h4)])))
        begin
          if ({reg1731})
            begin
              reg1859 = {$unsigned($signed((^(reg1686 ? reg1632 : reg1787)))),
                  wire1482,
                  ((((^reg1581) ?
                          (~^wire1652) : {reg1838,
                              reg1586}) ^~ (reg1496[(3'h5):(1'h1)] << (reg1706 ?
                          (7'h41) : reg1805))) ?
                      $signed(reg1839[(4'hb):(3'h5)]) : (($signed(reg1605) ?
                          (~&(8'ha4)) : (reg1673 >>> reg1773)) | {(reg1691 >>> (8'hb1)),
                          reg1715}))};
              reg1860 = $signed($unsigned(((8'hb4) || (reg1542 & (^reg1719)))));
              reg1861 = (^(|($signed((reg1571 ? (7'h4f) : (8'hbe))) ?
                  wire1813 : (reg1581 ? reg1846 : (^reg1854)))));
            end
          else
            begin
              reg1862 <= (|($signed($unsigned($unsigned(reg1736))) > $signed((~(reg1777 || reg1664)))));
              reg1863 <= ((~|(~&($signed(reg1829) ?
                  $unsigned(reg1742) : $unsigned(reg1498)))) || ({$unsigned((reg1773 ?
                          reg1571 : reg1756))} ?
                  reg1750 : $signed($unsigned((8'hbc)))));
              reg1864 <= (~^(&(!(~|((8'hae) ? reg1780 : reg1700)))));
            end
          reg1865 <= $unsigned($unsigned($unsigned(wire1483[(4'hc):(3'h7)])));
          reg1866 <= (($signed(reg1595) ?
              reg1822 : (&(^~$unsigned(reg1517)))) | reg1671);
          reg1867 <= $signed(reg1864[(5'h16):(3'h4)]);
          reg1868 = reg1574[(1'h1):(1'h0)];
          for (forvar1869 = (1'h0); (forvar1869 < (2'h3)); forvar1869 = (forvar1869 + (1'h1)))
            begin
              reg1870 <= (^~$unsigned((|($signed(reg1643) ?
                  $unsigned(reg1847) : reg1657))));
              reg1871 = (&reg1847[(3'h4):(1'h1)]);
            end
          reg1872 <= (8'hb8);
        end
      else
        begin
          for (forvar1859 = (1'h0); (forvar1859 < (1'h1)); forvar1859 = (forvar1859 + (1'h1)))
            begin
              reg1862 <= (~|reg1618);
              reg1863 <= reg1686[(4'ha):(3'h4)];
              reg1864 <= (~|reg1582);
              reg1868 = (~&reg1542[(3'h5):(2'h2)]);
            end
          for (forvar1869 = (1'h0); (forvar1869 < (3'h6)); forvar1869 = (forvar1869 + (1'h1)))
            begin
              reg1871 = reg1617;
              reg1873 = reg1625;
              reg1874 = $unsigned((7'h49));
              reg1875 <= $unsigned(($signed(reg1574[(4'he):(2'h2)]) > ($signed((~^wire1484)) || $signed((~&wire1484)))));
              reg1876 = reg1731;
              reg1877 = reg1651[(2'h2):(1'h0)];
              reg1878 = reg1588;
            end
        end
      for (forvar1879 = (1'h0); (forvar1879 < (1'h1)); forvar1879 = (forvar1879 + (1'h1)))
        begin
          for (forvar1880 = (1'h0); (forvar1880 < (1'h1)); forvar1880 = (forvar1880 + (1'h1)))
            begin
              reg1881 = $signed(((reg1587 == reg1721[(3'h5):(2'h3)]) < ($signed((~^wire1835)) ?
                  reg1586 : {$unsigned((8'haa)), $signed(reg1760)})));
              reg1882 = (reg1690[(4'hc):(4'ha)] ^~ (~^((reg1593 || (reg1665 > reg1829)) ?
                  {(reg1872 + reg1760), reg1829} : (8'hb6))));
              reg1883 = $unsigned(reg1698[(3'h7):(1'h0)]);
              reg1884 = $unsigned(reg1582);
              reg1885 <= (8'hb1);
            end
          reg1886 = $unsigned((~^reg1698));
          reg1887 = $signed(reg1833[(4'h8):(3'h5)]);
          reg1888 = $unsigned((reg1703[(2'h2):(1'h0)] != ((reg1571[(4'h8):(1'h1)] != reg1716) ?
              ({reg1600, reg1498} & (!(8'hb9))) : reg1882)));
        end
      for (forvar1889 = (1'h0); (forvar1889 < (2'h3)); forvar1889 = (forvar1889 + (1'h1)))
        begin
          for (forvar1890 = (1'h0); (forvar1890 < (3'h6)); forvar1890 = (forvar1890 + (1'h1)))
            begin
              reg1891 <= $unsigned((reg1773[(5'h15):(3'h6)] < $signed($signed((reg1688 || wire1834)))));
            end
          for (forvar1892 = (1'h0); (forvar1892 < (2'h3)); forvar1892 = (forvar1892 + (1'h1)))
            begin
              reg1893 <= $signed($signed((($signed(wire1485) && $signed(reg1847)) & $unsigned(reg1632))));
              reg1894 <= (reg1852 ?
                  (reg1886 & {$signed((reg1617 ? reg1690 : reg1588)),
                      reg1829,
                      {(wire1812 ?
                              (7'h47) : (7'h57))}}) : (reg1748[(1'h0):(1'h0)] || $signed(reg1847[(1'h1):(1'h0)])));
            end
          reg1895 = reg1871;
          reg1896 <= $signed((((+$unsigned((8'hbb))) >> ($unsigned((7'h52)) + $signed(wire1482))) ?
              ({(forvar1859 != (7'h4a)),
                  (reg1895 || reg1794),
                  (!reg1599)} >>> $signed($signed((7'h43)))) : (8'hbf)));
          if ((~^reg1894[(1'h0):(1'h0)]))
            begin
              reg1897 <= reg1760[(4'hc):(4'hb)];
            end
          else
            begin
              reg1897 <= (({$signed({reg1690})} ?
                  reg1866 : {((~^reg1855) ?
                          $unsigned(reg1523) : {reg1827,
                              reg1768})}) | reg1550[(3'h4):(2'h2)]);
              reg1898 = (($signed((~^(reg1715 ^ reg1688))) ?
                      $signed(($signed(reg1517) ?
                          (reg1864 > reg1807) : {(8'ha8)})) : $signed(reg1846[(1'h1):(1'h1)])) ?
                  reg1678 : reg1588);
              reg1899 <= reg1841;
              reg1900 <= (reg1895[(1'h1):(1'h0)] >= reg1605);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1901 = (1'h0); (forvar1901 < (1'h1)); forvar1901 = (forvar1901 + (1'h1)))
        begin
          if ($signed(reg1826[(5'h10):(4'he)]))
            begin
              reg1902 <= $signed($signed($unsigned((-(reg1618 ?
                  reg1669 : reg1758)))));
              reg1903 <= ((((~&reg1751) >>> (reg1591 && reg1844[(4'h9):(1'h0)])) ^~ {reg1793,
                  (!(reg1767 ? (8'hbd) : (7'h45))),
                  (~|reg1827)}) ^~ ((+reg1683[(1'h0):(1'h0)]) == reg1844));
              reg1904 = $signed((reg1719 ^~ reg1793[(4'h8):(1'h0)]));
              reg1905 <= $signed((-(|(reg1858 ?
                  {reg1560, reg1617} : (reg1505 && reg1723)))));
              reg1906 = $signed((+$unsigned(({(7'h50), reg1517, (7'h54)} ?
                  (reg1593 ? (8'hb1) : reg1820) : {(7'h46)}))));
            end
          else
            begin
              reg1902 <= ((~^$unsigned(reg1751[(1'h0):(1'h0)])) ?
                  $unsigned(wire1770[(1'h1):(1'h1)]) : $signed(wire1770[(1'h1):(1'h1)]));
              reg1904 = reg1521;
              reg1906 = (8'hb0);
              reg1907 <= $signed((reg1642[(4'hf):(4'he)] > reg1803));
              reg1908 = {(!reg1673)};
              reg1909 = $unsigned(($unsigned(({reg1907} ?
                      $unsigned(reg1496) : (reg1833 ? reg1719 : reg1831))) ?
                  ({$unsigned(reg1706),
                      reg1493[(4'h9):(3'h7)],
                      {reg1597, (7'h57)}} >>> wire1482) : (reg1700 ?
                      ((wire1485 + reg1536) == (-reg1748)) : $signed(reg1600[(4'hb):(4'hb)]))));
              reg1910 = reg1512;
            end
          if ((-(reg1800 ?
              (((reg1796 ? reg1758 : reg1688) ?
                  reg1904 : (7'h57)) ^ reg1829) : reg1694)))
            begin
              reg1911 <= (((!(+(7'h56))) <= $unsigned(reg1555[(1'h1):(1'h1)])) >>> $signed((!reg1863)));
              reg1912 <= reg1585[(4'h8):(2'h3)];
              reg1913 <= reg1572[(1'h0):(1'h0)];
              reg1914 = ((((^$unsigned(reg1649)) != (reg1582 ?
                          $unsigned(reg1605) : $signed((7'h54)))) ?
                      $signed(wire1652[(1'h0):(1'h0)]) : (^~reg1712[(3'h5):(1'h0)])) ?
                  $signed($signed({reg1731[(2'h2):(2'h2)]})) : reg1894);
            end
          else
            begin
              reg1911 <= ((wire1563 * reg1865) ?
                  reg1683 : {$signed(reg1691), reg1900, $unsigned((7'h43))});
              reg1914 = reg1706;
              reg1915 <= reg1850[(2'h2):(1'h0)];
              reg1916 <= reg1748;
              reg1917 <= reg1610[(4'hc):(4'h9)];
              reg1918 = $signed($signed($unsigned((&(reg1600 <= (7'h52))))));
              reg1919 <= {wire1563[(3'h5):(1'h1)],
                  ($signed($unsigned(reg1600[(4'hf):(4'he)])) * (+($unsigned(reg1600) ?
                      reg1746[(1'h0):(1'h0)] : (~^reg1493))))};
            end
          reg1920 <= reg1665;
          for (forvar1921 = (1'h0); (forvar1921 < (3'h6)); forvar1921 = (forvar1921 + (1'h1)))
            begin
              reg1922 <= ($signed(((^~{reg1669}) < (reg1690 ~^ (reg1713 ?
                  (8'hb8) : reg1726)))) != {reg1822[(3'h4):(1'h1)],
                  ({reg1588[(2'h3):(1'h1)]} >> reg1768)});
              reg1923 = {reg1902};
              reg1924 <= reg1905;
              reg1925 <= (+(reg1758 < $signed((+reg1870[(2'h3):(2'h3)]))));
            end
          reg1926 = (reg1691[(5'h12):(4'hc)] >> reg1631);
          for (forvar1927 = (1'h0); (forvar1927 < (3'h4)); forvar1927 = (forvar1927 + (1'h1)))
            begin
              reg1928 = (~|(~|($unsigned(reg1572) && (7'h40))));
              reg1929 <= (^~($unsigned((reg1706[(5'h10):(2'h2)] - (!(8'hae)))) ?
                  (^reg1891) : $unsigned((^~wire1482))));
              reg1930 = $signed($unsigned((^((^~reg1642) > reg1691[(5'h10):(1'h1)]))));
              reg1931 <= reg1845;
              reg1932 <= ($signed($signed($signed((|reg1796)))) > (+$signed({reg1718,
                  reg1571})));
              reg1933 <= (^~(^~$unsigned(($signed(reg1800) ?
                  $signed((7'h46)) : $unsigned(wire1652)))));
              reg1934 <= $unsigned(({$signed((reg1542 || reg1787)),
                  (~&(reg1694 * reg1705))} >= (8'ha2)));
            end
          reg1935 <= ((~&reg1841) ^ wire1652);
        end
    end
  assign wire1936 = {reg1826[(2'h2):(1'h0)]};
  always
    @(posedge clk) begin
      for (forvar1937 = (1'h0); (forvar1937 < (2'h3)); forvar1937 = (forvar1937 + (1'h1)))
        begin
          reg1938 <= (8'hb9);
          if ($signed($signed(reg1718[(1'h0):(1'h0)])))
            begin
              reg1939 = {$signed((($signed(reg1596) ?
                      $unsigned(reg1492) : reg1618[(1'h0):(1'h0)]) <<< reg1875)),
                  reg1515,
                  ($signed((-(reg1793 ? (7'h57) : reg1858))) + reg1553)};
            end
          else
            begin
              reg1939 = (|{$unsigned($unsigned(reg1694[(2'h2):(1'h1)]))});
            end
          for (forvar1940 = (1'h0); (forvar1940 < (3'h6)); forvar1940 = (forvar1940 + (1'h1)))
            begin
              reg1941 = ((|$unsigned((7'h43))) ?
                  (|$unsigned(reg1758)) : reg1561);
              reg1942 = ($unsigned(($signed($unsigned(reg1715)) | reg1705[(1'h0):(1'h0)])) | ((({reg1600,
                              reg1870} ?
                          (reg1512 ? reg1503 : (8'ha9)) : (reg1715 ?
                              reg1700 : reg1864)) ?
                      ({(8'hb1)} ?
                          reg1746[(1'h0):(1'h0)] : reg1939) : (~|reg1915[(1'h1):(1'h1)])) ?
                  wire1936 : reg1665[(4'ha):(1'h1)]));
              reg1943 = $signed((8'ha1));
              reg1944 = reg1807[(4'h9):(1'h1)];
              reg1945 = wire1770[(1'h1):(1'h0)];
              reg1946 = (reg1609[(3'h5):(1'h0)] >>> reg1872[(4'hd):(1'h0)]);
            end
        end
      if ((7'h54))
        begin
          reg1947 = ({reg1715[(3'h5):(3'h4)],
                  $signed((|(reg1615 ? reg1885 : reg1787))),
                  (~&{$unsigned(reg1931), (reg1525 & reg1650)})} ?
              (~|((^reg1807[(3'h5):(3'h4)]) ?
                  (reg1932 ~^ $signed(reg1632)) : $signed((reg1872 != reg1642)))) : {reg1870,
                  reg1711});
          for (forvar1948 = (1'h0); (forvar1948 < (3'h4)); forvar1948 = (forvar1948 + (1'h1)))
            begin
              reg1949 <= ((reg1933[(4'h8):(2'h2)] ?
                      reg1839[(4'hc):(3'h5)] : (7'h40)) ?
                  ((|(!$unsigned(reg1676))) ?
                      reg1715[(2'h3):(1'h1)] : ((forvar1937[(1'h1):(1'h0)] | reg1855[(4'hb):(3'h6)]) ?
                          $unsigned((~|reg1582)) : reg1578)) : (~|reg1588));
              reg1950 = $signed((-($unsigned({reg1894, reg1643, reg1900}) ?
                  reg1913[(5'h13):(4'h8)] : (^~$unsigned(reg1803)))));
              reg1951 = (reg1657 ?
                  (~&reg1777[(1'h1):(1'h0)]) : (-($signed({wire1834,
                      reg1933,
                      reg1515}) <<< (reg1919 + $unsigned(reg1950)))));
              reg1952 <= (+(~^$signed((reg1651[(1'h0):(1'h0)] ?
                  (reg1502 ? reg1905 : reg1705) : (~reg1543)))));
              reg1953 <= reg1657[(1'h1):(1'h1)];
              reg1954 <= reg1715;
              reg1955 = (($unsigned(reg1899) * (((!reg1896) ?
                      $unsigned((8'hba)) : (wire1482 ?
                          reg1846 : reg1493)) > {$unsigned(reg1944),
                      reg1903})) ?
                  reg1931 : ($unsigned(reg1867[(3'h4):(2'h3)]) != $unsigned(({reg1756} <<< reg1707[(2'h2):(1'h0)]))));
            end
          reg1956 = {$signed(reg1538)};
          reg1957 = $signed((-{reg1855[(2'h3):(1'h1)],
              ((|reg1866) ?
                  reg1855[(2'h3):(2'h3)] : {reg1912, reg1939, reg1726})}));
        end
      else
        begin
          reg1948 <= reg1518;
          reg1949 <= ($unsigned(($signed((reg1931 ? wire1562 : reg1899)) ?
                  (reg1831[(3'h4):(1'h1)] ?
                      $signed(reg1561) : $unsigned((8'hbe))) : reg1731)) ?
              $unsigned(reg1643) : ($unsigned((wire1484 != $unsigned(reg1673))) ?
                  (&reg1687[(1'h1):(1'h0)]) : (reg1705[(3'h7):(2'h3)] ?
                      ($unsigned(reg1864) ?
                          reg1922 : $unsigned(reg1576)) : {reg1850})));
          reg1952 <= reg1524[(2'h3):(1'h1)];
          reg1953 <= ($signed(({reg1945[(2'h2):(1'h1)],
                  $signed(reg1896),
                  reg1678[(4'h8):(3'h5)]} == reg1939)) ?
              $unsigned(reg1847[(2'h2):(1'h1)]) : (!{reg1637[(3'h4):(3'h4)]}));
        end
      for (forvar1958 = (1'h0); (forvar1958 < (2'h2)); forvar1958 = (forvar1958 + (1'h1)))
        begin
          for (forvar1959 = (1'h0); (forvar1959 < (1'h0)); forvar1959 = (forvar1959 + (1'h1)))
            begin
              reg1960 = reg1736[(4'h8):(3'h4)];
            end
          for (forvar1961 = (1'h0); (forvar1961 < (1'h1)); forvar1961 = (forvar1961 + (1'h1)))
            begin
              reg1962 <= (&(~|(+{((8'hbc) ? wire1769 : reg1581)})));
              reg1963 <= (^$signed($unsigned($signed(((8'hb9) == wire1813)))));
              reg1964 <= ((^~$signed(reg1955[(5'h12):(4'hb)])) && ((((reg1832 ?
                              reg1489 : reg1827) ?
                          (reg1542 ? reg1960 : reg1683) : reg1827) ?
                      (((7'h50) ? reg1924 : reg1512) ?
                          reg1913[(3'h6):(2'h3)] : $unsigned((8'hac))) : $signed((+(8'ha5)))) ?
                  $unsigned($unsigned((8'had))) : ($signed($signed(reg1610)) <= $unsigned(reg1524))));
              reg1965 <= reg1793[(4'h8):(3'h5)];
            end
          reg1966 = reg1845[(2'h3):(2'h2)];
          reg1967 <= reg1922[(4'hb):(4'h8)];
        end
    end
  always
    @(posedge clk) begin
      if ((($unsigned(((^(7'h4a)) ? (~&reg1706) : (wire1812 << reg1581))) ?
              (reg1731[(1'h1):(1'h0)] >> $signed(reg1608)) : (reg1841[(5'h13):(4'h9)] + $unsigned($signed((8'ha5))))) ?
          $unsigned(($signed((reg1772 ? reg1686 : reg1867)) ?
              $signed(reg1872) : ((reg1556 - reg1542) ?
                  $unsigned((8'hb8)) : {(7'h50),
                      reg1748}))) : ({$signed(((8'h9d) ? (7'h45) : wire1483))} ?
              ((reg1920 <= (8'hb4)) ?
                  reg1608 : ((-reg1586) == (~&reg1781))) : ((!$signed((7'h46))) ?
                  ((reg1752 ? reg1571 : reg1649) ?
                      $unsigned(reg1782) : (~^reg1595)) : $unsigned({reg1772})))))
        begin
          for (forvar1968 = (1'h0); (forvar1968 < (3'h4)); forvar1968 = (forvar1968 + (1'h1)))
            begin
              reg1969 = {(($unsigned($signed(reg1953)) && $unsigned((reg1862 && (8'ha6)))) == ($signed((-reg1760)) ?
                      $signed(reg1727) : (reg1931 ^ ((8'hab) ?
                          reg1954 : reg1952)))),
                  ($signed(reg1907) <<< reg1964[(5'h18):(4'hf)]),
                  (!reg1593)};
              reg1970 = (reg1552 ?
                  reg1525[(5'h13):(4'h9)] : reg1864[(4'hd):(4'h9)]);
              reg1971 <= (reg1615[(1'h0):(1'h0)] ?
                  reg1718 : $unsigned(((^reg1736[(1'h0):(1'h0)]) ?
                      {reg1803,
                          $unsigned(reg1870),
                          (^reg1903)} : {reg1793[(2'h2):(2'h2)], {(8'h9c)}})));
            end
          reg1972 <= ((-reg1605[(2'h3):(2'h2)]) ?
              ({$signed($signed((8'ha7))),
                  reg1807[(4'hc):(4'h8)]} ~^ (^~{(reg1550 ?
                      (8'hac) : reg1687)})) : $unsigned((((reg1512 + (8'hac)) & (reg1572 || reg1814)) ?
                  reg1962 : reg1777)));
          reg1973 = $unsigned(({$unsigned((-reg1916)),
                  (^~reg1702[(4'hb):(3'h6)])} ?
              $unsigned((|{reg1726,
                  (7'h4d),
                  reg1543})) : reg1736[(3'h6):(2'h3)]));
          reg1974 <= (reg1615[(2'h3):(1'h0)] ?
              reg1586[(5'h15):(5'h13)] : reg1867);
        end
      else
        begin
          reg1968 = ($signed(reg1847) <<< $signed((&{wire1812, reg1727})));
          if (((wire1812 >> (8'ha6)) >>> reg1716))
            begin
              reg1969 = (reg1932 ?
                  ((+$unsigned(reg1740[(3'h6):(1'h0)])) > (^~$signed(reg1578))) : $unsigned($signed(reg1571)));
              reg1971 <= reg1753[(4'hd):(3'h4)];
              reg1973 = {(!$signed((+reg1525))), (^reg1521), reg1591};
              reg1975 = reg1841[(1'h0):(1'h0)];
              reg1976 <= $signed($signed(reg1931[(3'h6):(3'h6)]));
              reg1977 <= {$signed($unsigned(($signed(reg1750) ?
                      (reg1651 >> reg1625) : reg1698[(3'h6):(3'h6)]))),
                  $unsigned({$unsigned((reg1517 > reg1913)),
                      {$signed(reg1907), (~&(8'hb7)), reg1864}})};
              reg1978 <= (-((~&reg1793[(3'h7):(3'h5)]) ?
                  {((reg1949 ? reg1493 : reg1637) ?
                          reg1844[(3'h5):(2'h2)] : {reg1727})} : (!$unsigned(reg1748[(5'h10):(3'h4)]))));
            end
          else
            begin
              reg1971 <= $unsigned(($signed($unsigned(reg1712)) ?
                  ((8'hb1) ?
                      ($signed(reg1971) << reg1805) : (8'haf)) : reg1511));
              reg1973 = reg1781;
            end
          reg1979 <= (&((reg1649 ?
              reg1493 : (reg1807[(4'ha):(4'h9)] ?
                  $signed(reg1489) : (reg1618 ?
                      reg1919 : (7'h53)))) == $unsigned($signed((reg1506 >> reg1683)))));
          reg1980 <= {wire1834};
        end
      reg1981 = ((~|{reg1891, $signed(reg1581)}) ?
          {$signed(reg1967),
              (reg1561[(1'h1):(1'h1)] <= $signed(wire1483[(4'he):(3'h7)]))} : $signed(reg1833));
      reg1982 = $signed(reg1676);
      reg1983 <= reg1662[(5'h19):(4'hb)];
      reg1984 <= {({reg1814[(3'h4):(1'h0)],
                  $unsigned($signed(reg1983)),
                  ($signed(reg1494) <= $signed(reg1686))} ?
              ($signed(reg1931[(4'h9):(1'h0)]) ?
                  (~^(-wire1769)) : reg1875[(1'h1):(1'h1)]) : reg1847[(3'h4):(3'h4)]),
          (~|reg1703[(4'he):(4'hb)]),
          (~|$unsigned(($signed(reg1550) <<< ((7'h48) ^~ reg1673))))};
    end
  assign wire1985 = $signed(reg1974);
  assign wire1986 = reg1596[(2'h3):(2'h3)];
  assign wire1987 = reg1627[(4'ha):(1'h1)];
  assign wire1988 = (reg1814[(1'h0):(1'h0)] * $signed(reg1595));
  assign wire1989 = reg1502;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1387
#(parameter param1477 = {(~|(8'hae))})
(y, clk, wire1391, wire1390, wire1389, wire1388);
  output wire [(32'h633):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire1391;
  input wire [(5'h1a):(1'h0)] wire1390;
  input wire [(5'h1c):(1'h0)] wire1389;
  input wire [(4'hb):(1'h0)] wire1388;
  wire signed [(5'h1f):(1'h0)] wire1476;
  wire [(3'h6):(1'h0)] wire1473;
  wire signed [(3'h5):(1'h0)] wire1472;
  wire [(3'h4):(1'h0)] wire1471;
  wire [(3'h7):(1'h0)] wire1470;
  wire signed [(5'h1f):(1'h0)] wire1394;
  reg signed [(4'h8):(1'h0)] reg1475 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1467 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1466 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1461 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1458 = (1'h0);
  reg [(5'h12):(1'h0)] reg1456 = (1'h0);
  reg [(5'h14):(1'h0)] reg1455 = (1'h0);
  reg [(4'he):(1'h0)] reg1454 = (1'h0);
  reg [(3'h5):(1'h0)] reg1452 = (1'h0);
  reg [(5'h16):(1'h0)] reg1451 = (1'h0);
  reg [(4'he):(1'h0)] reg1450 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1449 = (1'h0);
  reg [(4'hd):(1'h0)] reg1448 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1447 = (1'h0);
  reg [(5'h12):(1'h0)] reg1445 = (1'h0);
  reg [(5'h11):(1'h0)] reg1443 = (1'h0);
  reg [(5'h15):(1'h0)] reg1439 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1438 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1437 = (1'h0);
  reg [(4'hf):(1'h0)] reg1436 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1433 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1432 = (1'h0);
  reg [(4'h9):(1'h0)] reg1430 = (1'h0);
  reg [(4'hc):(1'h0)] reg1424 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1422 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1417 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1416 = (1'h0);
  reg [(2'h2):(1'h0)] reg1415 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1410 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1404 = (1'h0);
  reg [(5'h10):(1'h0)] reg1401 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1400 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1399 = (1'h0);
  reg [(4'hf):(1'h0)] reg1397 = (1'h0);
  reg [(5'h18):(1'h0)] reg1396 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1393 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1392 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1474 = (1'h0);
  reg [(5'h15):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1468 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1465 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1464 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1463 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1462 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1454 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1460 = (1'h0);
  reg [(5'h15):(1'h0)] reg1459 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1457 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1453 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1446 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1444 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar1442 = (1'h0);
  reg [(2'h3):(1'h0)] reg1441 = (1'h0);
  reg [(4'h9):(1'h0)] reg1440 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1435 = (1'h0);
  reg [(5'h11):(1'h0)] reg1434 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1431 = (1'h0);
  reg [(3'h7):(1'h0)] reg1429 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1428 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1427 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1426 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1425 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1423 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar1421 = (1'h0);
  reg [(2'h2):(1'h0)] reg1420 = (1'h0);
  reg [(5'h12):(1'h0)] reg1419 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1418 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1414 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1413 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1412 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1411 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1409 = (1'h0);
  reg [(4'hc):(1'h0)] reg1408 = (1'h0);
  reg [(5'h11):(1'h0)] reg1407 = (1'h0);
  reg [(5'h14):(1'h0)] reg1406 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1405 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1403 = (1'h0);
  reg [(4'hf):(1'h0)] reg1402 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1398 = (1'h0);
  reg [(4'hb):(1'h0)] reg1395 = (1'h0);
  assign y = {wire1476,
                 wire1473,
                 wire1472,
                 wire1471,
                 wire1470,
                 wire1394,
                 reg1475,
                 reg1467,
                 reg1466,
                 reg1461,
                 reg1458,
                 reg1456,
                 reg1455,
                 reg1454,
                 reg1452,
                 reg1451,
                 reg1450,
                 reg1449,
                 reg1448,
                 reg1447,
                 reg1445,
                 reg1443,
                 reg1439,
                 reg1438,
                 reg1437,
                 reg1436,
                 reg1433,
                 reg1432,
                 reg1430,
                 reg1424,
                 reg1422,
                 reg1417,
                 reg1416,
                 reg1415,
                 reg1410,
                 reg1404,
                 reg1401,
                 reg1400,
                 reg1399,
                 reg1397,
                 reg1396,
                 reg1393,
                 reg1392,
                 reg1474,
                 reg1469,
                 reg1468,
                 reg1465,
                 reg1464,
                 reg1463,
                 reg1462,
                 forvar1454,
                 reg1460,
                 reg1459,
                 reg1457,
                 reg1453,
                 forvar1446,
                 reg1444,
                 forvar1442,
                 reg1441,
                 reg1440,
                 reg1435,
                 reg1434,
                 reg1431,
                 reg1429,
                 forvar1428,
                 reg1427,
                 forvar1426,
                 reg1425,
                 reg1423,
                 forvar1421,
                 reg1420,
                 reg1419,
                 reg1418,
                 reg1414,
                 reg1413,
                 reg1412,
                 reg1411,
                 forvar1409,
                 reg1408,
                 reg1407,
                 reg1406,
                 reg1405,
                 reg1403,
                 reg1402,
                 reg1398,
                 reg1395,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1392 <= ($unsigned($unsigned((~&(wire1391 & wire1390)))) ?
          ($signed($signed($signed(wire1389))) ?
              (^~wire1390[(5'h11):(2'h2)]) : ($signed((^wire1390)) ?
                  {$signed(wire1390),
                      $signed(wire1390),
                      wire1391} : ($signed(wire1389) ?
                      (wire1388 <<< wire1388) : wire1390))) : wire1391);
      reg1393 <= ({{{(reg1392 ^~ wire1389), (^~wire1388), $signed(reg1392)}},
              wire1388[(4'h9):(1'h1)]} ?
          (~^wire1388) : $unsigned(wire1389));
    end
  assign wire1394 = ($unsigned((8'ha7)) != reg1393);
  always
    @(posedge clk) begin
      reg1395 = {wire1389[(5'h10):(1'h0)]};
      if (wire1390[(5'h14):(4'hb)])
        begin
          if ({(wire1394 ^~ $signed(wire1388[(1'h1):(1'h1)])),
              $signed($unsigned(wire1389[(5'h12):(4'hb)]))})
            begin
              reg1396 <= (~^(wire1388[(4'h9):(4'h9)] != (-(8'ha8))));
              reg1397 <= ((reg1393 ?
                  ({wire1389[(5'h19):(3'h7)]} ^~ (~^wire1394)) : (wire1394[(5'h1d):(5'h14)] | (~wire1388))) || $unsigned((wire1394[(4'ha):(4'ha)] > reg1392)));
              reg1398 = (^wire1391);
            end
          else
            begin
              reg1396 <= $signed($signed((|reg1396[(5'h10):(4'h8)])));
              reg1398 = $unsigned({$unsigned($unsigned((wire1390 ?
                      reg1395 : reg1398)))});
              reg1399 <= (reg1398[(4'hd):(2'h2)] >>> ({($unsigned(wire1390) ^~ {(7'h53),
                      reg1392,
                      wire1391}),
                  $unsigned($signed(wire1389))} || ((reg1397 >> $signed(wire1391)) == reg1395)));
            end
          if (((!reg1397[(3'h4):(1'h1)]) ?
              reg1398[(5'h17):(5'h17)] : (|{(^~(reg1398 ?
                      (8'ha4) : (8'hac)))})))
            begin
              reg1400 <= (!wire1389[(4'hf):(3'h5)]);
              reg1401 <= ({reg1393[(3'h5):(1'h0)],
                      $signed($signed((reg1397 ^~ wire1391)))} ?
                  (wire1391 > (reg1400[(5'h11):(2'h2)] ?
                      reg1398[(5'h11):(3'h7)] : wire1394[(3'h4):(3'h4)])) : $signed(wire1391));
              reg1402 = (((|(reg1393 ? (&reg1396) : $signed(wire1388))) ?
                      $unsigned((~|reg1401[(3'h7):(1'h0)])) : reg1395[(4'hb):(4'h9)]) ?
                  reg1400[(3'h6):(1'h0)] : $unsigned(({$signed((8'h9f))} ^ wire1390[(5'h14):(3'h6)])));
              reg1403 = $signed((-$signed({$signed(reg1402),
                  {(8'ha1), wire1388, reg1398},
                  $signed(reg1402)})));
              reg1404 <= ((~&({$unsigned((8'ha8))} ?
                      reg1399[(2'h2):(1'h1)] : (+wire1391))) ?
                  (reg1397[(1'h1):(1'h0)] <= $signed({$unsigned(reg1392),
                      $unsigned(reg1399),
                      $signed((7'h49))})) : reg1401);
            end
          else
            begin
              reg1402 = $unsigned((({((8'ha1) || (8'hbf))} ?
                      $unsigned(reg1400[(3'h6):(1'h0)]) : $unsigned(reg1397)) ?
                  (reg1400 ?
                      (!(+reg1397)) : $unsigned($signed(reg1398))) : reg1395));
              reg1403 = {reg1397[(4'h8):(3'h7)],
                  $signed(reg1402[(1'h1):(1'h1)]),
                  $unsigned(reg1404)};
              reg1404 <= ((reg1395[(4'hb):(1'h1)] ?
                  (+reg1400) : $unsigned($unsigned($unsigned(wire1389)))) ~^ $signed($unsigned(($unsigned(reg1397) - {reg1400,
                  wire1390,
                  reg1399}))));
              reg1405 = ($signed((7'h47)) ?
                  (reg1403[(4'hc):(4'h9)] ?
                      $unsigned((~wire1391)) : $signed((^~{wire1389}))) : (|reg1395));
              reg1406 = ($signed(($signed($unsigned(reg1396)) == ((reg1404 ?
                  reg1396 : wire1390) < $unsigned(reg1402)))) < (-$unsigned($unsigned((^~reg1404)))));
              reg1407 = {$signed($signed(((wire1389 >>> reg1397) == $signed(wire1390)))),
                  $unsigned($signed(((reg1403 | reg1392) ^ (reg1397 & (8'hb4)))))};
              reg1408 = $signed(($signed((8'ha5)) ?
                  $unsigned(((|reg1393) || $signed(reg1401))) : ((wire1394[(3'h6):(1'h1)] << (wire1390 ?
                          wire1391 : reg1396)) ?
                      $unsigned(reg1392[(2'h2):(1'h1)]) : reg1393[(3'h4):(1'h1)])));
            end
          for (forvar1409 = (1'h0); (forvar1409 < (3'h4)); forvar1409 = (forvar1409 + (1'h1)))
            begin
              reg1410 <= reg1397;
              reg1411 = (~&(8'ha1));
            end
          reg1412 = (+$signed(wire1388));
          reg1413 = (~&(reg1410[(2'h2):(2'h2)] ^~ (&$unsigned((reg1396 ?
              reg1405 : reg1393)))));
        end
      else
        begin
          reg1398 = reg1410;
        end
      if ($unsigned(((8'hbb) ?
          (~|((|reg1412) ?
              (reg1410 - reg1400) : (reg1393 ? reg1397 : reg1406))) : reg1408)))
        begin
          reg1414 = (reg1393[(1'h0):(1'h0)] ?
              $unsigned((((8'hae) ?
                  reg1393[(2'h3):(1'h0)] : (forvar1409 + reg1393)) < $signed(((7'h54) ?
                  wire1389 : reg1400)))) : ($signed(reg1407) ?
                  reg1392[(3'h5):(3'h4)] : (reg1395 ?
                      reg1407[(4'hf):(4'h8)] : (reg1413 ?
                          reg1397 : (reg1396 || reg1400)))));
        end
      else
        begin
          reg1414 = reg1397;
          if (((&($signed(reg1406) ^ {$signed(reg1413)})) ~^ (7'h52)))
            begin
              reg1415 <= reg1405[(4'h9):(3'h7)];
            end
          else
            begin
              reg1415 <= reg1398[(5'h11):(3'h5)];
              reg1416 <= (-$signed(reg1413[(5'h1a):(5'h17)]));
              reg1417 <= reg1402;
              reg1418 = {(~&(+(reg1393 & (~|reg1416))))};
            end
          reg1419 = $unsigned($unsigned({(^$signed(wire1389)),
              wire1389[(2'h3):(2'h2)]}));
          reg1420 = reg1399;
          for (forvar1421 = (1'h0); (forvar1421 < (3'h6)); forvar1421 = (forvar1421 + (1'h1)))
            begin
              reg1422 <= $unsigned((~|$signed(reg1405[(4'hd):(3'h6)])));
              reg1423 = reg1412[(2'h3):(2'h3)];
              reg1424 <= forvar1421;
              reg1425 = wire1391;
            end
        end
      for (forvar1426 = (1'h0); (forvar1426 < (3'h6)); forvar1426 = (forvar1426 + (1'h1)))
        begin
          reg1427 = (~&(~^$signed(wire1394)));
          for (forvar1428 = (1'h0); (forvar1428 < (3'h4)); forvar1428 = (forvar1428 + (1'h1)))
            begin
              reg1429 = wire1391;
              reg1430 <= reg1417;
              reg1431 = (~|(^((reg1404[(1'h0):(1'h0)] ?
                      (&reg1422) : $unsigned(reg1413)) ?
                  (+(reg1416 ^~ (8'hac))) : ((reg1411 >> reg1403) == (|reg1407)))));
              reg1432 <= $signed(({reg1422[(1'h1):(1'h0)],
                      {forvar1421[(5'h19):(5'h18)], $unsigned((7'h53))},
                      reg1420} ?
                  $unsigned($unsigned({reg1402,
                      (7'h4f)})) : {((wire1394 * reg1411) + (7'h48)),
                      (reg1402 ? reg1393 : $unsigned(reg1422))}));
              reg1433 <= $signed($unsigned(($signed($unsigned(reg1424)) - (+reg1393))));
              reg1434 = reg1422[(1'h1):(1'h0)];
              reg1435 = reg1415;
            end
          reg1436 <= reg1435[(1'h0):(1'h0)];
          if ($unsigned((|reg1398[(5'h1a):(5'h16)])))
            begin
              reg1437 <= $unsigned($unsigned(reg1395));
              reg1438 <= $unsigned((~&((reg1422 <<< $signed(reg1417)) ?
                  (reg1401 ?
                      (reg1437 || reg1396) : (reg1424 ?
                          (8'ha2) : reg1429)) : forvar1426[(2'h2):(2'h2)])));
              reg1439 <= ({{forvar1428[(4'h8):(2'h2)],
                          {reg1414[(5'h1a):(5'h12)], (8'hbf)}},
                      {$signed($signed(forvar1428))},
                      (-reg1422[(4'ha):(3'h6)])} ?
                  $signed(((wire1389 ? (-reg1415) : (reg1414 < wire1391)) ?
                      $signed((|forvar1428)) : $unsigned((-(8'hbc))))) : $unsigned((reg1432 ?
                      $signed(reg1402) : reg1420[(2'h2):(1'h1)])));
            end
          else
            begin
              reg1437 <= reg1417[(2'h3):(2'h3)];
              reg1440 = ((&($signed((|reg1408)) ?
                  $unsigned(((8'ha4) ^~ reg1404)) : $unsigned((~|reg1403)))) ^~ (~|(~(7'h43))));
              reg1441 = ($signed((wire1389[(5'h10):(4'h8)] ~^ reg1413)) ?
                  (reg1438[(5'h15):(3'h6)] ?
                      wire1394 : $unsigned(wire1391)) : reg1414[(5'h12):(3'h4)]);
            end
          for (forvar1442 = (1'h0); (forvar1442 < (1'h0)); forvar1442 = (forvar1442 + (1'h1)))
            begin
              reg1443 <= reg1403;
              reg1444 = ((|reg1438[(4'ha):(4'ha)]) ?
                  $unsigned($unsigned(((reg1415 | reg1404) ?
                      $unsigned(reg1422) : $signed(reg1398)))) : ($signed($signed((reg1437 >= reg1437))) ?
                      ((reg1408[(2'h3):(2'h3)] ?
                          (!reg1413) : $signed((8'h9d))) <<< $unsigned($unsigned((8'hb2)))) : reg1403[(1'h0):(1'h0)]));
              reg1445 <= $unsigned((reg1410 == (^reg1393)));
            end
          for (forvar1446 = (1'h0); (forvar1446 < (3'h6)); forvar1446 = (forvar1446 + (1'h1)))
            begin
              reg1447 <= $unsigned($signed((reg1411[(5'h17):(4'hb)] == reg1435[(2'h2):(1'h0)])));
              reg1448 <= {$unsigned($unsigned(((reg1435 <<< reg1434) ?
                      (^reg1425) : {reg1424, reg1412}))),
                  ((~&{(forvar1409 ? reg1414 : reg1437),
                      (wire1390 ? wire1388 : reg1433),
                      (wire1391 <<< (7'h56))}) <<< {(reg1414[(4'h9):(3'h6)] ?
                          reg1432[(4'hc):(4'hc)] : (reg1427 >> reg1410)),
                      ((reg1432 < (7'h43)) >= (|reg1434))}),
                  $unsigned(reg1414)};
              reg1449 <= reg1403;
              reg1450 <= (!(forvar1442 - ((reg1436[(2'h3):(1'h0)] ~^ (reg1393 >= reg1434)) ?
                  ((7'h58) || (8'haf)) : reg1422[(4'h8):(2'h3)])));
            end
        end
      reg1451 <= $unsigned($signed(({(reg1447 ? reg1392 : reg1425)} ?
          reg1433[(3'h4):(1'h0)] : ({(8'hb8)} <<< wire1389))));
    end
  always
    @(posedge clk) begin
      reg1452 <= reg1399;
      reg1453 = (+(8'hbe));
      if (((|$unsigned((reg1400 ? $unsigned(reg1401) : reg1443))) ?
          wire1390[(4'h9):(3'h5)] : (+reg1436[(1'h1):(1'h1)])))
        begin
          reg1454 <= $unsigned(wire1390);
          reg1455 <= $signed((-(&($signed((8'hb8)) ?
              $signed(reg1454) : $unsigned((7'h50))))));
          if ((reg1397[(3'h7):(2'h3)] + reg1399[(2'h2):(1'h1)]))
            begin
              reg1456 <= ((((~^reg1448) ?
                      ({reg1450} && (^~reg1430)) : (|(^~reg1392))) ?
                  {reg1422[(3'h7):(1'h1)],
                      reg1450[(2'h3):(1'h1)]} : $unsigned(((reg1415 - (7'h4b)) >> $unsigned(wire1390)))) | $unsigned($unsigned(((reg1448 ^ (8'hbc)) ~^ ((7'h58) ?
                  reg1452 : reg1410)))));
            end
          else
            begin
              reg1457 = (~$signed($unsigned($unsigned((reg1456 >= reg1439)))));
              reg1458 <= ((7'h53) ? reg1396 : wire1394);
              reg1459 = reg1456;
              reg1460 = (|$unsigned((~&reg1399)));
            end
          reg1461 <= reg1416;
        end
      else
        begin
          for (forvar1454 = (1'h0); (forvar1454 < (1'h0)); forvar1454 = (forvar1454 + (1'h1)))
            begin
              reg1457 = reg1438[(5'h1f):(5'h14)];
              reg1459 = (7'h4f);
              reg1460 = ((reg1432 ?
                      ($unsigned((reg1458 ? (8'had) : reg1448)) == ({wire1388,
                              forvar1454,
                              (8'ha5)} ?
                          reg1416 : $unsigned((8'h9e)))) : $unsigned($unsigned(reg1452))) ?
                  $unsigned(reg1450) : ((+((reg1410 ? reg1397 : reg1432) ?
                      reg1459[(5'h10):(1'h1)] : $unsigned(reg1451))) << $unsigned((|$signed((8'ha1))))));
              reg1462 = ((~&reg1458[(3'h5):(1'h0)]) ?
                  {$unsigned(wire1388),
                      reg1461[(4'ha):(3'h6)]} : reg1459[(4'hf):(4'ha)]);
            end
          if ($unsigned({$signed((reg1436[(3'h5):(2'h2)] ?
                  {reg1443, reg1439} : (reg1397 ? (7'h48) : wire1394))),
              reg1410[(5'h15):(5'h12)]}))
            begin
              reg1463 = wire1389;
              reg1464 = $signed((reg1430[(2'h2):(1'h0)] >= $signed((&reg1422[(4'h9):(4'h9)]))));
              reg1465 = $signed($signed($unsigned(({reg1433} ?
                  $signed(reg1399) : (reg1417 ? (7'h52) : (7'h4f))))));
              reg1466 <= $unsigned($unsigned((($unsigned(reg1450) ?
                      (wire1391 + reg1438) : $unsigned(reg1424)) ?
                  reg1452 : {reg1438})));
              reg1467 <= reg1453;
              reg1468 = $unsigned({$unsigned((7'h46))});
              reg1469 = wire1389;
            end
          else
            begin
              reg1463 = $signed((-reg1399[(4'hd):(3'h6)]));
              reg1464 = (+reg1452);
              reg1466 <= (8'hb2);
              reg1467 <= {$unsigned($signed(reg1410[(2'h2):(1'h0)])),
                  (($unsigned((reg1396 ? (7'h4b) : (8'hb4))) ?
                          $unsigned((reg1424 ?
                              (8'h9d) : reg1454)) : {$unsigned(reg1461),
                              $signed((7'h4b))}) ?
                      $signed({reg1417[(1'h0):(1'h0)]}) : ((!$signed(reg1459)) ?
                          (^~reg1439) : $signed((&reg1437))))};
              reg1468 = ($unsigned((&reg1462[(5'h14):(5'h13)])) * (reg1458[(5'h1c):(5'h15)] ?
                  $signed((~|wire1394)) : (~^reg1430)));
            end
        end
    end
  assign wire1470 = (reg1422[(3'h6):(3'h5)] ? reg1454 : $signed((|reg1400)));
  assign wire1471 = $signed($signed($unsigned(reg1397[(3'h4):(1'h1)])));
  assign wire1472 = ($unsigned($signed({(reg1410 > reg1399),
                        (reg1448 ? reg1416 : wire1389)})) >>> reg1456);
  assign wire1473 = (^~{(((wire1389 <= reg1456) > (wire1394 <= (7'h4a))) ?
                            wire1389 : {$signed(reg1417),
                                (reg1424 ? wire1388 : wire1388),
                                (reg1466 ? wire1390 : reg1415)}),
                        reg1448,
                        ($unsigned(reg1449[(5'h17):(4'he)]) - $unsigned($signed(reg1452)))});
  always
    @(posedge clk) begin
      reg1474 = reg1415[(1'h0):(1'h0)];
      reg1475 <= reg1396[(4'hc):(4'hb)];
    end
  assign wire1476 = ($signed(((~|reg1437) == $unsigned(((8'hb3) < reg1401)))) < (8'ha5));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1060
#(parameter param1242 = ((|(~&{(~|(8'ha3)), ((8'hb7) ? (8'hac) : (7'h57)), ((8'hbb) & (8'hb8))})) & (({{(8'h9c), (8'hb2), (8'hbd)}} ? {(~|(8'haf)), {(8'ha3), (7'h50), (8'hb2)}, {(7'h53), (8'ha4)}} : (|{(8'hbf), (8'hb2)})) ? ((((7'h51) ? (8'hb2) : (8'h9f)) ? ((7'h44) ? (8'hbf) : (8'haa)) : ((7'h4b) ^ (8'had))) ? (~^((8'ha9) ? (7'h49) : (8'hb3))) : (^(7'h4f))) : ((((7'h47) != (8'hb5)) ^~ ((8'ha9) <= (8'had))) ? (((7'h4b) ? (8'hab) : (7'h54)) ^ (^(7'h56))) : (((7'h58) ^ (7'h4b)) & (~|(8'ha7)))))), 
parameter param1243 = param1242)
(y, clk, wire1066, wire1065, wire1064, wire1063, wire1062, wire1061);
  output wire [(32'hc84):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire1066;
  input wire [(5'h1c):(1'h0)] wire1065;
  input wire signed [(4'hf):(1'h0)] wire1064;
  input wire [(5'h19):(1'h0)] wire1063;
  input wire [(5'h10):(1'h0)] wire1062;
  input wire [(2'h2):(1'h0)] wire1061;
  wire [(3'h4):(1'h0)] wire1241;
  wire signed [(3'h7):(1'h0)] wire1147;
  wire signed [(3'h7):(1'h0)] wire1067;
  reg [(5'h1d):(1'h0)] reg1240 = (1'h0);
  reg [(4'hb):(1'h0)] reg1239 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1237 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1236 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1234 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1230 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1229 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1226 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1225 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1223 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1222 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1221 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1212 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1216 = (1'h0);
  reg [(4'he):(1'h0)] reg1214 = (1'h0);
  reg [(5'h13):(1'h0)] reg1211 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1209 = (1'h0);
  reg [(5'h18):(1'h0)] reg1205 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1204 = (1'h0);
  reg [(4'h8):(1'h0)] reg1199 = (1'h0);
  reg [(5'h16):(1'h0)] reg1198 = (1'h0);
  reg [(4'hb):(1'h0)] reg1197 = (1'h0);
  reg [(4'hd):(1'h0)] reg1193 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1192 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1190 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1187 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1186 = (1'h0);
  reg [(5'h10):(1'h0)] reg1184 = (1'h0);
  reg [(4'hd):(1'h0)] reg1183 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1182 = (1'h0);
  reg [(5'h14):(1'h0)] reg1180 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1179 = (1'h0);
  reg [(5'h15):(1'h0)] reg1175 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1171 = (1'h0);
  reg [(5'h16):(1'h0)] reg1169 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1168 = (1'h0);
  reg [(3'h5):(1'h0)] reg1165 = (1'h0);
  reg [(5'h16):(1'h0)] reg1163 = (1'h0);
  reg [(4'h8):(1'h0)] reg1161 = (1'h0);
  reg [(5'h14):(1'h0)] reg1160 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1158 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1157 = (1'h0);
  reg [(5'h17):(1'h0)] reg1154 = (1'h0);
  reg [(4'hb):(1'h0)] reg1151 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1144 = (1'h0);
  reg [(5'h19):(1'h0)] reg1140 = (1'h0);
  reg [(4'hc):(1'h0)] reg1138 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1136 = (1'h0);
  reg [(5'h15):(1'h0)] reg1134 = (1'h0);
  reg [(3'h4):(1'h0)] reg1133 = (1'h0);
  reg [(3'h5):(1'h0)] reg1129 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1126 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1125 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1123 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1122 = (1'h0);
  reg [(3'h4):(1'h0)] reg1121 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1120 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1117 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1111 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1105 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1104 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1101 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1100 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1099 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1097 = (1'h0);
  reg [(3'h7):(1'h0)] reg1092 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1091 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1090 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1089 = (1'h0);
  reg [(4'h8):(1'h0)] reg1087 = (1'h0);
  reg [(4'hd):(1'h0)] reg1085 = (1'h0);
  reg [(5'h17):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1081 = (1'h0);
  reg [(4'hf):(1'h0)] reg1079 = (1'h0);
  reg [(5'h15):(1'h0)] reg1078 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1076 = (1'h0);
  reg [(3'h7):(1'h0)] reg1075 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1074 = (1'h0);
  reg [(3'h7):(1'h0)] reg1073 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1071 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1070 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1232 = (1'h0);
  reg [(5'h19):(1'h0)] reg1231 = (1'h0);
  reg [(4'ha):(1'h0)] reg1238 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1235 = (1'h0);
  reg [(2'h3):(1'h0)] reg1233 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1232 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1231 = (1'h0);
  reg [(5'h18):(1'h0)] reg1228 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1227 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1224 = (1'h0);
  reg [(5'h13):(1'h0)] reg1220 = (1'h0);
  reg [(4'h9):(1'h0)] reg1219 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1218 = (1'h0);
  reg [(4'h8):(1'h0)] reg1217 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1216 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1205 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1215 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1213 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1212 = (1'h0);
  reg [(4'h9):(1'h0)] reg1210 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1208 = (1'h0);
  reg [(3'h7):(1'h0)] reg1207 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1206 = (1'h0);
  reg [(5'h13):(1'h0)] reg1203 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1202 = (1'h0);
  reg [(4'h9):(1'h0)] reg1201 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1200 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1196 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1195 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1194 = (1'h0);
  reg [(5'h16):(1'h0)] reg1191 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1189 = (1'h0);
  reg [(3'h4):(1'h0)] reg1188 = (1'h0);
  reg [(5'h18):(1'h0)] reg1185 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1176 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1169 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1181 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1178 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1177 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1176 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1174 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1173 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1172 = (1'h0);
  reg [(5'h12):(1'h0)] reg1170 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1167 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1166 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1164 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1162 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1159 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1156 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1155 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1153 = (1'h0);
  reg [(4'hf):(1'h0)] reg1152 = (1'h0);
  reg [(4'ha):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1149 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1148 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1146 = (1'h0);
  reg [(4'h8):(1'h0)] reg1145 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1143 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1142 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1141 = (1'h0);
  reg [(5'h15):(1'h0)] reg1139 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1137 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1135 = (1'h0);
  reg [(5'h19):(1'h0)] reg1132 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1131 = (1'h0);
  reg [(2'h3):(1'h0)] reg1130 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1128 = (1'h0);
  reg [(5'h19):(1'h0)] reg1127 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1124 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1113 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1119 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1118 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1117 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1116 = (1'h0);
  reg [(5'h11):(1'h0)] reg1115 = (1'h0);
  reg [(2'h3):(1'h0)] reg1114 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1113 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1112 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1110 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1109 = (1'h0);
  reg [(3'h6):(1'h0)] reg1108 = (1'h0);
  reg [(2'h2):(1'h0)] reg1107 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1106 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1103 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1102 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1098 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1096 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1095 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1094 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1093 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1088 = (1'h0);
  reg [(4'h9):(1'h0)] reg1086 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1083 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1082 = (1'h0);
  reg [(5'h12):(1'h0)] reg1080 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1077 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1072 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1069 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1068 = (1'h0);
  assign y = {wire1241,
                 wire1147,
                 wire1067,
                 reg1240,
                 reg1239,
                 reg1237,
                 reg1236,
                 reg1234,
                 reg1230,
                 reg1229,
                 reg1226,
                 reg1225,
                 reg1223,
                 reg1222,
                 reg1221,
                 reg1212,
                 reg1216,
                 reg1214,
                 reg1211,
                 reg1209,
                 reg1205,
                 reg1204,
                 reg1199,
                 reg1198,
                 reg1197,
                 reg1193,
                 reg1192,
                 reg1190,
                 reg1187,
                 reg1186,
                 reg1184,
                 reg1183,
                 reg1182,
                 reg1180,
                 reg1179,
                 reg1175,
                 reg1171,
                 reg1169,
                 reg1168,
                 reg1165,
                 reg1163,
                 reg1161,
                 reg1160,
                 reg1158,
                 reg1157,
                 reg1154,
                 reg1151,
                 reg1144,
                 reg1140,
                 reg1138,
                 reg1136,
                 reg1134,
                 reg1133,
                 reg1129,
                 reg1126,
                 reg1125,
                 reg1123,
                 reg1122,
                 reg1121,
                 reg1120,
                 reg1117,
                 reg1111,
                 reg1105,
                 reg1104,
                 reg1101,
                 reg1100,
                 reg1099,
                 reg1097,
                 reg1092,
                 reg1091,
                 reg1090,
                 reg1089,
                 reg1087,
                 reg1085,
                 reg1084,
                 reg1081,
                 reg1079,
                 reg1078,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1073,
                 reg1071,
                 reg1070,
                 forvar1232,
                 reg1231,
                 reg1238,
                 reg1235,
                 reg1233,
                 reg1232,
                 forvar1231,
                 reg1228,
                 reg1227,
                 reg1224,
                 reg1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 forvar1216,
                 forvar1205,
                 reg1215,
                 reg1213,
                 forvar1212,
                 reg1210,
                 reg1208,
                 reg1207,
                 reg1206,
                 reg1203,
                 reg1202,
                 reg1201,
                 reg1200,
                 reg1196,
                 reg1195,
                 reg1194,
                 reg1191,
                 reg1189,
                 reg1188,
                 reg1185,
                 forvar1176,
                 forvar1169,
                 reg1181,
                 forvar1178,
                 reg1177,
                 reg1176,
                 reg1174,
                 reg1173,
                 reg1172,
                 reg1170,
                 reg1167,
                 forvar1166,
                 reg1164,
                 reg1162,
                 reg1159,
                 forvar1156,
                 reg1155,
                 reg1153,
                 reg1152,
                 reg1150,
                 forvar1149,
                 forvar1148,
                 reg1146,
                 reg1145,
                 reg1143,
                 reg1142,
                 reg1141,
                 reg1139,
                 reg1137,
                 reg1135,
                 reg1132,
                 reg1131,
                 reg1130,
                 forvar1128,
                 reg1127,
                 reg1124,
                 reg1113,
                 reg1119,
                 reg1118,
                 forvar1117,
                 reg1116,
                 reg1115,
                 reg1114,
                 forvar1113,
                 reg1112,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1107,
                 reg1106,
                 reg1103,
                 reg1102,
                 reg1098,
                 reg1096,
                 reg1095,
                 reg1094,
                 reg1093,
                 reg1088,
                 reg1086,
                 reg1083,
                 forvar1082,
                 reg1080,
                 reg1077,
                 reg1072,
                 forvar1069,
                 reg1068,
                 (1'h0)};
  assign wire1067 = $unsigned(wire1063[(5'h10):(4'hf)]);
  always
    @(posedge clk) begin
      reg1068 = $signed($unsigned((|$signed(wire1063[(5'h17):(3'h4)]))));
      for (forvar1069 = (1'h0); (forvar1069 < (3'h4)); forvar1069 = (forvar1069 + (1'h1)))
        begin
          reg1070 <= (wire1067[(1'h1):(1'h1)] && (wire1065 == ($signed((wire1067 ^ wire1061)) ?
              ((wire1067 <= wire1063) ?
                  (wire1067 ?
                      wire1064 : wire1066) : $signed(reg1068)) : {(wire1063 ?
                      forvar1069 : wire1064),
                  (~^wire1067),
                  ((7'h57) <= reg1068)})));
          reg1071 <= $signed($unsigned((!(~wire1066[(1'h1):(1'h1)]))));
          reg1072 = $unsigned((~&((~^(reg1068 != wire1064)) || (^~$signed(wire1061)))));
          reg1073 <= (~&(wire1061[(1'h1):(1'h0)] ?
              (7'h40) : ($unsigned({(8'hb9),
                  reg1072,
                  wire1061}) || ($signed(wire1063) ?
                  (-wire1067) : $unsigned(reg1070)))));
          reg1074 <= (~^({(~(wire1066 ? forvar1069 : reg1068)),
                  ($signed(forvar1069) ?
                      reg1068[(5'h13):(3'h4)] : $signed(reg1072)),
                  (reg1071[(5'h15):(2'h2)] >= (|(7'h48)))} ?
              $signed((+{reg1073,
                  reg1068})) : $unsigned((^~$unsigned(wire1065)))));
          if ($signed($unsigned($unsigned(forvar1069[(4'hf):(4'hf)]))))
            begin
              reg1075 <= reg1071;
            end
          else
            begin
              reg1075 <= $signed((~&$unsigned($unsigned(wire1067[(3'h6):(3'h5)]))));
              reg1076 <= ($signed(reg1071) < wire1063[(5'h14):(5'h14)]);
              reg1077 = ({reg1071[(5'h13):(4'h9)],
                  reg1076,
                  ((!$signed(reg1071)) ?
                      ((^wire1067) ?
                          wire1066[(2'h3):(2'h2)] : (~|(7'h51))) : wire1066)} && (!wire1065[(4'hb):(4'h9)]));
              reg1078 <= wire1061[(1'h1):(1'h1)];
              reg1079 <= $unsigned(reg1068);
              reg1080 = reg1079[(4'h9):(3'h6)];
              reg1081 <= (({{$unsigned(wire1067)},
                      $signed(reg1076[(5'h11):(3'h5)]),
                      (reg1077[(4'he):(1'h0)] ?
                          (!wire1067) : (wire1067 * reg1078))} ^~ $unsigned(reg1068)) ?
                  $signed((wire1062 + $signed(reg1068[(4'h8):(3'h7)]))) : $unsigned(wire1067[(3'h7):(1'h0)]));
            end
        end
      for (forvar1082 = (1'h0); (forvar1082 < (2'h3)); forvar1082 = (forvar1082 + (1'h1)))
        begin
          reg1083 = {($signed(wire1061) ?
                  (+(8'hb9)) : {(~&{reg1076, forvar1082, reg1073}),
                      ((reg1072 ? wire1066 : reg1074) ?
                          $signed(reg1080) : reg1081)}),
              wire1062[(4'ha):(3'h6)],
              {{{(~|wire1067), (7'h47)}}}};
          reg1084 <= (reg1079[(2'h3):(2'h2)] & $unsigned($unsigned($unsigned((reg1070 * reg1068)))));
          reg1085 <= $signed({reg1079});
          if ((reg1084[(3'h5):(1'h1)] ?
              ($unsigned($signed((8'had))) ?
                  $signed(({reg1081,
                      wire1067,
                      reg1070} & reg1071[(4'he):(1'h0)])) : reg1085) : (($signed(wire1064[(4'hd):(4'hb)]) ?
                      (~((8'h9d) ? wire1065 : (8'hba))) : (~|(reg1076 ?
                          reg1073 : wire1064))) ?
                  $signed((-(|(8'hbb)))) : $signed(($signed(reg1068) ?
                      (-reg1077) : $signed(wire1064))))))
            begin
              reg1086 = (($signed(wire1064) < $signed($unsigned(reg1076[(2'h2):(1'h1)]))) ?
                  wire1063[(3'h4):(1'h0)] : $signed(wire1067));
              reg1087 <= wire1063[(2'h3):(1'h1)];
              reg1088 = reg1074[(3'h7):(1'h0)];
              reg1089 <= reg1080;
              reg1090 <= $unsigned({$unsigned(reg1086[(3'h6):(2'h3)]),
                  $unsigned(reg1068[(5'h16):(4'he)]),
                  {(~|{reg1089, (7'h47), wire1065}),
                      $unsigned($signed(wire1063))}});
            end
          else
            begin
              reg1087 <= reg1070;
              reg1089 <= ({$unsigned(reg1075),
                  $unsigned(((reg1084 ? reg1090 : reg1074) * wire1065)),
                  wire1063} & ($unsigned($unsigned(reg1084)) ?
                  reg1073 : $signed((-reg1071))));
              reg1090 <= reg1080[(5'h11):(4'h8)];
              reg1091 <= (wire1061 ?
                  reg1072 : (reg1076 >>> $unsigned((reg1068 ?
                      wire1064 : reg1081[(3'h5):(1'h0)]))));
              reg1092 <= ((wire1061 < (7'h4b)) ?
                  wire1064[(4'hc):(2'h3)] : {($signed($unsigned(wire1061)) ?
                          reg1088[(5'h1f):(5'h1f)] : (8'haf)),
                      $unsigned(reg1079[(2'h3):(1'h0)]),
                      reg1081});
              reg1093 = (8'h9f);
              reg1094 = $signed({reg1091[(5'h14):(5'h10)]});
            end
          if (reg1087)
            begin
              reg1095 = {$signed(reg1077[(1'h0):(1'h0)]),
                  reg1081[(3'h4):(2'h2)]};
              reg1096 = $signed((wire1064 ^ {$unsigned(reg1088[(5'h11):(3'h7)]),
                  $signed(reg1093)}));
              reg1097 <= wire1066;
              reg1098 = $signed($unsigned($unsigned(((!reg1074) > reg1091[(4'hb):(4'h8)]))));
              reg1099 <= reg1091;
              reg1100 <= (^$unsigned($unsigned($unsigned(reg1094))));
              reg1101 <= (!(&$signed(((wire1064 != (7'h56)) && (~&wire1066)))));
            end
          else
            begin
              reg1095 = $signed($unsigned($signed($unsigned(((8'had) << reg1074)))));
              reg1096 = (((8'hb1) ?
                      ((-reg1083[(4'hf):(4'ha)]) >>> {(reg1080 ?
                              reg1076 : reg1071)}) : (7'h41)) ?
                  (reg1073 * (^~(((8'ha9) ?
                      reg1089 : (7'h43)) & reg1071[(1'h0):(1'h0)]))) : ($unsigned($unsigned($signed(reg1086))) > {((reg1068 ?
                              reg1068 : forvar1069) ?
                          $unsigned(reg1084) : $unsigned(wire1067))}));
              reg1097 <= wire1061;
              reg1098 = $signed((!$signed($signed(wire1063[(2'h3):(2'h3)]))));
              reg1102 = reg1080;
              reg1103 = reg1090[(5'h18):(5'h17)];
            end
          if ($signed(wire1065[(3'h7):(3'h5)]))
            begin
              reg1104 <= reg1086[(3'h5):(3'h4)];
              reg1105 <= $unsigned(($unsigned(($signed(reg1087) ?
                  reg1103[(4'hc):(3'h5)] : reg1090[(5'h10):(1'h0)])) * (reg1083[(4'h9):(1'h1)] - reg1077)));
            end
          else
            begin
              reg1106 = (+$unsigned((8'haf)));
              reg1107 = (!(~&(^~(~^(reg1095 >>> reg1095)))));
              reg1108 = $unsigned($signed(wire1064[(4'he):(4'hd)]));
              reg1109 = reg1100;
              reg1110 = reg1100[(3'h5):(1'h0)];
            end
        end
      reg1111 <= (~$unsigned(((reg1070 <<< {reg1094}) ?
          ((reg1106 <= reg1079) ?
              {reg1102,
                  reg1081} : (reg1103 | reg1090)) : reg1105[(4'he):(2'h2)])));
      reg1112 = (!(reg1087 <= reg1076));
      if ((!reg1099[(5'h13):(4'hf)]))
        begin
          for (forvar1113 = (1'h0); (forvar1113 < (1'h1)); forvar1113 = (forvar1113 + (1'h1)))
            begin
              reg1114 = wire1066;
              reg1115 = (-$signed(((reg1070[(3'h4):(1'h0)] ?
                      (reg1092 == reg1106) : (reg1096 || wire1063)) ?
                  (~&reg1083[(3'h5):(2'h2)]) : ((reg1077 ? reg1083 : reg1090) ?
                      $unsigned(wire1063) : (reg1088 || forvar1082)))));
              reg1116 = ((&(((reg1110 >> reg1109) ?
                          {reg1090, reg1115} : reg1099[(5'h1a):(5'h18)]) ?
                      {{reg1114},
                          ((8'haa) ? forvar1082 : wire1062),
                          (~|(8'hb1))} : ((reg1071 + (7'h47)) != (-(8'h9c))))) ?
                  reg1112 : $unsigned($unsigned($signed($unsigned(reg1096)))));
            end
          for (forvar1117 = (1'h0); (forvar1117 < (1'h1)); forvar1117 = (forvar1117 + (1'h1)))
            begin
              reg1118 = reg1106;
            end
          reg1119 = $unsigned(($signed($signed(reg1103[(5'h1a):(5'h18)])) ?
              $signed((8'hac)) : reg1072[(1'h0):(1'h0)]));
        end
      else
        begin
          if (((+reg1115) ?
              (reg1074[(5'h12):(2'h2)] != (7'h47)) : ($unsigned($unsigned((^wire1066))) & ($unsigned(wire1061[(2'h2):(1'h1)]) ?
                  ((!reg1118) >= wire1063) : (!reg1100[(1'h1):(1'h0)])))))
            begin
              reg1113 = (wire1061 ?
                  $signed($unsigned(reg1093[(3'h7):(1'h1)])) : (^$signed({(reg1077 > reg1071),
                      (reg1096 & reg1070),
                      forvar1069[(4'ha):(2'h2)]})));
              reg1114 = $signed({(((^~(7'h49)) ? reg1108 : wire1065) ?
                      reg1113[(4'hc):(1'h0)] : (-reg1100[(2'h3):(1'h0)])),
                  $signed((^~forvar1117))});
              reg1117 <= $signed((|$signed(($signed((8'hbe)) >= wire1061[(1'h0):(1'h0)]))));
              reg1118 = {$signed($unsigned(($unsigned(reg1085) ?
                      ((8'hbf) ? reg1103 : reg1071) : (reg1075 ^~ wire1061)))),
                  $signed((((reg1114 ? reg1073 : reg1099) ?
                      wire1063 : (reg1099 ?
                          reg1100 : (7'h43))) != (~|$signed((8'hbb)))))};
              reg1119 = {reg1097,
                  ((({reg1079, (8'ha8)} | $unsigned(reg1093)) ?
                          ($unsigned(reg1109) <= (~reg1071)) : reg1106) ?
                      reg1110 : $unsigned(($unsigned(reg1108) ?
                          {(8'ha1), reg1113, reg1106} : $signed(wire1063)))),
                  reg1116[(4'he):(4'hb)]};
            end
          else
            begin
              reg1117 <= $unsigned(reg1093[(5'h13):(1'h1)]);
              reg1118 = $unsigned(reg1088);
              reg1120 <= $unsigned($unsigned(wire1066[(4'hc):(4'h9)]));
            end
          if (reg1078[(4'h9):(1'h0)])
            begin
              reg1121 <= ((+wire1067) ? reg1085 : (^$unsigned((~|(!(7'h41))))));
              reg1122 <= ($unsigned(wire1066[(4'hc):(3'h4)]) <<< $signed(($unsigned((reg1092 <= reg1084)) <= reg1075)));
              reg1123 <= forvar1113[(5'h11):(4'hc)];
            end
          else
            begin
              reg1124 = $signed($unsigned((~$unsigned(reg1070[(3'h4):(1'h1)]))));
              reg1125 <= reg1083[(3'h4):(2'h3)];
              reg1126 <= $signed($signed((~{reg1084[(4'hc):(3'h4)],
                  (~^(7'h46))})));
              reg1127 = $signed($unsigned(reg1088[(4'hd):(4'ha)]));
            end
          for (forvar1128 = (1'h0); (forvar1128 < (1'h1)); forvar1128 = (forvar1128 + (1'h1)))
            begin
              reg1129 <= {$unsigned($unsigned(reg1124))};
              reg1130 = reg1114[(1'h1):(1'h1)];
              reg1131 = $signed($signed({reg1119[(1'h0):(1'h0)],
                  $unsigned(reg1110),
                  $signed($unsigned(reg1081))}));
              reg1132 = reg1122[(5'h1b):(4'hd)];
              reg1133 <= (~({$unsigned(reg1081[(4'hd):(4'hb)])} || $unsigned(($signed(reg1070) != reg1087[(3'h5):(3'h4)]))));
            end
          reg1134 <= ($signed(({wire1065,
                  $unsigned(wire1063),
                  reg1118[(1'h1):(1'h0)]} ^~ reg1070[(4'hc):(1'h1)])) ?
              (((7'h56) ?
                      (reg1076[(5'h1b):(2'h3)] ?
                          (reg1118 & reg1075) : $unsigned(reg1088)) : reg1070) ?
                  $signed($unsigned(reg1084[(4'ha):(4'h8)])) : (^~(^(^reg1088)))) : $signed(reg1105));
          if (({$unsigned(($unsigned(reg1102) || reg1095)),
                  ({$unsigned(reg1094),
                      $unsigned(reg1131)} || (reg1089 && $signed(wire1063)))} ?
              {$signed(reg1102[(4'hd):(3'h4)]),
                  ((~|(~|(7'h56))) ?
                      ($signed(reg1125) > (reg1115 << reg1068)) : reg1078)} : (reg1123 ?
                  reg1115[(2'h3):(1'h1)] : reg1122[(5'h1b):(5'h1b)])))
            begin
              reg1135 = $unsigned(reg1086[(2'h3):(1'h1)]);
              reg1136 <= (|$unsigned($signed($signed($signed(reg1086)))));
              reg1137 = reg1097[(1'h1):(1'h0)];
              reg1138 <= reg1098[(5'h10):(2'h2)];
              reg1139 = (~&reg1122[(4'hc):(4'hb)]);
              reg1140 <= reg1102[(4'hf):(1'h0)];
            end
          else
            begin
              reg1135 = (~{(^reg1108),
                  (reg1081[(2'h2):(1'h1)] ?
                      ({(7'h41), wire1065, reg1114} ?
                          (~&(7'h58)) : $unsigned((8'haa))) : reg1085),
                  $signed(reg1092[(3'h7):(1'h0)])});
              reg1136 <= (^((&((^wire1062) ?
                  (^reg1111) : $unsigned(reg1081))) < $signed(($unsigned(reg1085) ^~ (7'h4f)))));
              reg1137 = forvar1117[(5'h14):(1'h0)];
              reg1138 <= reg1083;
              reg1140 <= reg1119;
              reg1141 = {({wire1067} ?
                      $unsigned($unsigned(reg1083[(4'hd):(3'h4)])) : reg1116[(3'h4):(2'h3)])};
              reg1142 = {$unsigned({(((7'h48) ?
                          (8'hbd) : reg1086) << {wire1062})}),
                  $signed(reg1139[(3'h6):(1'h1)]),
                  {({(~|wire1061), (+reg1139)} ?
                          ((forvar1117 != reg1074) ?
                              (reg1141 ?
                                  reg1086 : reg1121) : (8'hb1)) : $unsigned((reg1124 > reg1103))),
                      ((7'h4f) <<< $unsigned((+reg1134)))}};
            end
          reg1143 = reg1137;
          if ({$unsigned(((((8'ha0) ? reg1129 : reg1134) ?
                  reg1091[(4'h8):(2'h3)] : (wire1061 ?
                      (7'h4c) : (8'ha7))) << forvar1069))})
            begin
              reg1144 <= ($unsigned(({$unsigned(reg1078)} ?
                  (~reg1076[(5'h12):(2'h2)]) : ((+reg1139) ?
                      {reg1098} : reg1138[(3'h6):(3'h4)]))) << reg1142);
              reg1145 = reg1112;
            end
          else
            begin
              reg1145 = wire1061;
              reg1146 = reg1084[(4'he):(4'ha)];
            end
        end
    end
  assign wire1147 = wire1063;
  always
    @(posedge clk) begin
      for (forvar1148 = (1'h0); (forvar1148 < (1'h1)); forvar1148 = (forvar1148 + (1'h1)))
        begin
          for (forvar1149 = (1'h0); (forvar1149 < (2'h2)); forvar1149 = (forvar1149 + (1'h1)))
            begin
              reg1150 = (reg1092[(2'h3):(2'h2)] - reg1070[(4'hf):(4'h8)]);
              reg1151 <= (~reg1074);
              reg1152 = (reg1151 ?
                  (reg1099 ?
                      reg1073 : wire1067[(3'h4):(1'h1)]) : (!reg1100[(3'h4):(1'h1)]));
              reg1153 = $unsigned((~reg1121));
              reg1154 <= (reg1111[(1'h0):(1'h0)] ? (~(~|(8'h9d))) : reg1091);
              reg1155 = $signed((^$signed((|reg1140))));
            end
          for (forvar1156 = (1'h0); (forvar1156 < (1'h0)); forvar1156 = (forvar1156 + (1'h1)))
            begin
              reg1157 <= ($signed(wire1063[(3'h6):(3'h5)]) && (~^$signed((|(8'hae)))));
              reg1158 <= $unsigned($signed(reg1085));
              reg1159 = reg1074;
              reg1160 <= ((-(~$unsigned({reg1074, reg1071, reg1071}))) ?
                  ($signed((8'haf)) ?
                      $unsigned(reg1079) : $unsigned((-(~reg1091)))) : ($unsigned(reg1123) == (($signed(reg1081) ?
                          {reg1085, reg1138} : {forvar1148, reg1071}) ?
                      reg1090[(3'h6):(3'h6)] : ((&(8'ha0)) ?
                          (reg1155 <= reg1129) : (-reg1126)))));
            end
          reg1161 <= ((reg1134 > $signed(reg1071[(5'h10):(3'h6)])) > {(reg1136[(1'h0):(1'h0)] >> (!reg1111))});
          if ($unsigned(reg1158))
            begin
              reg1162 = reg1126[(3'h5):(3'h5)];
              reg1163 <= ({$unsigned($unsigned((7'h53))),
                      (~reg1134[(4'hc):(4'hb)])} ?
                  reg1151 : $unsigned(wire1067[(3'h6):(2'h2)]));
              reg1164 = $unsigned($unsigned(reg1076[(4'h9):(3'h4)]));
            end
          else
            begin
              reg1162 = wire1066;
            end
          reg1165 <= (reg1070[(1'h1):(1'h1)] ?
              reg1081[(4'hf):(3'h5)] : reg1074);
          for (forvar1166 = (1'h0); (forvar1166 < (2'h3)); forvar1166 = (forvar1166 + (1'h1)))
            begin
              reg1167 = (~|($unsigned(($unsigned(reg1152) ?
                  (reg1161 ?
                      reg1092 : reg1125) : $signed(reg1165))) >>> (+(&reg1159[(5'h15):(3'h4)]))));
            end
        end
      reg1168 <= ((!(^~$signed($signed(reg1079)))) ?
          $signed(reg1129) : (-((^$signed(reg1099)) ?
              reg1157[(5'h17):(5'h17)] : $signed((reg1120 << reg1144)))));
      if (((($signed($signed(reg1133)) ? reg1160 : reg1125) ?
              reg1154[(4'ha):(3'h4)] : $unsigned((!(8'hb6)))) ?
          (($signed($signed(reg1165)) | ((-reg1087) << $signed(reg1133))) * ($signed((|reg1168)) & ((~(7'h4d)) ?
              wire1062 : (!reg1120)))) : ($signed($unsigned($unsigned(reg1158))) ?
              (^~({reg1151, reg1160} ?
                  reg1159[(4'hf):(1'h1)] : {reg1087})) : forvar1149[(4'ha):(1'h1)])))
        begin
          if ((($unsigned(((^~reg1105) ?
              (reg1144 ?
                  reg1165 : reg1151) : reg1079[(4'ha):(2'h2)])) - ($signed((reg1163 != reg1105)) ?
              {$unsigned((8'hb1)),
                  $unsigned(reg1167)} : {reg1125[(2'h3):(1'h1)]})) | wire1063[(4'hc):(4'ha)]))
            begin
              reg1169 <= (&(reg1076 ?
                  ((~&$unsigned(reg1099)) << (reg1140 >= (~(8'hb0)))) : (reg1104 - $signed(reg1138))));
              reg1170 = reg1084;
              reg1171 <= {$signed(({(reg1101 - reg1076), {wire1147, reg1105}} ?
                      $signed((reg1074 ?
                          reg1168 : (7'h4c))) : $signed(reg1100))),
                  ((-((reg1144 ? reg1151 : forvar1166) ?
                          reg1162[(5'h12):(4'h9)] : {forvar1148,
                              wire1067,
                              reg1150})) ?
                      (+(~$signed(reg1101))) : (+($unsigned(reg1075) > reg1158[(2'h3):(2'h2)]))),
                  reg1152};
            end
          else
            begin
              reg1170 = $unsigned(reg1099[(3'h5):(1'h1)]);
              reg1172 = ($unsigned({reg1117[(2'h2):(1'h0)]}) && (($signed(reg1122[(4'he):(3'h7)]) - reg1099[(5'h18):(4'hc)]) ?
                  reg1081[(1'h1):(1'h0)] : ($signed(reg1155) ?
                      (reg1075[(3'h6):(3'h6)] * (|(8'hba))) : (~|(reg1164 ?
                          reg1153 : wire1063)))));
              reg1173 = $unsigned(forvar1148);
              reg1174 = (reg1168[(3'h4):(1'h1)] + $unsigned(forvar1166[(4'hc):(3'h7)]));
              reg1175 <= reg1099;
              reg1176 = wire1147[(3'h4):(2'h3)];
              reg1177 = (7'h41);
            end
          for (forvar1178 = (1'h0); (forvar1178 < (2'h3)); forvar1178 = (forvar1178 + (1'h1)))
            begin
              reg1179 <= $signed((~|reg1087));
              reg1180 <= $unsigned(reg1105[(5'h13):(4'he)]);
              reg1181 = (^~((((|reg1071) << (reg1159 ?
                  reg1150 : reg1120)) - reg1180) << reg1164));
            end
        end
      else
        begin
          for (forvar1169 = (1'h0); (forvar1169 < (3'h5)); forvar1169 = (forvar1169 + (1'h1)))
            begin
              reg1171 <= $signed($unsigned(reg1089));
              reg1172 = $unsigned($unsigned(reg1167[(1'h1):(1'h0)]));
              reg1175 <= $unsigned(reg1170[(4'hf):(2'h3)]);
            end
          for (forvar1176 = (1'h0); (forvar1176 < (3'h4)); forvar1176 = (forvar1176 + (1'h1)))
            begin
              reg1177 = (~|((reg1081[(4'hb):(4'h8)] < reg1175) != $signed($signed($unsigned(reg1071)))));
            end
          for (forvar1178 = (1'h0); (forvar1178 < (1'h0)); forvar1178 = (forvar1178 + (1'h1)))
            begin
              reg1181 = ({{(reg1158[(1'h0):(1'h0)] << (reg1174 < reg1071))},
                  (-{reg1151[(4'h9):(3'h4)]})} < $unsigned((7'h58)));
              reg1182 <= ((reg1089 ?
                  reg1162[(1'h0):(1'h0)] : (~&$signed((wire1063 ?
                      reg1177 : reg1155)))) ~^ {(|$signed((reg1079 ?
                      reg1078 : wire1063)))});
              reg1183 <= {((~^$unsigned((reg1159 ? (8'ha0) : reg1090))) ?
                      ($signed(wire1066) ?
                          (reg1122[(5'h10):(3'h7)] >> ((7'h49) <<< reg1085)) : forvar1148) : reg1167[(1'h1):(1'h0)]),
                  $signed((reg1074[(5'h12):(1'h0)] ?
                      reg1129[(2'h3):(2'h2)] : (8'h9d))),
                  {($unsigned(reg1122) ?
                          reg1179[(3'h5):(3'h5)] : $signed({reg1157}))}};
              reg1184 <= $unsigned({($signed(((7'h53) - reg1179)) ?
                      reg1100 : wire1064[(3'h6):(3'h6)]),
                  $signed((((7'h58) ? reg1172 : reg1105) ?
                      (reg1167 ? reg1092 : reg1123) : forvar1166)),
                  (&$signed((reg1172 ? reg1168 : reg1165)))});
              reg1185 = ($signed(reg1171[(5'h10):(2'h3)]) ?
                  (&{{{reg1111, reg1151}, $signed(reg1162)}}) : reg1081);
            end
          if ((reg1097[(1'h1):(1'h0)] != ((8'hb3) ?
              $signed(({wire1061,
                  (7'h42)} >>> $signed((8'ha3)))) : (~(!(~forvar1148))))))
            begin
              reg1186 <= (((reg1079[(2'h3):(1'h1)] ?
                      (~|$unsigned(reg1183)) : ({wire1067} ?
                          (~reg1168) : (8'ha2))) ?
                  reg1157[(3'h7):(3'h6)] : $unsigned(($signed(reg1087) ^ (8'hbe)))) & $signed(reg1167[(1'h0):(1'h0)]));
              reg1187 <= $signed(((!$unsigned(forvar1156[(3'h4):(2'h3)])) >> ((reg1152[(4'hc):(4'ha)] ?
                  $signed(wire1067) : reg1140[(4'hb):(2'h2)]) && (^(wire1061 ?
                  (7'h46) : reg1179)))));
              reg1188 = reg1099[(4'h9):(3'h7)];
            end
          else
            begin
              reg1186 <= (~&(reg1117 ?
                  ($signed((reg1175 ? reg1158 : reg1117)) ?
                      reg1171[(4'h9):(3'h6)] : reg1129[(2'h2):(2'h2)]) : reg1133[(1'h0):(1'h0)]));
              reg1188 = ({(((reg1074 != (8'ha7)) ?
                          reg1155[(5'h12):(3'h7)] : (^(8'haa))) * (~^{reg1186,
                          reg1169})),
                      ((~^$signed(forvar1176)) ?
                          reg1097[(2'h3):(1'h0)] : $signed((wire1067 ?
                              reg1154 : (8'hb6))))} ?
                  reg1170[(3'h7):(3'h5)] : $signed((^~reg1161[(4'h8):(3'h6)])));
              reg1189 = $unsigned(((|reg1085[(4'h9):(1'h1)]) ?
                  $signed($unsigned(forvar1176)) : reg1174));
              reg1190 <= ($signed($unsigned(reg1187)) ?
                  (!(!$unsigned($unsigned((7'h4a))))) : ($unsigned(reg1167) ?
                      $signed((reg1073[(1'h0):(1'h0)] >>> {reg1136,
                          reg1111,
                          (8'ha4)})) : forvar1176[(4'h8):(1'h0)]));
              reg1191 = $unsigned((^~reg1126[(2'h3):(1'h0)]));
              reg1192 <= (-reg1101[(4'he):(3'h7)]);
            end
          if ((reg1075[(1'h0):(1'h0)] ?
              reg1182 : $signed($unsigned(({reg1134, reg1085} ?
                  forvar1149 : $signed(wire1062))))))
            begin
              reg1193 <= (+$signed((reg1182 >> reg1188[(1'h1):(1'h1)])));
              reg1194 = (({(~&(~&reg1179))} ?
                      $unsigned((!(reg1121 ?
                          reg1175 : reg1140))) : $signed($signed(((8'haf) ?
                          reg1144 : reg1136)))) ?
                  reg1073 : (reg1172 <= (reg1079 ^ (8'h9c))));
              reg1195 = (reg1101 ^~ reg1185[(4'hb):(3'h7)]);
            end
          else
            begin
              reg1193 <= $unsigned(((!(reg1185 == (|reg1071))) & reg1076));
            end
          if (reg1184)
            begin
              reg1196 = reg1111[(1'h1):(1'h1)];
              reg1197 <= wire1065[(4'hb):(4'hb)];
              reg1198 <= $unsigned({((^~(reg1175 || reg1197)) && (((8'hbf) ?
                      reg1144 : reg1179) <= reg1144)),
                  forvar1156});
              reg1199 <= $unsigned((&(^~reg1185[(5'h14):(3'h7)])));
            end
          else
            begin
              reg1197 <= (~(($unsigned(reg1117[(5'h13):(3'h7)]) ^ {reg1078[(1'h0):(1'h0)],
                      $signed(reg1081)}) ?
                  reg1155[(4'hb):(4'h8)] : {(reg1176 ?
                          (!reg1159) : {(7'h4a), reg1198}),
                      (^(reg1198 >> reg1085)),
                      ($unsigned(reg1155) ? reg1144 : $unsigned(reg1170))}));
            end
        end
      if ((({((^reg1164) ? (reg1153 ? reg1122 : reg1188) : $unsigned(wire1066)),
              $unsigned((!reg1158))} ?
          wire1064[(4'h9):(2'h3)] : $unsigned((7'h53))) < $signed(((-reg1121) ^ $unsigned(((8'hbb) ?
          reg1157 : reg1122))))))
        begin
          if ((!forvar1178[(3'h5):(2'h2)]))
            begin
              reg1200 = (reg1194 ?
                  (($unsigned(reg1092) ? reg1151 : (^~reg1182[(3'h6):(3'h6)])) ?
                      ((((8'hb5) * (8'hae)) ?
                          (reg1165 != reg1079) : $signed((8'hb6))) >>> reg1070[(3'h6):(2'h2)]) : reg1117) : (7'h47));
            end
          else
            begin
              reg1200 = $signed((reg1134[(3'h5):(1'h1)] >> $signed(($unsigned(reg1071) ?
                  reg1151[(4'h9):(3'h6)] : (!reg1187)))));
              reg1201 = ((8'hbc) ?
                  $signed($signed(((reg1097 ? reg1153 : reg1089) ?
                      reg1150 : {(8'hbd)}))) : ($unsigned($signed(reg1087[(3'h4):(2'h3)])) ?
                      $signed($unsigned($signed(wire1063))) : {(~^$unsigned(reg1136)),
                          forvar1156[(3'h5):(2'h3)],
                          ($unsigned(reg1121) ?
                              (reg1133 ?
                                  reg1168 : reg1194) : $signed(wire1147))}));
              reg1202 = ((~&(wire1064[(3'h5):(3'h5)] ?
                  ($unsigned(reg1192) ~^ (wire1063 ?
                      reg1100 : reg1117)) : ((&reg1186) ?
                      $signed(reg1140) : $signed((7'h40))))) && forvar1166);
              reg1203 = {($signed({reg1121, reg1188[(1'h0):(1'h0)]}) ?
                      reg1129 : $unsigned(reg1197)),
                  $signed((wire1147[(1'h0):(1'h0)] ?
                      $signed((forvar1169 | reg1181)) : {$unsigned(reg1155)})),
                  (8'hba)};
            end
          if ((~reg1189))
            begin
              reg1204 <= $signed((^reg1078[(5'h11):(2'h3)]));
              reg1205 <= ($unsigned(reg1199[(3'h4):(3'h4)]) | reg1174);
            end
          else
            begin
              reg1206 = reg1154[(4'he):(2'h2)];
              reg1207 = {$signed((^~({reg1193} ?
                      (^reg1122) : (reg1176 >> (7'h4d)))))};
              reg1208 = (($unsigned(reg1075[(3'h5):(3'h5)]) || {{reg1175[(5'h13):(4'h8)],
                      (reg1152 ? reg1201 : (7'h4c))},
                  ($unsigned(forvar1169) ?
                      (~^reg1161) : reg1159[(4'ha):(2'h2)])}) ^~ reg1157);
              reg1209 <= ((reg1191 + reg1167) ?
                  {$unsigned((^reg1192)),
                      $signed({wire1065[(3'h6):(2'h3)]}),
                      (reg1122 ?
                          $signed(wire1065[(5'h12):(4'h8)]) : $signed(reg1151))} : reg1196[(2'h3):(1'h0)]);
            end
          reg1210 = ({$unsigned($unsigned(((7'h4b) ? reg1084 : reg1203))),
              reg1201} <= ((~(8'hb2)) ?
              (+$unsigned(reg1090)) : $signed((~&{(7'h4a), forvar1148}))));
          reg1211 <= $signed($unsigned($unsigned(((&reg1097) ?
              (~^reg1179) : $signed(reg1209)))));
          for (forvar1212 = (1'h0); (forvar1212 < (2'h2)); forvar1212 = (forvar1212 + (1'h1)))
            begin
              reg1213 = $signed(((($signed(reg1192) != $signed(reg1152)) == (~(!reg1157))) * (reg1182 | {(reg1129 ?
                      (8'hb4) : reg1153)})));
              reg1214 <= $unsigned($signed((7'h56)));
              reg1215 = ((!reg1179[(2'h2):(2'h2)]) <<< $unsigned(reg1125[(5'h11):(4'hf)]));
              reg1216 <= (((&$signed((reg1104 ?
                      reg1179 : reg1070))) ^ reg1071[(3'h6):(3'h4)]) ?
                  (reg1181[(4'hd):(4'ha)] & $signed($signed(reg1171))) : forvar1178);
            end
        end
      else
        begin
          reg1204 <= ((((wire1063[(3'h4):(2'h3)] ? reg1153 : reg1090) ?
              $signed((forvar1176 ?
                  reg1214 : reg1085)) : $unsigned(reg1164)) <<< ((reg1189[(2'h3):(2'h3)] ?
                  $signed(reg1100) : ((8'hb9) - wire1147)) ?
              reg1172[(4'hd):(1'h0)] : $signed($signed(reg1125)))) <<< $signed((~^{forvar1178,
              reg1208})));
          for (forvar1205 = (1'h0); (forvar1205 < (1'h1)); forvar1205 = (forvar1205 + (1'h1)))
            begin
              reg1206 = {(8'hb5), reg1184, reg1174};
              reg1209 <= reg1215[(1'h1):(1'h0)];
              reg1211 <= reg1183;
              reg1212 <= $unsigned(reg1161);
              reg1214 <= ($unsigned($unsigned(reg1215)) && ((reg1177 ~^ reg1172[(2'h3):(1'h1)]) <<< (|$unsigned($signed(forvar1205)))));
            end
          reg1215 = reg1211;
          for (forvar1216 = (1'h0); (forvar1216 < (3'h6)); forvar1216 = (forvar1216 + (1'h1)))
            begin
              reg1217 = ($unsigned((($signed(forvar1205) ?
                      (8'hb6) : (|(7'h4d))) ?
                  reg1120[(3'h5):(3'h5)] : reg1180)) - (-wire1065[(4'hf):(4'hf)]));
              reg1218 = ($signed($unsigned(($unsigned((8'h9d)) ^~ $unsigned((8'ha7))))) >>> (~^$signed((~&$unsigned(reg1194)))));
            end
          reg1219 = {reg1117[(5'h11):(4'hd)]};
          if ({$unsigned(forvar1166[(4'hb):(2'h3)])})
            begin
              reg1220 = ((^reg1185[(5'h13):(2'h3)]) ?
                  $unsigned((((reg1154 ? forvar1176 : reg1084) ?
                          $unsigned(reg1181) : $signed(reg1129)) ?
                      (reg1084 ?
                          reg1133[(1'h1):(1'h0)] : reg1168) : $signed(reg1157))) : reg1087);
              reg1221 <= reg1163[(1'h1):(1'h1)];
            end
          else
            begin
              reg1221 <= reg1220;
              reg1222 <= {(&($signed(reg1197[(1'h0):(1'h0)]) ?
                      ($unsigned(reg1089) * (reg1091 ?
                          wire1066 : reg1190)) : (~reg1202[(2'h3):(1'h0)]))),
                  ((~^wire1064) || (8'hb2)),
                  forvar1176};
              reg1223 <= (({reg1217, reg1087} ?
                  wire1147 : (reg1199[(1'h0):(1'h0)] >>> forvar1216)) ^ ($signed(((reg1159 ?
                  reg1187 : reg1105) ^~ reg1092)) - reg1208[(3'h5):(1'h0)]));
              reg1224 = reg1193;
              reg1225 <= (~&(8'hbe));
              reg1226 <= $signed(($unsigned((~reg1071)) ^ $unsigned({reg1134[(3'h7):(3'h7)],
                  (reg1126 ? wire1147 : reg1075)})));
              reg1227 = (~|$signed((((reg1152 != reg1091) == (^~reg1073)) ?
                  {reg1075[(3'h6):(1'h0)]} : $unsigned(((8'hb1) < (8'ha0))))));
            end
          reg1228 = reg1099;
        end
      reg1229 <= reg1220;
      reg1230 <= $unsigned($unsigned(($unsigned($signed(reg1183)) && ($unsigned(reg1184) ^ {reg1202}))));
      if ({reg1079,
          ((($signed(reg1174) ? $signed(reg1075) : (+reg1100)) ?
                  (((8'hb3) >> (7'h57)) ?
                      (^~reg1085) : reg1174[(1'h0):(1'h0)]) : {(reg1126 ?
                          reg1174 : forvar1178),
                      reg1099[(3'h6):(3'h6)]}) ?
              (reg1090[(5'h13):(5'h12)] || ((reg1189 ?
                  reg1225 : reg1206) >= $unsigned(reg1196))) : $unsigned({$unsigned((7'h43))}))})
        begin
          for (forvar1231 = (1'h0); (forvar1231 < (3'h6)); forvar1231 = (forvar1231 + (1'h1)))
            begin
              reg1232 = ((($signed($signed(reg1193)) - reg1079) != reg1089[(4'h8):(3'h5)]) ?
                  (($signed($unsigned(reg1217)) < (~^(^reg1228))) >= ($unsigned((reg1230 ?
                          reg1221 : wire1061)) ?
                      (~forvar1176[(3'h7):(1'h1)]) : {$signed(forvar1205)})) : ((((reg1152 ?
                          reg1200 : reg1223) <= {(8'h9e),
                          (7'h48)}) == ((reg1209 < reg1150) ?
                          $signed(reg1168) : (~&reg1097))) ?
                      $signed($unsigned($signed(reg1202))) : $signed({(reg1196 ?
                              reg1123 : (8'hb1)),
                          $unsigned((8'hb6)),
                          ((8'hbd) | (7'h4f))})));
              reg1233 = {(~{$unsigned(reg1120), reg1071[(4'ha):(4'ha)]}),
                  $unsigned((!(^$signed(forvar1166))))};
              reg1234 <= reg1155[(5'h19):(3'h6)];
              reg1235 = $signed(reg1089[(3'h5):(3'h5)]);
            end
          reg1236 <= $signed($signed($unsigned(((&reg1160) ?
              $unsigned(reg1138) : $unsigned(reg1161)))));
          reg1237 <= {$unsigned(($unsigned($signed(reg1158)) ?
                  $unsigned({reg1224,
                      reg1129,
                      reg1126}) : (reg1208[(3'h5):(2'h3)] ?
                      $unsigned(reg1138) : (reg1099 ? reg1121 : reg1227)))),
              reg1223};
          reg1238 = $unsigned($signed($signed($signed(reg1089[(3'h5):(1'h1)]))));
        end
      else
        begin
          reg1231 = reg1216;
          for (forvar1232 = (1'h0); (forvar1232 < (1'h1)); forvar1232 = (forvar1232 + (1'h1)))
            begin
              reg1233 = (7'h40);
              reg1234 <= ((8'haf) - {(~&(~((7'h4d) ? reg1111 : reg1081))),
                  $unsigned(forvar1205)});
              reg1235 = {(+{$signed((reg1220 ? reg1078 : (8'ha5))),
                      (wire1065[(1'h1):(1'h1)] != reg1075),
                      $unsigned(reg1085[(4'h8):(3'h6)])}),
                  reg1234[(3'h7):(3'h6)]};
              reg1238 = $signed($unsigned(($unsigned(reg1121[(2'h3):(1'h0)]) ?
                  (&reg1111[(2'h2):(1'h0)]) : reg1192)));
              reg1239 <= reg1179;
              reg1240 <= (~&$signed(($signed(((7'h44) && (7'h50))) ?
                  ($unsigned(reg1187) ?
                      (reg1236 <= reg1193) : reg1208[(3'h6):(3'h5)]) : ({(8'haa),
                          (7'h55),
                          reg1089} ?
                      (~(7'h4d)) : (~^reg1239)))));
            end
        end
    end
  assign wire1241 = ((^reg1079[(1'h1):(1'h1)]) ?
                        (reg1104 ?
                            $signed(reg1081[(1'h0):(1'h0)]) : reg1190) : {((~|$signed(reg1165)) >= (~&reg1226)),
                            $signed($signed($unsigned(wire1147))),
                            $signed({(reg1169 != reg1084)})});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module543
#(parameter param837 = ((((((8'ha3) ? (8'hb4) : (8'ha8)) <<< ((7'h4b) <= (8'ha8))) * (((8'hb3) & (8'hb3)) ? ((8'ha7) ? (8'ha7) : (7'h55)) : (~&(8'ha1)))) ? ((^((7'h52) != (8'hac))) ? (((8'hb1) ? (8'hb9) : (7'h45)) ? ((8'hb0) ? (7'h51) : (8'hb8)) : {(7'h52), (7'h57)}) : (!((8'h9d) ^~ (7'h40)))) : (~^(((7'h51) & (7'h4d)) ? {(8'h9d), (8'hac)} : ((7'h58) || (8'h9d))))) ^~ ((~&{((8'hbb) ? (8'hae) : (8'hb4))}) ? ((^~(^~(8'ha9))) ? (((7'h50) <<< (8'h9d)) ? {(8'haa)} : ((7'h45) >>> (7'h57))) : (7'h42)) : ({((7'h48) ? (7'h43) : (7'h4c))} ? (^{(8'hae), (8'haa), (7'h43)}) : (+(!(7'h52)))))))
(y, clk, wire547, wire546, wire545, wire544);
  output wire [(32'h12fe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire547;
  input wire [(4'h9):(1'h0)] wire546;
  input wire signed [(2'h2):(1'h0)] wire545;
  input wire [(3'h4):(1'h0)] wire544;
  wire signed [(4'h8):(1'h0)] wire836;
  wire signed [(3'h4):(1'h0)] wire835;
  wire [(2'h3):(1'h0)] wire816;
  wire signed [(5'h19):(1'h0)] wire815;
  wire [(5'h13):(1'h0)] wire814;
  wire [(5'h14):(1'h0)] wire813;
  wire signed [(5'h1f):(1'h0)] wire636;
  wire [(2'h2):(1'h0)] wire579;
  reg signed [(5'h14):(1'h0)] reg833 = (1'h0);
  reg signed [(4'he):(1'h0)] reg832 = (1'h0);
  reg [(5'h19):(1'h0)] reg831 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg830 = (1'h0);
  reg [(5'h17):(1'h0)] reg826 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg825 = (1'h0);
  reg [(4'ha):(1'h0)] reg821 = (1'h0);
  reg [(4'ha):(1'h0)] reg820 = (1'h0);
  reg [(4'hc):(1'h0)] reg819 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg818 = (1'h0);
  reg [(4'hf):(1'h0)] reg812 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg811 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg806 = (1'h0);
  reg [(5'h11):(1'h0)] reg802 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg801 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg797 = (1'h0);
  reg [(4'ha):(1'h0)] reg796 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg795 = (1'h0);
  reg [(5'h13):(1'h0)] reg792 = (1'h0);
  reg [(4'h8):(1'h0)] reg787 = (1'h0);
  reg [(5'h18):(1'h0)] reg782 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg779 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg777 = (1'h0);
  reg [(2'h2):(1'h0)] reg772 = (1'h0);
  reg [(4'hb):(1'h0)] reg769 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg768 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg767 = (1'h0);
  reg [(4'hf):(1'h0)] reg766 = (1'h0);
  reg [(5'h14):(1'h0)] reg763 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg756 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg755 = (1'h0);
  reg [(4'hb):(1'h0)] reg753 = (1'h0);
  reg [(5'h18):(1'h0)] reg752 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg750 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg748 = (1'h0);
  reg [(5'h15):(1'h0)] reg743 = (1'h0);
  reg [(5'h10):(1'h0)] reg742 = (1'h0);
  reg [(5'h12):(1'h0)] reg741 = (1'h0);
  reg [(4'hd):(1'h0)] reg736 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg734 = (1'h0);
  reg [(5'h16):(1'h0)] reg731 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg729 = (1'h0);
  reg [(4'ha):(1'h0)] reg728 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg727 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg726 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg722 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg720 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg719 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg716 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg711 = (1'h0);
  reg [(5'h10):(1'h0)] reg708 = (1'h0);
  reg [(5'h11):(1'h0)] reg706 = (1'h0);
  reg [(5'h15):(1'h0)] reg703 = (1'h0);
  reg [(4'hc):(1'h0)] reg702 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg701 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg699 = (1'h0);
  reg [(2'h3):(1'h0)] reg697 = (1'h0);
  reg [(2'h2):(1'h0)] reg696 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg695 = (1'h0);
  reg [(4'h9):(1'h0)] reg694 = (1'h0);
  reg [(5'h18):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg692 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg690 = (1'h0);
  reg [(4'ha):(1'h0)] reg688 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg687 = (1'h0);
  reg [(5'h16):(1'h0)] reg686 = (1'h0);
  reg [(2'h2):(1'h0)] reg683 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg682 = (1'h0);
  reg [(5'h10):(1'h0)] reg679 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg675 = (1'h0);
  reg [(5'h13):(1'h0)] reg672 = (1'h0);
  reg [(4'he):(1'h0)] reg671 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg666 = (1'h0);
  reg [(5'h16):(1'h0)] reg665 = (1'h0);
  reg [(4'ha):(1'h0)] reg661 = (1'h0);
  reg [(4'hb):(1'h0)] reg657 = (1'h0);
  reg [(5'h12):(1'h0)] reg656 = (1'h0);
  reg [(5'h1b):(1'h0)] reg655 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg653 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg647 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg642 = (1'h0);
  reg [(2'h2):(1'h0)] reg639 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg635 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg626 = (1'h0);
  reg [(2'h2):(1'h0)] reg615 = (1'h0);
  reg [(5'h1d):(1'h0)] reg619 = (1'h0);
  reg [(5'h17):(1'h0)] reg618 = (1'h0);
  reg [(5'h14):(1'h0)] reg617 = (1'h0);
  reg [(4'h9):(1'h0)] reg613 = (1'h0);
  reg [(5'h11):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg611 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg606 = (1'h0);
  reg [(5'h1c):(1'h0)] reg605 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg604 = (1'h0);
  reg signed [(4'he):(1'h0)] reg601 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg598 = (1'h0);
  reg [(4'hf):(1'h0)] reg596 = (1'h0);
  reg [(5'h16):(1'h0)] reg595 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg594 = (1'h0);
  reg [(5'h15):(1'h0)] reg593 = (1'h0);
  reg [(5'h17):(1'h0)] reg590 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg589 = (1'h0);
  reg [(2'h3):(1'h0)] reg582 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg588 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg585 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg584 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg581 = (1'h0);
  reg [(4'hf):(1'h0)] reg578 = (1'h0);
  reg [(4'ha):(1'h0)] reg573 = (1'h0);
  reg [(5'h19):(1'h0)] reg572 = (1'h0);
  reg signed [(4'he):(1'h0)] reg566 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg565 = (1'h0);
  reg [(5'h1a):(1'h0)] reg562 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg834 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg829 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg828 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg827 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg824 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar823 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg822 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar817 = (1'h0);
  reg [(5'h1e):(1'h0)] reg810 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar809 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg808 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg807 = (1'h0);
  reg [(5'h18):(1'h0)] reg805 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg803 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg800 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg799 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg798 = (1'h0);
  reg [(4'hb):(1'h0)] forvar794 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg793 = (1'h0);
  reg [(4'he):(1'h0)] reg791 = (1'h0);
  reg [(4'he):(1'h0)] forvar790 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg789 = (1'h0);
  reg [(3'h6):(1'h0)] reg788 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg786 = (1'h0);
  reg [(4'hd):(1'h0)] forvar785 = (1'h0);
  reg [(5'h1c):(1'h0)] reg784 = (1'h0);
  reg [(5'h15):(1'h0)] reg783 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar781 = (1'h0);
  reg [(4'hd):(1'h0)] forvar778 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg776 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg775 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg774 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg773 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg771 = (1'h0);
  reg [(4'hf):(1'h0)] reg770 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg765 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg764 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar762 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg761 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg760 = (1'h0);
  reg [(4'hd):(1'h0)] reg759 = (1'h0);
  reg [(5'h17):(1'h0)] reg758 = (1'h0);
  reg [(4'hd):(1'h0)] forvar755 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg757 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar756 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar728 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg754 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar751 = (1'h0);
  reg [(2'h2):(1'h0)] reg749 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg747 = (1'h0);
  reg [(5'h1d):(1'h0)] reg746 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg745 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar744 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg740 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg739 = (1'h0);
  reg [(5'h14):(1'h0)] reg738 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg737 = (1'h0);
  reg [(5'h13):(1'h0)] reg735 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg733 = (1'h0);
  reg [(5'h19):(1'h0)] reg732 = (1'h0);
  reg [(3'h4):(1'h0)] reg730 = (1'h0);
  reg [(3'h5):(1'h0)] reg725 = (1'h0);
  reg [(5'h19):(1'h0)] reg724 = (1'h0);
  reg [(5'h18):(1'h0)] reg723 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg721 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg718 = (1'h0);
  reg [(3'h5):(1'h0)] reg717 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg714 = (1'h0);
  reg [(5'h14):(1'h0)] forvar713 = (1'h0);
  reg [(4'hc):(1'h0)] reg712 = (1'h0);
  reg [(5'h12):(1'h0)] reg710 = (1'h0);
  reg [(4'ha):(1'h0)] reg709 = (1'h0);
  reg [(5'h1f):(1'h0)] reg707 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg705 = (1'h0);
  reg signed [(4'he):(1'h0)] reg704 = (1'h0);
  reg [(4'hd):(1'h0)] reg700 = (1'h0);
  reg [(3'h4):(1'h0)] reg698 = (1'h0);
  reg [(4'hd):(1'h0)] reg691 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar689 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar685 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg684 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg681 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg680 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar667 = (1'h0);
  reg [(5'h1e):(1'h0)] reg678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg677 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg676 = (1'h0);
  reg [(5'h12):(1'h0)] reg674 = (1'h0);
  reg [(5'h11):(1'h0)] reg673 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg669 = (1'h0);
  reg [(4'h8):(1'h0)] forvar668 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg664 = (1'h0);
  reg [(5'h12):(1'h0)] forvar663 = (1'h0);
  reg [(4'h8):(1'h0)] reg662 = (1'h0);
  reg [(5'h1e):(1'h0)] reg660 = (1'h0);
  reg [(5'h19):(1'h0)] reg659 = (1'h0);
  reg [(5'h1f):(1'h0)] reg658 = (1'h0);
  reg [(5'h15):(1'h0)] reg654 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar652 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg650 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg649 = (1'h0);
  reg [(2'h3):(1'h0)] forvar648 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg648 = (1'h0);
  reg [(5'h17):(1'h0)] reg646 = (1'h0);
  reg [(5'h12):(1'h0)] reg645 = (1'h0);
  reg [(5'h18):(1'h0)] reg644 = (1'h0);
  reg [(5'h1f):(1'h0)] reg643 = (1'h0);
  reg [(5'h1a):(1'h0)] reg641 = (1'h0);
  reg [(4'h8):(1'h0)] forvar640 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar638 = (1'h0);
  reg [(5'h19):(1'h0)] reg637 = (1'h0);
  reg [(5'h19):(1'h0)] reg634 = (1'h0);
  reg [(2'h2):(1'h0)] reg633 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg631 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg630 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg629 = (1'h0);
  reg [(2'h2):(1'h0)] reg628 = (1'h0);
  reg [(4'hd):(1'h0)] reg627 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg625 = (1'h0);
  reg [(4'hb):(1'h0)] reg624 = (1'h0);
  reg [(5'h19):(1'h0)] reg623 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar622 = (1'h0);
  reg [(2'h3):(1'h0)] reg621 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg620 = (1'h0);
  reg [(5'h14):(1'h0)] forvar609 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar606 = (1'h0);
  reg [(4'h9):(1'h0)] reg616 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar615 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg614 = (1'h0);
  reg [(3'h7):(1'h0)] reg610 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg609 = (1'h0);
  reg [(5'h13):(1'h0)] reg607 = (1'h0);
  reg [(5'h16):(1'h0)] reg603 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg602 = (1'h0);
  reg [(5'h1c):(1'h0)] reg600 = (1'h0);
  reg [(5'h15):(1'h0)] forvar599 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg597 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg592 = (1'h0);
  reg [(5'h13):(1'h0)] reg591 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg587 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg586 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg583 = (1'h0);
  reg [(5'h13):(1'h0)] forvar582 = (1'h0);
  reg [(4'hf):(1'h0)] reg580 = (1'h0);
  reg [(5'h1e):(1'h0)] reg577 = (1'h0);
  reg [(5'h1b):(1'h0)] reg576 = (1'h0);
  reg [(4'ha):(1'h0)] reg575 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg574 = (1'h0);
  reg [(5'h19):(1'h0)] reg571 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg570 = (1'h0);
  reg [(5'h14):(1'h0)] reg569 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg568 = (1'h0);
  reg [(3'h6):(1'h0)] reg567 = (1'h0);
  reg [(5'h1b):(1'h0)] reg564 = (1'h0);
  reg [(4'hf):(1'h0)] reg563 = (1'h0);
  reg [(4'h9):(1'h0)] reg561 = (1'h0);
  reg [(4'h8):(1'h0)] reg560 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar559 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg558 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg557 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg556 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar555 = (1'h0);
  reg [(4'hc):(1'h0)] forvar554 = (1'h0);
  reg [(4'he):(1'h0)] reg553 = (1'h0);
  reg [(5'h15):(1'h0)] reg552 = (1'h0);
  reg signed [(4'he):(1'h0)] reg551 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg549 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar548 = (1'h0);
  assign y = {wire836,
                 wire835,
                 wire816,
                 wire815,
                 wire814,
                 wire813,
                 wire636,
                 wire579,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 reg826,
                 reg825,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 reg812,
                 reg811,
                 reg806,
                 reg802,
                 reg801,
                 reg797,
                 reg796,
                 reg795,
                 reg792,
                 reg787,
                 reg782,
                 reg780,
                 reg779,
                 reg777,
                 reg772,
                 reg769,
                 reg768,
                 reg767,
                 reg766,
                 reg763,
                 reg756,
                 reg755,
                 reg753,
                 reg752,
                 reg750,
                 reg748,
                 reg743,
                 reg742,
                 reg741,
                 reg736,
                 reg734,
                 reg731,
                 reg729,
                 reg728,
                 reg727,
                 reg726,
                 reg722,
                 reg720,
                 reg719,
                 reg716,
                 reg715,
                 reg711,
                 reg708,
                 reg706,
                 reg703,
                 reg702,
                 reg701,
                 reg699,
                 reg697,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg690,
                 reg688,
                 reg687,
                 reg686,
                 reg683,
                 reg682,
                 reg679,
                 reg668,
                 reg675,
                 reg672,
                 reg671,
                 reg670,
                 reg667,
                 reg666,
                 reg665,
                 reg661,
                 reg657,
                 reg656,
                 reg655,
                 reg653,
                 reg647,
                 reg642,
                 reg639,
                 reg635,
                 reg632,
                 reg626,
                 reg615,
                 reg619,
                 reg618,
                 reg617,
                 reg613,
                 reg612,
                 reg611,
                 reg608,
                 reg606,
                 reg605,
                 reg604,
                 reg601,
                 reg598,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg590,
                 reg589,
                 reg582,
                 reg588,
                 reg585,
                 reg584,
                 reg581,
                 reg578,
                 reg573,
                 reg572,
                 reg566,
                 reg565,
                 reg562,
                 reg834,
                 reg829,
                 reg828,
                 reg827,
                 reg824,
                 forvar823,
                 reg822,
                 forvar817,
                 reg810,
                 forvar809,
                 reg808,
                 reg807,
                 reg805,
                 reg804,
                 reg803,
                 reg800,
                 reg799,
                 reg798,
                 forvar794,
                 reg793,
                 reg791,
                 forvar790,
                 reg789,
                 reg788,
                 reg786,
                 forvar785,
                 reg784,
                 reg783,
                 forvar781,
                 forvar778,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 reg771,
                 reg770,
                 reg765,
                 reg764,
                 forvar762,
                 reg761,
                 reg760,
                 reg759,
                 reg758,
                 forvar755,
                 reg757,
                 forvar756,
                 forvar728,
                 reg754,
                 forvar751,
                 reg749,
                 reg747,
                 reg746,
                 reg745,
                 forvar744,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 reg735,
                 reg733,
                 reg732,
                 reg730,
                 reg725,
                 reg724,
                 reg723,
                 reg721,
                 reg718,
                 reg717,
                 reg714,
                 forvar713,
                 reg712,
                 reg710,
                 reg709,
                 reg707,
                 reg705,
                 reg704,
                 reg700,
                 reg698,
                 reg691,
                 forvar689,
                 forvar685,
                 reg684,
                 reg681,
                 reg680,
                 forvar667,
                 reg678,
                 reg677,
                 reg676,
                 reg674,
                 reg673,
                 reg669,
                 forvar668,
                 reg664,
                 forvar663,
                 reg662,
                 reg660,
                 reg659,
                 reg658,
                 reg654,
                 forvar652,
                 reg651,
                 reg650,
                 reg649,
                 forvar648,
                 reg648,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 reg641,
                 forvar640,
                 forvar638,
                 reg637,
                 reg634,
                 reg633,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg625,
                 reg624,
                 reg623,
                 forvar622,
                 reg621,
                 reg620,
                 forvar609,
                 forvar606,
                 reg616,
                 forvar615,
                 reg614,
                 reg610,
                 reg609,
                 reg607,
                 reg603,
                 reg602,
                 reg600,
                 forvar599,
                 reg597,
                 reg592,
                 reg591,
                 reg587,
                 reg586,
                 reg583,
                 forvar582,
                 reg580,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg564,
                 reg563,
                 reg561,
                 reg560,
                 forvar559,
                 reg558,
                 reg557,
                 reg556,
                 forvar555,
                 forvar554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 forvar548,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar548 = (1'h0); (forvar548 < (3'h6)); forvar548 = (forvar548 + (1'h1)))
        begin
          reg549 = $signed($unsigned($unsigned($unsigned(((7'h41) * (8'hb7))))));
          reg550 = (~|((wire546[(3'h6):(3'h5)] ?
              {wire545,
                  $unsigned(reg549)} : wire544[(1'h0):(1'h0)]) && ($unsigned((wire547 ^ reg549)) ?
              {{forvar548},
                  (wire546 ? reg549 : (7'h58)),
                  {wire545, (8'ha2), forvar548}} : wire545[(1'h1):(1'h1)])));
          reg551 = $unsigned(((($unsigned(reg549) | (|wire545)) - (~|(+wire544))) || (~$signed((~|wire547)))));
        end
      reg552 = $signed($signed(wire546[(1'h0):(1'h0)]));
      reg553 = (+$signed((+reg551[(4'hd):(3'h5)])));
      for (forvar554 = (1'h0); (forvar554 < (2'h3)); forvar554 = (forvar554 + (1'h1)))
        begin
          for (forvar555 = (1'h0); (forvar555 < (1'h0)); forvar555 = (forvar555 + (1'h1)))
            begin
              reg556 = reg553;
              reg557 = (-((~((forvar554 + reg550) ?
                      $unsigned((7'h54)) : (reg553 ? wire546 : (7'h57)))) ?
                  reg553 : reg549[(4'he):(4'ha)]));
              reg558 = (((!(+forvar554)) ?
                  (8'hb4) : reg551[(1'h0):(1'h0)]) * wire544);
            end
          for (forvar559 = (1'h0); (forvar559 < (3'h6)); forvar559 = (forvar559 + (1'h1)))
            begin
              reg560 = (^~$signed(reg551[(1'h0):(1'h0)]));
              reg561 = (|{(wire545 ?
                      {(reg560 ? wire546 : reg553)} : $unsigned({forvar559,
                          reg557,
                          (8'ha4)}))});
              reg562 <= ((reg553 ?
                      $unsigned(forvar555[(3'h4):(2'h3)]) : $signed((+reg552[(4'he):(2'h3)]))) ?
                  $unsigned((^~(~^(forvar559 || reg560)))) : (|({(8'ha5),
                      (7'h40),
                      (reg560 ?
                          (7'h54) : reg561)} & $signed(((8'haa) >> wire547)))));
              reg563 = $signed(wire547);
              reg564 = $unsigned(((~|((forvar559 ?
                  reg561 : wire547) + $unsigned(reg557))) > forvar548[(1'h1):(1'h1)]));
              reg565 <= reg563;
              reg566 <= reg561;
            end
          if (reg556[(3'h5):(3'h4)])
            begin
              reg567 = $unsigned((8'haf));
              reg568 = (7'h4a);
              reg569 = wire546;
              reg570 = (~|(((reg561[(1'h0):(1'h0)] ?
                      ((7'h4f) || wire547) : (|reg558)) && ((!(8'hb1)) ?
                      {reg564, (8'hae), reg566} : (reg553 <= reg568))) ?
                  ($unsigned((~^reg557)) ?
                      reg558 : (|((7'h50) & reg562))) : $signed((&(+(8'hb6))))));
              reg571 = wire545;
            end
          else
            begin
              reg572 <= (reg552 >> (($unsigned(forvar559) ?
                  reg560 : $signed(reg564)) > wire545));
              reg573 <= $signed($signed(forvar548[(5'h12):(4'hf)]));
              reg574 = forvar559[(3'h4):(1'h0)];
              reg575 = (~reg572[(4'h8):(3'h6)]);
              reg576 = $unsigned(($signed(((~|reg551) ?
                      (+forvar555) : {wire544, reg575, reg575})) ?
                  (7'h51) : reg561[(3'h7):(3'h7)]));
              reg577 = reg553[(3'h7):(3'h7)];
            end
        end
      reg578 <= reg572;
    end
  assign wire579 = $unsigned((wire544[(1'h0):(1'h0)] << $signed(wire545)));
  always
    @(posedge clk) begin
      if ((((reg562 << reg566[(3'h4):(2'h2)]) ?
              wire547[(4'ha):(3'h7)] : ($signed(reg565[(1'h0):(1'h0)]) ?
                  $signed(reg573[(1'h1):(1'h1)]) : ($signed((7'h57)) ?
                      wire544 : (+reg573)))) ?
          reg578 : (7'h4a)))
        begin
          reg580 = $unsigned(({(!(wire544 << reg573))} ~^ $unsigned($unsigned(wire546[(3'h5):(1'h0)]))));
          reg581 <= $unsigned(((~reg573[(4'ha):(4'ha)]) && ((7'h52) ?
              ((reg573 ? wire547 : reg565) ?
                  ((8'hbb) ?
                      reg572 : wire544) : reg566[(3'h5):(3'h4)]) : reg573)));
          for (forvar582 = (1'h0); (forvar582 < (3'h5)); forvar582 = (forvar582 + (1'h1)))
            begin
              reg583 = $signed($signed(reg580[(4'hd):(4'hc)]));
              reg584 <= (reg565 ?
                  wire547 : ($unsigned($signed(reg573[(1'h1):(1'h1)])) ?
                      ({(!forvar582), (reg581 ^~ reg581)} ?
                          ($signed(reg562) >= wire544[(2'h2):(1'h0)]) : reg566[(4'he):(4'h9)]) : {reg581[(4'h8):(3'h7)],
                          ((reg573 && wire546) ?
                              wire545[(1'h1):(1'h0)] : (~|reg573)),
                          $signed({reg572, wire547, (7'h44)})}));
            end
          reg585 <= ((wire547 ~^ (wire544 <<< wire544[(3'h4):(1'h1)])) || reg578[(1'h1):(1'h0)]);
          reg586 = ($unsigned(reg565) ?
              $signed(wire547[(1'h0):(1'h0)]) : $unsigned(($signed((reg578 ?
                      (8'ha9) : reg580)) ?
                  ($signed(reg562) ?
                      {(8'hbd),
                          reg583} : (reg584 & forvar582)) : {$unsigned((7'h49)),
                      ((7'h48) == reg565),
                      $signed((8'haa))})));
          reg587 = ((((reg583 ?
                  (~^reg583) : $unsigned(wire579)) << (wire547 << (forvar582 ?
                  forvar582 : forvar582))) >= wire579) ?
              ((~$signed(reg580[(2'h2):(2'h2)])) ?
                  ($unsigned($unsigned(wire545)) | wire547) : {((^forvar582) ?
                          $unsigned(reg562) : $signed(wire545)),
                      {(reg566 ? reg580 : reg585),
                          reg581,
                          $signed(wire547)}}) : $signed($signed(reg565[(1'h0):(1'h0)])));
          reg588 <= {((-(reg580 ?
                  reg581[(1'h1):(1'h1)] : $signed((7'h57)))) | $signed($signed(wire544))),
              $unsigned((|reg573)),
              (~({(^reg566)} ?
                  (reg583[(2'h3):(2'h3)] >= {reg580,
                      (8'hb2),
                      reg565}) : (((8'hb0) - reg581) - (reg562 ?
                      reg572 : reg586))))};
        end
      else
        begin
          if (reg566)
            begin
              reg580 = (({reg585[(1'h0):(1'h0)],
                          ((-reg562) != ((8'h9e) || (8'had))),
                          ((8'hab) ?
                              (wire545 ? wire544 : (7'h43)) : (reg565 ?
                                  reg572 : (7'h56)))} ?
                      ((~{reg578, (7'h53), reg581}) ?
                          $unsigned((wire546 ?
                              reg578 : wire544)) : ($unsigned((8'ha2)) ?
                              reg562[(5'h12):(4'hf)] : $unsigned(wire579))) : ($unsigned(wire579[(1'h0):(1'h0)]) ^ $signed(reg584))) ?
                  (-(|wire545[(1'h1):(1'h1)])) : ((^~$signed((^~reg562))) ?
                      (reg580 + ((^~forvar582) >>> wire545)) : (~^{$signed((8'hbd))})));
              reg581 <= wire545[(2'h2):(2'h2)];
              reg582 <= wire544;
              reg583 = $signed((&reg586[(5'h11):(4'hb)]));
              reg586 = {$signed(({reg562[(1'h0):(1'h0)],
                          {(8'ha2), (8'hb1), (8'ha3)}} ?
                      $signed(reg584[(2'h3):(1'h1)]) : ((reg572 ?
                              reg562 : reg580) ?
                          $unsigned(reg578) : (reg566 <<< wire545)))),
                  reg585,
                  (reg573 ?
                      ($unsigned((reg584 > reg586)) >= reg565[(2'h3):(2'h3)]) : forvar582[(4'h9):(2'h2)])};
              reg588 <= reg585[(1'h0):(1'h0)];
            end
          else
            begin
              reg581 <= reg580[(4'h8):(3'h7)];
              reg582 <= reg578[(4'ha):(1'h1)];
            end
        end
      if ({wire547,
          (~&reg562[(5'h12):(4'hb)]),
          $signed($signed(($unsigned(forvar582) ?
              (reg580 ? reg578 : reg562) : (!reg588))))})
        begin
          if ($unsigned(($signed($signed($signed((8'hbd)))) ?
              $signed($unsigned({reg586})) : reg588)))
            begin
              reg589 <= {((!(wire579 || $unsigned(reg562))) ?
                      {$signed($signed(reg588))} : (((reg566 >>> reg583) ?
                          reg565[(2'h2):(2'h2)] : (!reg587)) <<< ((-forvar582) >> wire544))),
                  {$unsigned($unsigned({(7'h50), reg582, reg562})),
                      ({(reg587 <= reg584),
                          $signed(reg585),
                          $unsigned(reg587)} || $signed($signed(reg578)))}};
              reg590 <= {$unsigned((|($unsigned(reg580) ~^ $signed(reg572)))),
                  wire579,
                  {{(+{reg584, reg566, wire547}), (!$unsigned(reg566))},
                      $signed($signed((7'h47))),
                      (((wire579 << reg583) ?
                          (8'hb6) : (-reg573)) < $signed((wire546 * reg586)))}};
              reg591 = $signed((~^{((reg581 ? reg581 : reg589) ?
                      wire545[(2'h2):(1'h0)] : (wire545 <<< (8'h9d))),
                  $signed((-reg562)),
                  $unsigned((wire544 ? (8'hb8) : reg572))}));
              reg592 = $signed((~reg589[(4'h8):(4'h8)]));
              reg593 <= {(~^wire546)};
            end
          else
            begin
              reg591 = {wire547,
                  $unsigned((~^(~^(reg592 ? (8'hbc) : (7'h4f))))),
                  $signed(reg593[(3'h5):(1'h0)])};
              reg593 <= ({wire544} ?
                  $unsigned(((^~{reg583, reg583}) ?
                      reg592 : $unsigned($unsigned(reg593)))) : reg585);
              reg594 <= ((~^$signed(((8'h9e) != reg587))) <<< ($unsigned(((reg583 ?
                  reg585 : forvar582) >= reg588)) + reg587));
              reg595 <= (-wire547);
              reg596 <= (-reg588);
            end
        end
      else
        begin
          if ((($signed(($signed(reg596) + $unsigned(reg582))) != (((!wire545) ^ ((8'h9e) ?
              reg578 : (7'h4f))) != ($unsigned(reg578) <<< reg566[(3'h7):(3'h6)]))) || (~&($signed((|reg573)) ?
              ((&wire544) << {(8'hb4), reg583, reg591}) : reg591))))
            begin
              reg589 <= $signed(wire547);
              reg590 <= ({reg562} <= reg591[(3'h7):(2'h2)]);
            end
          else
            begin
              reg589 <= $signed($signed($unsigned(reg592)));
              reg590 <= (~|$signed(reg593[(4'hc):(3'h4)]));
              reg593 <= forvar582;
              reg597 = (+reg573);
              reg598 <= reg597[(4'ha):(1'h1)];
            end
          for (forvar599 = (1'h0); (forvar599 < (1'h0)); forvar599 = (forvar599 + (1'h1)))
            begin
              reg600 = ($unsigned((~|(reg597 * (wire579 ? reg584 : (7'h48))))) ?
                  ($unsigned($signed((reg566 ?
                      reg572 : reg590))) < reg597[(2'h3):(1'h0)]) : ((+{$signed(reg595),
                          reg591[(4'hc):(3'h4)]}) ?
                      reg562[(5'h13):(2'h3)] : ((^~$unsigned(reg572)) ?
                          $unsigned($unsigned(reg583)) : $unsigned(reg597[(4'h8):(1'h1)]))));
              reg601 <= $unsigned((+(8'ha0)));
              reg602 = (^$signed(($signed((reg593 << reg584)) ?
                  $unsigned((8'ha3)) : reg584[(2'h2):(1'h1)])));
              reg603 = $signed(((-(~|(reg580 ? (8'hb5) : reg584))) ?
                  $signed(((&reg592) | (-(8'hae)))) : (reg590[(5'h15):(3'h5)] >= {(reg600 - wire544),
                      reg562[(2'h2):(1'h1)]})));
              reg604 <= (reg591[(5'h11):(4'hd)] ?
                  (|($unsigned($unsigned(wire579)) ?
                      ({reg591, reg593} ? (reg588 ^ reg602) : reg565) : {reg586,
                          reg596})) : {(!((reg578 ?
                          (8'ha9) : reg596) ^~ reg573[(3'h5):(1'h0)]))});
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned((^$signed($unsigned((wire579 >> reg601))))))
        begin
          if ($signed($signed((8'h9c))))
            begin
              reg605 <= $unsigned(($unsigned($unsigned((~&(7'h4a)))) ?
                  $unsigned((^(reg604 ?
                      (8'hbe) : reg598))) : {($signed(reg565) <<< (reg598 ?
                          (8'hab) : (8'ha6)))}));
              reg606 <= (reg578[(3'h4):(2'h2)] ?
                  (&(reg605 ? {(!wire579)} : $signed((7'h48)))) : wire547);
            end
          else
            begin
              reg607 = ($signed($signed(((reg604 >> reg593) ?
                  reg565[(1'h0):(1'h0)] : $unsigned(reg578)))) & ($unsigned((~&reg581[(3'h5):(3'h4)])) <<< {(~|(reg566 < reg584))}));
              reg608 <= (~&$signed(reg582));
              reg609 = (&$signed((($unsigned(reg594) || $signed(reg581)) && wire547)));
              reg610 = (reg606 <<< reg598);
              reg611 <= (reg596 || {{{$signed(reg608), reg601}},
                  (reg573 ?
                      $signed((reg595 ?
                          (8'ha5) : reg606)) : $unsigned(((8'hb0) ?
                          reg598 : (8'hb3))))});
              reg612 <= ($unsigned($signed(reg595[(4'hd):(4'hb)])) ?
                  (reg605 ?
                      ($unsigned($signed(reg609)) ^~ reg594[(4'hc):(4'h8)]) : $unsigned($unsigned(((8'h9e) || reg608)))) : wire546);
              reg613 <= (((reg593[(5'h10):(2'h2)] >> reg601[(1'h1):(1'h0)]) ~^ (~reg598[(3'h4):(2'h3)])) - (-reg609));
            end
          reg614 = wire579[(2'h2):(1'h1)];
          for (forvar615 = (1'h0); (forvar615 < (1'h1)); forvar615 = (forvar615 + (1'h1)))
            begin
              reg616 = ($unsigned(reg566) - wire546);
              reg617 <= ($signed(reg566) > {reg596,
                  (reg606 >>> reg606[(4'h9):(2'h2)]),
                  (reg578[(3'h4):(3'h4)] ^ reg582[(2'h3):(1'h0)])});
            end
          reg618 <= reg604;
          reg619 <= reg572[(5'h18):(2'h3)];
        end
      else
        begin
          reg605 <= (|reg595);
          for (forvar606 = (1'h0); (forvar606 < (3'h4)); forvar606 = (forvar606 + (1'h1)))
            begin
              reg608 <= reg618;
            end
          for (forvar609 = (1'h0); (forvar609 < (3'h5)); forvar609 = (forvar609 + (1'h1)))
            begin
              reg611 <= {reg594[(3'h6):(2'h3)],
                  (reg595[(5'h14):(3'h7)] ?
                      (~&(&(reg593 ? (7'h52) : reg581))) : (7'h51)),
                  (-$unsigned(wire547[(4'hd):(4'h9)]))};
              reg614 = {($signed((reg585[(2'h3):(2'h3)] != reg613[(4'h8):(3'h7)])) <= reg566[(3'h4):(2'h2)]),
                  (+$unsigned({reg612, reg581[(1'h0):(1'h0)], reg565})),
                  (^reg611)};
              reg615 <= $signed($signed(((reg616[(4'h8):(1'h1)] <= reg588) ?
                  ($signed(reg613) >>> (reg562 ?
                      reg601 : (8'ha7))) : $unsigned(wire545))));
              reg616 = wire547[(4'he):(4'hd)];
              reg617 <= (7'h4f);
              reg620 = ((((forvar606[(1'h0):(1'h0)] ?
                              reg584[(2'h2):(1'h1)] : {reg606}) ?
                          reg565 : (((8'h9d) ? reg604 : reg601) ?
                              (~|reg606) : (wire546 ? reg565 : reg617))) ?
                      {$unsigned((reg608 >>> reg590)),
                          (&(reg578 <<< reg612))} : ($signed((reg572 <<< reg562)) ?
                          reg612[(4'hf):(3'h6)] : ((7'h53) >> $unsigned(reg598)))) ?
                  $unsigned(reg584[(2'h3):(2'h3)]) : ((reg615[(1'h0):(1'h0)] + $unsigned($signed(forvar609))) ^ reg573[(2'h2):(2'h2)]));
            end
          reg621 = (!$unsigned($signed((^~reg578[(2'h3):(2'h2)]))));
          for (forvar622 = (1'h0); (forvar622 < (2'h2)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 = (^~reg578);
              reg624 = {forvar622[(3'h6):(3'h6)], (~&reg578)};
              reg625 = reg619;
              reg626 <= $signed(reg601[(1'h0):(1'h0)]);
              reg627 = reg615[(2'h2):(2'h2)];
              reg628 = (&reg615[(2'h2):(1'h0)]);
              reg629 = $signed($signed(($signed((-wire547)) | (^~reg623))));
            end
          if ({(reg612[(4'ha):(2'h2)] ?
                  {(reg616[(3'h6):(2'h3)] ?
                          $unsigned(wire545) : $signed(reg593))} : reg601),
              ((+$signed($signed(forvar615))) ?
                  (~($signed(reg572) ?
                      reg566 : reg566[(4'hd):(3'h7)])) : $unsigned(reg606[(5'h11):(1'h1)])),
              reg584[(1'h0):(1'h0)]})
            begin
              reg630 = ($unsigned(($unsigned($unsigned(wire545)) - reg616)) << ((($signed(reg608) - ((7'h41) ?
                          reg582 : reg588)) ?
                      $unsigned((wire547 ? forvar615 : wire579)) : ((reg598 ?
                          reg584 : (8'hb9)) > reg617)) ?
                  forvar606 : reg614));
              reg631 = $signed((((reg610 ?
                      $unsigned(reg629) : $unsigned(reg606)) < $unsigned((reg630 ^~ reg629))) ?
                  {reg594[(4'h8):(1'h1)],
                      (^~(wire546 ? reg585 : reg572)),
                      ($unsigned(reg620) << (!reg627))} : (8'ha6)));
              reg632 <= reg625;
              reg633 = (!$signed((reg584 == reg578[(4'hb):(1'h0)])));
              reg634 = {wire544[(2'h2):(1'h1)]};
              reg635 <= $unsigned((reg581[(3'h4):(1'h0)] * forvar615));
            end
          else
            begin
              reg632 <= (reg632[(1'h1):(1'h0)] ?
                  reg615 : {reg582[(1'h0):(1'h0)],
                      (+(wire546 == reg628[(2'h2):(1'h1)])),
                      (($unsigned(reg601) && $signed((8'h9f))) != ($signed(reg605) * $unsigned(reg615)))});
              reg633 = reg596[(3'h6):(3'h4)];
            end
        end
    end
  assign wire636 = (reg598[(4'hb):(3'h5)] > (&(reg635 ?
                       reg604 : ((reg595 ?
                           reg608 : reg632) ^ $signed((7'h54))))));
  always
    @(posedge clk) begin
      reg637 = (8'hb1);
      for (forvar638 = (1'h0); (forvar638 < (1'h1)); forvar638 = (forvar638 + (1'h1)))
        begin
          reg639 <= (reg612[(3'h6):(1'h0)] <= $signed((7'h54)));
          for (forvar640 = (1'h0); (forvar640 < (3'h5)); forvar640 = (forvar640 + (1'h1)))
            begin
              reg641 = $signed(reg613);
            end
          reg642 <= ($signed(wire546) ?
              ($signed(wire545) & {$unsigned((reg604 ^~ reg605)),
                  (^wire579)}) : $signed(({((8'hb4) ~^ wire579),
                  $signed((7'h44)),
                  {reg639}} < reg566)));
          reg643 = $unsigned((~^reg572[(5'h13):(4'hf)]));
        end
      if ($signed(($unsigned($unsigned(reg604)) ?
          (((-reg595) ?
              ((8'ha2) < (7'h46)) : reg593[(2'h2):(1'h1)]) >= (forvar638 ?
              (reg606 >>> (7'h42)) : (+reg578))) : {$unsigned($signed(reg606))})))
        begin
          if ($signed($unsigned($unsigned(($unsigned(reg641) ?
              (|reg604) : (~|reg566))))))
            begin
              reg644 = (~reg590);
              reg645 = (8'hb3);
              reg646 = ({(reg562[(1'h0):(1'h0)] > (8'ha8)),
                      (($signed(reg566) ~^ $unsigned(reg642)) | reg595),
                      (^$unsigned((-(8'haf))))} ?
                  (reg598 <<< $signed({{wire544},
                      $signed(reg626),
                      $signed(reg598)})) : $unsigned((((&reg593) ?
                          $unsigned(reg588) : $signed(reg604)) ?
                      ($signed(reg584) ?
                          (reg593 ?
                              (8'ha3) : wire579) : (reg566 ^~ reg608)) : (&(reg590 ?
                          reg643 : reg619)))));
            end
          else
            begin
              reg647 <= wire545[(2'h2):(1'h1)];
              reg648 = (&$signed((~|(&$unsigned(wire636)))));
            end
        end
      else
        begin
          reg647 <= (^~$unsigned(reg632[(2'h2):(1'h0)]));
          for (forvar648 = (1'h0); (forvar648 < (1'h1)); forvar648 = (forvar648 + (1'h1)))
            begin
              reg649 = $unsigned(($unsigned($unsigned((reg618 * reg595))) << $signed(reg578[(2'h3):(2'h2)])));
            end
          reg650 = ($unsigned(reg626) ? $signed(reg613) : reg562);
        end
      reg651 = (reg593[(5'h13):(4'hd)] ?
          (reg619 ?
              forvar640 : $signed($unsigned((^reg643)))) : $signed({(~|(reg566 ?
                  reg632 : reg585))}));
      for (forvar652 = (1'h0); (forvar652 < (3'h5)); forvar652 = (forvar652 + (1'h1)))
        begin
          reg653 <= $unsigned($signed((reg626[(4'hb):(4'h8)] ?
              ((reg632 ? reg595 : reg642) < reg646[(5'h10):(4'h9)]) : reg615)));
          if ({$signed(reg585[(3'h4):(1'h1)]),
              reg632[(3'h6):(2'h2)],
              $signed((!$unsigned((^~(8'h9c)))))})
            begin
              reg654 = reg595;
              reg655 <= reg642[(3'h7):(1'h1)];
              reg656 <= {(~$signed(((-reg573) ~^ wire545[(1'h0):(1'h0)])))};
            end
          else
            begin
              reg655 <= $unsigned($unsigned(reg643[(4'ha):(3'h7)]));
            end
          if ((reg585 ? $signed($unsigned(reg649)) : reg651[(2'h3):(2'h2)]))
            begin
              reg657 <= $unsigned((reg604 ?
                  reg584[(1'h1):(1'h1)] : $unsigned(($unsigned(reg581) ?
                      reg651 : (reg584 ? reg598 : reg611)))));
              reg658 = reg618[(4'ha):(4'h9)];
              reg659 = ((^$signed($signed($signed(reg581)))) ?
                  reg649[(5'h16):(3'h6)] : ((wire547 * $signed($signed(wire547))) >> (reg649[(4'h9):(1'h0)] ?
                      $signed((reg645 << reg619)) : (reg595[(4'hf):(2'h3)] ?
                          $unsigned(reg650) : $unsigned(reg608)))));
              reg660 = (((-reg655) >= {reg635[(3'h6):(3'h6)],
                  $signed(reg653[(1'h1):(1'h0)])}) >>> ($signed(reg641[(5'h14):(3'h6)]) - $unsigned(({reg585} ?
                  (forvar652 <<< (8'ha1)) : (reg613 ? reg646 : reg562)))));
            end
          else
            begin
              reg657 <= (~(8'hab));
              reg661 <= {wire636, reg581};
              reg662 = reg590[(4'hc):(2'h3)];
            end
          for (forvar663 = (1'h0); (forvar663 < (3'h6)); forvar663 = (forvar663 + (1'h1)))
            begin
              reg664 = ({(~|forvar648),
                      $signed(({wire545, (8'hb8), (8'hbf)} ?
                          (reg654 ? reg590 : reg637) : (!wire544))),
                      $unsigned((&{wire547, reg619, reg651}))} ?
                  (($signed($signed(reg615)) ?
                      {reg635[(2'h2):(2'h2)]} : (-$unsigned(reg653))) > (!(8'had))) : (~|(-reg584[(2'h3):(2'h3)])));
              reg665 <= reg657[(2'h3):(2'h2)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg666 <= $signed(reg655[(5'h11):(3'h4)]);
      if (reg653[(3'h4):(1'h0)])
        begin
          reg667 <= (wire545[(1'h1):(1'h0)] & $signed(reg589[(1'h1):(1'h0)]));
          for (forvar668 = (1'h0); (forvar668 < (1'h0)); forvar668 = (forvar668 + (1'h1)))
            begin
              reg669 = reg573[(4'ha):(4'h8)];
              reg670 <= reg566;
              reg671 <= (^~(($signed(reg669[(2'h2):(1'h1)]) + (8'hb7)) ?
                  ($unsigned((reg656 != reg647)) ?
                      (~&reg585) : wire636[(4'h9):(4'h8)]) : reg601[(4'hd):(3'h4)]));
              reg672 <= (^~$signed($signed(reg667[(5'h11):(4'h8)])));
              reg673 = {reg566[(4'ha):(1'h0)], reg593[(3'h6):(3'h5)], reg647};
              reg674 = (reg647[(2'h2):(2'h2)] ?
                  $unsigned($unsigned($unsigned(reg613[(3'h4):(2'h3)]))) : (reg667 != wire546));
            end
          reg675 <= $unsigned((~^($signed(wire636) ?
              (~^wire546[(1'h0):(1'h0)]) : {$unsigned((7'h4f)),
                  (!reg611),
                  reg653[(2'h3):(2'h2)]})));
          reg676 = ($unsigned(($unsigned($unsigned(reg611)) && (~^(8'ha1)))) ?
              ((&reg670) >> {((reg611 ?
                      reg665 : reg606) + $unsigned(reg615))}) : $unsigned((((reg635 ?
                      reg604 : wire579) ?
                  (reg595 >= reg608) : wire636[(5'h1d):(5'h13)]) == reg655)));
          reg677 = ((+$signed((((8'hae) ? reg593 : wire544) ?
                  (+wire579) : (reg578 ? reg585 : reg613)))) ?
              $unsigned((8'h9f)) : (^~{{reg594, $unsigned(wire546)},
                  (-(reg572 ? (8'h9c) : reg626)),
                  (~|(&reg615))}));
          reg678 = forvar668;
        end
      else
        begin
          for (forvar667 = (1'h0); (forvar667 < (3'h6)); forvar667 = (forvar667 + (1'h1)))
            begin
              reg668 <= ((reg661[(3'h7):(3'h4)] ?
                  ($signed($unsigned(reg594)) ?
                      reg584 : ({reg670,
                          reg572,
                          reg588} * (8'hba))) : reg653) * $signed((~&$unsigned((-reg595)))));
              reg669 = (-($signed(($unsigned(reg596) ?
                      reg585 : ((7'h49) << reg666))) ?
                  ((~|(reg606 ? reg671 : reg656)) - ({reg626, reg615, reg632} ?
                      (reg656 + reg605) : ((7'h4f) <= reg612))) : (~&((&reg675) == $unsigned(wire545)))));
              reg670 <= $unsigned(reg671[(2'h2):(1'h1)]);
              reg673 = reg653[(2'h3):(2'h2)];
              reg674 = (-reg596);
            end
          reg675 <= ($unsigned(reg604) >> (($unsigned({reg675, reg647}) ?
                  ((reg601 >>> reg612) ?
                      reg619[(3'h5):(2'h2)] : $unsigned(reg612)) : (~(~|(8'hb9)))) ?
              $signed(reg594[(4'h9):(2'h3)]) : $unsigned(($signed(reg665) << $signed(reg632)))));
          if (((((~(reg671 << reg606)) == $unsigned((reg670 ?
              reg626 : reg588))) ^~ reg573[(3'h4):(1'h0)]) < (+reg606[(4'hd):(4'hb)])))
            begin
              reg676 = (8'ha5);
              reg679 <= ((reg604[(4'hc):(4'h8)] ?
                  (!$signed(((8'hbc) < reg672))) : $signed({(~|reg582),
                      $signed(reg605),
                      reg588[(1'h1):(1'h0)]})) ^~ (~^reg670[(3'h4):(1'h0)]));
              reg680 = $unsigned(reg593[(5'h11):(1'h1)]);
              reg681 = (7'h52);
              reg682 <= reg581;
            end
          else
            begin
              reg679 <= (&reg626[(4'he):(3'h6)]);
            end
        end
      reg683 <= (^{$signed($signed(reg673))});
      reg684 = reg642;
      for (forvar685 = (1'h0); (forvar685 < (2'h2)); forvar685 = (forvar685 + (1'h1)))
        begin
          reg686 <= $unsigned({reg674, reg635[(2'h2):(1'h1)]});
          reg687 <= (&($unsigned((8'hb1)) ~^ $signed(reg656)));
          reg688 <= (&$signed(wire547[(2'h2):(1'h0)]));
          for (forvar689 = (1'h0); (forvar689 < (3'h6)); forvar689 = (forvar689 + (1'h1)))
            begin
              reg690 <= {({$signed(wire579[(1'h1):(1'h0)]),
                          ((reg565 ? reg639 : reg642) <<< $signed((8'hb3))),
                          $signed(reg655[(3'h7):(3'h7)])} ?
                      $unsigned((+reg605[(1'h0):(1'h0)])) : reg639[(1'h1):(1'h0)]),
                  (-reg688[(4'h9):(3'h5)])};
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg601[(3'h6):(3'h4)])
        begin
          reg691 = ({$signed(($unsigned(reg653) ?
                      (^(8'hb7)) : $unsigned(reg657)))} ?
              (~&reg612[(4'h8):(3'h7)]) : $unsigned(reg613));
          reg692 <= ((((-(wire545 ? (8'hba) : reg613)) ?
                  ($unsigned(reg606) * $unsigned(reg655)) : reg682[(5'h19):(2'h2)]) ?
              ((~reg672[(5'h10):(2'h2)]) <= ((^~(8'hb6)) ?
                  $unsigned(reg666) : (^reg690))) : ((reg605 >= (reg656 ?
                      wire545 : reg671)) ?
                  ($signed(reg666) << reg565) : reg626[(5'h13):(5'h10)])) | (^$signed(reg565)));
        end
      else
        begin
          if (($signed((reg653[(2'h3):(1'h1)] ?
                  ((reg690 ^~ reg683) ?
                      wire579 : $unsigned(wire544)) : reg601[(4'hc):(4'h8)])) ?
              reg618 : (-($signed(((7'h4b) ^ reg666)) ?
                  (reg690 ~^ reg672) : reg656))))
            begin
              reg692 <= $signed(reg584);
              reg693 <= (((-(((8'ha9) ?
                      reg619 : reg683) ^ (~&reg589))) | (reg593[(3'h6):(1'h0)] ?
                      $unsigned(reg672) : ((~|reg578) ~^ reg584[(2'h3):(2'h2)]))) ?
                  wire579[(1'h1):(1'h1)] : $unsigned($signed((-(reg692 >>> reg679)))));
              reg694 <= reg601[(4'hb):(3'h5)];
              reg695 <= ((8'hb1) ?
                  reg653 : (-(reg670[(3'h4):(1'h0)] >> $unsigned((reg612 < (8'hbe))))));
              reg696 <= reg593;
              reg697 <= $unsigned($signed(reg596));
              reg698 = wire545[(1'h0):(1'h0)];
            end
          else
            begin
              reg692 <= (&$signed(reg642));
              reg698 = (~$unsigned((wire545[(2'h2):(2'h2)] - reg670[(1'h0):(1'h0)])));
              reg699 <= (reg691[(3'h6):(1'h0)] ?
                  reg667 : ($unsigned($unsigned(reg670[(3'h4):(1'h1)])) ?
                      (((reg661 & reg690) ^~ (reg665 ? reg693 : reg608)) ?
                          ($signed((7'h51)) ?
                              (~&reg565) : reg601[(1'h0):(1'h0)]) : (-(reg668 ?
                              reg655 : reg604))) : (-$unsigned({(8'hab),
                          reg617}))));
              reg700 = $signed(reg573[(2'h3):(2'h3)]);
            end
          reg701 <= (~^(reg588 >>> {$unsigned(reg573),
              $unsigned(reg626[(5'h13):(4'ha)])}));
          if ((($signed(((reg671 != wire579) ?
                  (-(7'h58)) : reg699[(2'h3):(2'h2)])) || $signed(reg565[(2'h2):(1'h1)])) ?
              $signed($unsigned(reg604)) : $unsigned($unsigned(((reg679 ^ reg589) <<< (~&reg613))))))
            begin
              reg702 <= reg688;
              reg703 <= ($unsigned(($signed((reg695 & (7'h54))) ?
                  (^$signed(reg572)) : (7'h44))) ~^ ((reg672 ?
                  ((reg572 >> reg566) ?
                      $unsigned((8'ha2)) : (reg601 << reg617)) : ($signed(reg657) <= {reg695,
                      wire547,
                      reg608})) | (+($signed((8'hbf)) > (reg572 ?
                  (7'h47) : reg615)))));
            end
          else
            begin
              reg702 <= reg572;
              reg704 = $unsigned({((^~reg635[(2'h3):(2'h3)]) <= (!reg675)),
                  reg698,
                  (|($unsigned(reg668) <= reg598))});
              reg705 = ((~|$unsigned((~^(reg675 != reg700)))) ?
                  ({($signed(reg615) ? $unsigned((8'haa)) : $unsigned(reg593)),
                      $signed(((7'h4c) | reg588))} == reg593[(4'hc):(4'hc)]) : $unsigned((wire546 ?
                      reg675[(5'h10):(2'h3)] : reg596[(4'h8):(3'h4)])));
            end
          if ($unsigned($unsigned((|reg611))))
            begin
              reg706 <= (!(|wire545));
              reg707 = $signed($unsigned(({((8'hbf) == wire546), reg686} ?
                  $unsigned((reg584 == reg588)) : $unsigned($signed(reg565)))));
              reg708 <= ($signed({{{reg593, reg626},
                      reg691[(2'h3):(1'h1)],
                      $unsigned(reg612)},
                  $signed($signed(reg657))}) && reg706[(4'hc):(4'ha)]);
            end
          else
            begin
              reg707 = ((({$unsigned(reg584), $signed(reg657)} ?
                      reg679[(4'h9):(3'h7)] : (reg595[(2'h3):(1'h1)] ?
                          {(7'h54), reg701} : $signed((7'h41)))) ?
                  (reg604 <= ((reg707 ? reg656 : reg588) ^~ (reg688 ?
                      (7'h46) : reg562))) : ($unsigned(reg706) ?
                      ((reg601 & reg578) ~^ reg705[(2'h3):(1'h0)]) : (8'hb3))) != reg604);
              reg709 = {reg706[(2'h2):(2'h2)]};
              reg710 = $unsigned((~(-$signed((reg682 >> reg657)))));
              reg711 <= {(7'h49)};
              reg712 = ((^~reg617) == $unsigned((reg613 - reg682)));
            end
          for (forvar713 = (1'h0); (forvar713 < (2'h3)); forvar713 = (forvar713 + (1'h1)))
            begin
              reg714 = $unsigned({reg619,
                  ($signed($signed(reg653)) ^~ ((~|reg613) >= reg647[(1'h1):(1'h0)]))});
            end
          reg715 <= ((~&(^~reg706[(4'hd):(2'h2)])) < (8'hb5));
        end
      if ($signed(((reg657[(4'ha):(3'h4)] != reg667) | $signed(reg672[(4'h8):(3'h6)]))))
        begin
          if ($unsigned((^$signed(reg665[(5'h14):(4'ha)]))))
            begin
              reg716 <= $signed((-$signed((!$unsigned(reg615)))));
              reg717 = wire545[(1'h0):(1'h0)];
              reg718 = (8'h9d);
              reg719 <= {{$signed((^~reg692[(3'h5):(1'h1)])),
                      reg582,
                      reg612[(4'hb):(2'h3)]},
                  $unsigned({$signed($unsigned(reg687)),
                      reg701[(5'h10):(3'h4)],
                      (reg712 >> $unsigned(reg606))}),
                  ((reg572[(3'h5):(1'h0)] + ((reg688 ? (8'hba) : reg690) ?
                          reg715[(2'h3):(2'h2)] : reg703[(5'h10):(4'h9)])) ?
                      (reg595[(3'h5):(3'h4)] ?
                          $signed((reg667 ? (8'h9c) : (8'hb1))) : ({reg573,
                                  reg718} ?
                              reg691 : reg679)) : ($signed((reg565 ?
                          forvar713 : reg639)) & reg595))};
              reg720 <= reg635;
              reg721 = $signed((~($signed(reg670[(2'h2):(2'h2)]) ?
                  $unsigned((~&reg595)) : ((reg656 ?
                      reg716 : (8'hbc)) >>> (reg711 == reg686)))));
            end
          else
            begin
              reg717 = $unsigned({(|({reg668} ? reg675 : (~|(8'ha0)))),
                  {reg698}});
              reg719 <= {reg710};
              reg721 = reg710;
              reg722 <= {reg566[(4'h9):(3'h5)],
                  (reg712 ^~ reg604),
                  $unsigned((($unsigned((7'h41)) * reg683) >>> $unsigned({reg711})))};
              reg723 = $unsigned(((7'h4c) ~^ ($unsigned(((8'hbc) ?
                      reg613 : reg604)) ?
                  $signed(reg632) : reg712[(3'h7):(3'h4)])));
            end
          if ($signed($unsigned(reg581[(5'h10):(4'hd)])))
            begin
              reg724 = reg683[(2'h2):(1'h0)];
              reg725 = (reg682 >> $unsigned((8'hae)));
              reg726 <= ({$unsigned(reg667),
                      $signed($unsigned(reg601[(3'h6):(1'h1)])),
                      $signed(reg632[(1'h0):(1'h0)])} ?
                  (~^$unsigned((~&$signed(reg572)))) : ($signed((+$unsigned((8'haf)))) ?
                      (($unsigned(reg721) ?
                              (reg694 ? reg724 : reg721) : $signed(reg718)) ?
                          reg605[(5'h1c):(5'h13)] : (reg613[(2'h2):(2'h2)] ?
                              $signed(reg702) : (forvar713 > (8'ha7)))) : reg690[(5'h17):(2'h3)]));
              reg727 <= $unsigned($signed($unsigned((reg608[(1'h0):(1'h0)] ?
                  $unsigned(reg672) : (reg588 ? (8'hb9) : (8'ha1))))));
              reg728 <= (((reg721[(5'h15):(5'h10)] * $signed($signed(reg670))) ?
                  $unsigned($signed(reg719[(4'ha):(4'h9)])) : $signed((^~$unsigned(wire579)))) >> reg717[(1'h1):(1'h1)]);
              reg729 <= (-$unsigned($unsigned({wire544[(1'h1):(1'h1)],
                  (reg687 ? reg702 : reg690),
                  (reg725 ^~ reg655)})));
            end
          else
            begin
              reg726 <= (8'ha3);
              reg730 = $unsigned(reg716);
              reg731 <= reg635;
              reg732 = $signed($unsigned((($unsigned(reg714) >> $unsigned(wire544)) * reg725[(1'h1):(1'h0)])));
              reg733 = (&reg675[(5'h1f):(5'h1b)]);
              reg734 <= (~(reg626[(4'h9):(3'h5)] <<< {reg733[(4'he):(1'h0)],
                  ({reg707, reg718} ?
                      $signed(reg608) : (reg611 ? reg672 : reg647)),
                  reg594[(4'h8):(2'h2)]}));
            end
          reg735 = reg696[(1'h0):(1'h0)];
          if ((-(reg732 ?
              ($unsigned(wire545[(1'h0):(1'h0)]) ^~ (reg722[(3'h5):(1'h0)] <= $unsigned(reg694))) : $unsigned(((reg695 == reg717) - reg653)))))
            begin
              reg736 <= reg590;
              reg737 = ($signed(reg635) ?
                  $signed(reg666[(3'h7):(1'h0)]) : ((-($unsigned(reg606) ?
                          reg734[(4'h9):(2'h2)] : (-reg675))) ?
                      $unsigned($signed(reg722[(4'hf):(4'hd)])) : reg706[(3'h4):(1'h0)]));
            end
          else
            begin
              reg737 = reg635[(4'hb):(2'h3)];
              reg738 = (forvar713 >> (+((forvar713[(2'h2):(1'h0)] ^ reg626[(4'hf):(4'hd)]) || {(^reg588),
                  ((7'h4a) ? reg682 : (7'h54))})));
              reg739 = $signed(reg687[(5'h10):(4'hb)]);
              reg740 = reg573;
              reg741 <= ($signed(reg584[(1'h1):(1'h0)]) >> reg617);
              reg742 <= ($signed($signed((((7'h41) <<< reg728) || reg698[(3'h4):(2'h3)]))) ?
                  $signed((-{$signed(reg692),
                      (reg726 | wire544),
                      $signed(reg657)})) : reg682);
              reg743 <= forvar713;
            end
          for (forvar744 = (1'h0); (forvar744 < (2'h2)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 = $signed(((|reg670[(2'h2):(1'h0)]) ?
                  reg742[(1'h1):(1'h0)] : (~&$unsigned(reg612[(3'h5):(3'h5)]))));
              reg746 = (~|{(reg692 ?
                      reg582[(2'h2):(2'h2)] : reg584[(1'h1):(1'h0)]),
                  ((reg611[(2'h2):(2'h2)] >> reg626[(1'h1):(1'h1)]) ~^ reg697),
                  {$signed(reg737), $unsigned((7'h4d))}});
              reg747 = $signed($signed($signed($signed((wire547 ?
                  reg666 : reg690)))));
              reg748 <= reg723;
              reg749 = (-($signed($signed($signed(reg690))) ?
                  $signed($signed($unsigned((8'ha5)))) : ({(~reg670),
                      reg647[(1'h1):(1'h0)]} | $signed($signed((7'h47))))));
              reg750 <= (reg566 ?
                  $unsigned((reg590[(5'h13):(5'h13)] ^ reg720)) : (&reg739));
            end
          for (forvar751 = (1'h0); (forvar751 < (3'h5)); forvar751 = (forvar751 + (1'h1)))
            begin
              reg752 <= ((8'hb3) ?
                  ((+((+(8'ha9)) << (reg740 ?
                      reg604 : reg679))) + (~^$unsigned($unsigned(reg695)))) : reg692);
              reg753 <= (~$unsigned(({reg601[(4'he):(4'ha)],
                  (^~reg733),
                  reg708[(2'h2):(1'h1)]} <= $unsigned((reg590 + reg739)))));
              reg754 = reg749[(2'h2):(2'h2)];
            end
        end
      else
        begin
          if (reg741)
            begin
              reg716 <= (((~(forvar744[(3'h7):(2'h3)] && (~^reg734))) & {{reg653,
                          {reg601, (8'ha1)}},
                      $signed((reg639 ? reg589 : reg647)),
                      {(reg725 - reg715)}}) ?
                  {$unsigned((reg690 ~^ (^reg732))),
                      $signed(((^~reg753) != $signed(reg736))),
                      $unsigned((reg736 >> (reg736 ?
                          reg601 : reg723)))} : reg743[(3'h6):(1'h0)]);
              reg719 <= {($unsigned(reg707[(5'h1f):(4'hb)]) < wire546[(4'h9):(3'h4)]),
                  ((+(reg752[(4'hf):(3'h4)] ?
                      (reg596 >= reg613) : $signed(reg730))) != $unsigned(((~reg725) ?
                      (reg754 << reg702) : reg692))),
                  (+$signed((+$signed(reg653))))};
              reg720 <= (8'ha2);
              reg722 <= (~|(wire545[(1'h0):(1'h0)] == $unsigned(reg657)));
              reg723 = (8'haf);
              reg724 = $unsigned(reg742[(4'h8):(3'h4)]);
              reg726 <= {reg703[(4'hb):(4'hb)], reg679, (7'h40)};
            end
          else
            begin
              reg717 = (((-$signed($signed(reg668))) == {($signed((8'ha5)) ?
                      (!(7'h56)) : $unsigned(reg722))}) != reg727);
            end
          reg727 <= {$unsigned((reg715 << reg562[(3'h5):(3'h5)]))};
          for (forvar728 = (1'h0); (forvar728 < (3'h5)); forvar728 = (forvar728 + (1'h1)))
            begin
              reg729 <= (^~$unsigned({reg618[(4'ha):(3'h5)],
                  (+{reg696, (8'h9f), (7'h46)})}));
              reg731 <= $signed((reg581 != reg730[(3'h4):(1'h0)]));
            end
          reg732 = {{(|reg672), reg590}, (!$signed(reg714[(4'h8):(2'h3)]))};
          reg734 <= ($signed($unsigned((+reg738))) ?
              (8'hbf) : $unsigned($signed((+$unsigned(reg670)))));
          reg736 <= (|(reg675[(5'h1f):(5'h1e)] ?
              ({reg626[(3'h4):(1'h0)],
                  (~reg611)} << reg732[(5'h19):(5'h14)]) : $unsigned($signed($unsigned(wire546)))));
        end
      if ($signed(({(reg704 <= $signed(reg717))} ?
          $signed($signed($unsigned((7'h43)))) : reg707)))
        begin
          reg755 <= ((^($unsigned((^reg703)) ?
              $unsigned({reg718,
                  reg687,
                  forvar744}) : (~|$signed((8'hb5))))) ~^ (reg598 ?
              (reg657 >= ($unsigned(reg688) != (reg735 & reg722))) : reg687[(4'ha):(4'h9)]));
          for (forvar756 = (1'h0); (forvar756 < (2'h2)); forvar756 = (forvar756 + (1'h1)))
            begin
              reg757 = reg590;
            end
        end
      else
        begin
          for (forvar755 = (1'h0); (forvar755 < (3'h4)); forvar755 = (forvar755 + (1'h1)))
            begin
              reg756 <= $signed(reg601[(4'hb):(2'h3)]);
              reg757 = {(reg745 ?
                      reg590[(5'h10):(5'h10)] : ($unsigned((reg695 != reg679)) ?
                          (~&$signed(reg656)) : ({reg742} ?
                              (-reg742) : (7'h48)))),
                  reg618};
              reg758 = reg730[(1'h0):(1'h0)];
              reg759 = {forvar744};
              reg760 = reg632;
            end
          reg761 = ({(~reg731),
                  $signed({(reg588 ? reg582 : reg717), wire579}),
                  reg734[(4'hb):(2'h2)]} ?
              (~&$signed({(~|(8'hb4)),
                  reg704[(3'h6):(3'h4)],
                  (reg653 ?
                      reg606 : reg722)})) : (wire545[(1'h1):(1'h1)] ~^ (7'h4f)));
          for (forvar762 = (1'h0); (forvar762 < (1'h1)); forvar762 = (forvar762 + (1'h1)))
            begin
              reg763 <= reg661[(4'h8):(2'h3)];
              reg764 = $unsigned(reg595[(2'h3):(2'h2)]);
              reg765 = $signed((~|(~|{$unsigned((7'h4d))})));
              reg766 <= (((forvar756 ?
                  $unsigned((reg682 ? (8'hbd) : forvar744)) : ($signed(reg596) ?
                      reg590[(5'h11):(4'he)] : (reg682 && reg605))) < ($signed({reg606,
                      reg693,
                      reg720}) ?
                  $signed((reg721 ?
                      forvar751 : (7'h52))) : reg728)) * ($unsigned(reg595) < ((wire636[(5'h11):(4'hd)] && reg700) && ($unsigned(reg707) & reg736))));
              reg767 <= (-(7'h45));
              reg768 <= ($signed((reg746[(5'h13):(1'h0)] || ((reg759 >> reg605) ?
                      $signed(reg612) : (reg584 ? reg590 : reg672)))) ?
                  $signed(forvar728[(5'h16):(4'hc)]) : reg704[(2'h3):(2'h2)]);
              reg769 <= reg720;
            end
          if ((^$signed($unsigned((^reg757)))))
            begin
              reg770 = (8'h9c);
              reg771 = $signed(reg757[(5'h10):(1'h0)]);
              reg772 <= $unsigned(reg707[(5'h16):(4'hd)]);
              reg773 = ($unsigned((($signed((8'ha2)) ^~ reg590[(4'hb):(1'h0)]) + (~&$unsigned((7'h40))))) ?
                  (+reg698[(2'h3):(2'h2)]) : ({$unsigned((8'ha2))} ?
                      {(-reg595)} : $signed(reg693[(4'hf):(1'h1)])));
            end
          else
            begin
              reg772 <= ((reg618[(3'h5):(1'h0)] ?
                  $unsigned(reg729) : ((reg729 - $signed(reg565)) << $signed((~&reg670)))) << reg562[(3'h7):(2'h2)]);
              reg773 = {({$signed(reg710[(2'h2):(1'h1)]),
                      reg720,
                      (+(~reg738))} <= $unsigned(forvar728[(5'h1a):(5'h17)]))};
              reg774 = $signed($unsigned(({$unsigned(reg750),
                      $unsigned(reg578)} ?
                  reg697 : (((7'h56) ? (7'h4f) : reg672) ?
                      $unsigned(reg741) : $unsigned(reg734)))));
              reg775 = $signed({{$unsigned({reg687, reg735, reg749})},
                  $signed($signed((reg719 | reg682))),
                  $signed(reg728)});
              reg776 = (^reg605[(5'h12):(3'h7)]);
              reg777 <= reg755[(1'h0):(1'h0)];
            end
        end
      for (forvar778 = (1'h0); (forvar778 < (2'h2)); forvar778 = (forvar778 + (1'h1)))
        begin
          reg779 <= (7'h58);
          reg780 <= reg619;
          for (forvar781 = (1'h0); (forvar781 < (3'h6)); forvar781 = (forvar781 + (1'h1)))
            begin
              reg782 <= {wire544,
                  (-(reg738 && $unsigned($unsigned(reg667)))),
                  reg598[(3'h5):(3'h5)]};
              reg783 = (^~(&reg688));
              reg784 = $unsigned(($signed(reg632[(3'h6):(2'h3)]) + (~$unsigned({reg679,
                  (8'hbb)}))));
            end
          for (forvar785 = (1'h0); (forvar785 < (1'h0)); forvar785 = (forvar785 + (1'h1)))
            begin
              reg786 = $signed((($signed(((7'h4a) & reg732)) <<< $signed($unsigned(reg706))) ?
                  reg721[(4'hd):(3'h7)] : (&((reg720 > reg667) < $unsigned(reg745)))));
              reg787 <= (reg675 ?
                  ((~&reg611) <= reg748) : $signed(reg665[(4'h9):(3'h5)]));
              reg788 = ($signed($unsigned($unsigned((reg706 ?
                      reg647 : reg589)))) ?
                  reg705 : (~&(~&$unsigned($unsigned(reg702)))));
            end
          reg789 = $signed(({reg756,
              (+reg731[(4'hc):(4'hc)]),
              reg639} * $unsigned($unsigned(reg714[(3'h7):(2'h2)]))));
          for (forvar790 = (1'h0); (forvar790 < (2'h3)); forvar790 = (forvar790 + (1'h1)))
            begin
              reg791 = (^~reg698);
              reg792 <= reg683[(2'h2):(1'h1)];
              reg793 = (^$unsigned(reg716));
            end
        end
      for (forvar794 = (1'h0); (forvar794 < (3'h6)); forvar794 = (forvar794 + (1'h1)))
        begin
          if ($unsigned(reg584))
            begin
              reg795 <= reg747;
              reg796 <= (({$signed((+(7'h4e))),
                      (&(reg729 * reg708)),
                      ((wire547 >> reg647) ^~ (~^reg739))} ^~ (|reg687)) ?
                  $signed(reg578) : ({reg761,
                          ((&(8'ha5)) && (~|(7'h46))),
                          $signed((^(8'hb7)))} ?
                      (({(8'had), reg737} > reg742[(5'h10):(4'he)]) == (reg606 ?
                          (reg729 ? reg727 : reg705) : ((7'h4e) ?
                              (8'h9e) : reg709))) : $signed(((7'h4f) < reg795))));
              reg797 <= $signed($unsigned(($unsigned($unsigned(reg694)) ?
                  ($signed(wire544) ~^ $unsigned(reg666)) : reg706[(3'h7):(2'h3)])));
            end
          else
            begin
              reg795 <= (8'hb2);
              reg798 = (+{(7'h56)});
              reg799 = (~$signed($signed(reg734)));
              reg800 = (^~(reg765 + ((reg670 + $unsigned(reg793)) <= {$unsigned(reg582),
                  (reg774 >>> reg596),
                  (~|reg675)})));
              reg801 <= (reg679 ?
                  (+$unsigned(((forvar790 ? reg688 : reg779) ?
                      forvar728 : (reg741 ?
                          reg632 : reg763)))) : $unsigned(reg776));
              reg802 <= (reg691 ^~ ({reg745[(5'h10):(3'h7)],
                  forvar785,
                  (&$signed((7'h49)))} ^~ reg635));
            end
          if ($unsigned((reg595 ?
              reg593[(5'h15):(2'h2)] : ($signed((reg582 >= reg615)) ?
                  $unsigned($signed(reg739)) : $unsigned((~reg647))))))
            begin
              reg803 = $unsigned((reg776[(3'h5):(3'h4)] ?
                  {(~^(forvar744 ^ wire546)),
                      ($signed(wire545) ^~ reg756[(4'hc):(3'h4)])} : $signed(reg788[(3'h4):(1'h1)])));
              reg804 = $signed(reg723);
              reg805 = forvar755;
            end
          else
            begin
              reg806 <= $signed(($signed(forvar762[(4'hb):(3'h6)]) ?
                  $signed($signed((reg666 ?
                      reg696 : reg589))) : $unsigned($signed((reg758 ^ reg797)))));
            end
          reg807 = $signed($unsigned($signed(((reg717 != reg795) ?
              (7'h4d) : (reg726 - forvar713)))));
          reg808 = {reg656[(4'he):(4'ha)],
              reg772[(1'h1):(1'h1)],
              $unsigned((($unsigned(reg604) <= (^forvar781)) ^ $unsigned((reg760 ^ reg763))))};
          for (forvar809 = (1'h0); (forvar809 < (1'h0)); forvar809 = (forvar809 + (1'h1)))
            begin
              reg810 = $signed(($signed((forvar751 > (reg745 ?
                  (8'hb7) : reg808))) < $unsigned(forvar790)));
              reg811 <= $unsigned(($signed((8'hb0)) || (reg721[(4'hc):(2'h2)] ?
                  reg593 : ({(7'h4e), reg694} ?
                      ((7'h48) ? reg593 : reg765) : $signed(reg761)))));
            end
        end
      reg812 <= {{(reg714 | (-reg724)),
              ({$signed(reg679)} ^ reg769[(2'h2):(2'h2)]),
              reg702}};
    end
  assign wire813 = ((8'hbf) && reg769);
  assign wire814 = $unsigned($signed(($unsigned(reg711[(2'h2):(1'h1)]) > $signed((~reg578)))));
  assign wire815 = reg667;
  assign wire816 = ({reg690, $signed(reg606)} ?
                       $signed(reg734) : ({((reg598 + reg688) ?
                               {reg632,
                                   reg642,
                                   (7'h43)} : reg562[(2'h3):(2'h2)]),
                           (8'hba)} >>> reg661));
  always
    @(posedge clk) begin
      for (forvar817 = (1'h0); (forvar817 < (1'h1)); forvar817 = (forvar817 + (1'h1)))
        begin
          reg818 <= (reg795[(5'h15):(4'ha)] && ($signed((reg756 ?
                  reg706 : $unsigned(reg661))) ?
              (~^(~(~&reg593))) : (reg605 >> $signed({(8'hab), reg811}))));
          reg819 <= reg687;
          reg820 <= ((~reg682) ?
              (-$signed(reg585[(2'h2):(1'h1)])) : (&(7'h41)));
          reg821 <= $unsigned((~^$unsigned($unsigned($unsigned(reg772)))));
        end
      reg822 = (^~reg594);
      for (forvar823 = (1'h0); (forvar823 < (2'h3)); forvar823 = (forvar823 + (1'h1)))
        begin
          reg824 = $signed(($unsigned((~^(reg601 ? reg656 : reg581))) ?
              $signed($signed(reg639)) : $unsigned($unsigned($signed(reg688)))));
          if ({reg604,
              $signed(($unsigned(reg581) - ((~reg729) ?
                  (~^reg632) : (^reg665)))),
              $unsigned($signed((reg675 | $signed(reg806))))})
            begin
              reg825 <= reg702[(3'h4):(1'h0)];
              reg826 <= $unsigned((^~((^~$unsigned(reg639)) ?
                  reg766[(3'h7):(3'h7)] : ((&reg728) ?
                      ((8'ha8) | reg695) : (reg588 <<< (7'h56))))));
              reg827 = (8'hbe);
              reg828 = reg750[(4'h9):(3'h7)];
              reg829 = reg581;
            end
          else
            begin
              reg827 = (8'hbe);
              reg828 = wire636[(5'h12):(5'h11)];
              reg829 = ((reg755 ?
                      $signed({(~^reg692),
                          (&reg618)}) : wire636[(5'h1a):(5'h12)]) ?
                  $unsigned((&$unsigned((7'h43)))) : $unsigned($signed($signed((reg795 >> (7'h50))))));
              reg830 <= (~&reg584[(2'h3):(2'h3)]);
              reg831 <= (~^(reg720[(3'h5):(2'h3)] <<< (reg632[(1'h0):(1'h0)] ?
                  (&((8'hbc) ?
                      reg812 : reg687)) : ($unsigned(reg726) ^~ {(7'h4f),
                      reg596}))));
              reg832 <= ({$signed((~$signed((8'hb5)))),
                  (&reg590[(5'h14):(5'h12)])} ~^ ($signed(reg688) ?
                  reg743 : (-reg572)));
              reg833 <= (((~|(&reg601[(4'h8):(3'h6)])) ?
                  ($unsigned($signed(reg608)) ?
                      (&(wire814 ?
                          reg594 : reg701)) : reg706[(3'h7):(3'h7)]) : reg653) < $unsigned({((reg716 >> reg682) * $unsigned(reg688))}));
            end
          reg834 = (7'h4d);
        end
    end
  assign wire835 = ((reg665 & reg811[(5'h12):(4'hc)]) ?
                       reg728 : (!(reg593 ?
                           $signed(reg768) : $signed($signed((8'ha6))))));
  assign wire836 = $signed({$signed(reg777[(2'h2):(1'h0)]),
                       {(7'h51), $signed((~&reg588))},
                       reg777[(1'h1):(1'h0)]});
endmodule