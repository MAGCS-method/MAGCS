module top_1
#(parameter param411 = (8'ha3), 
parameter param412 = ((&((8'hbf) ? {(~param411), ((7'h42) > (7'h44))} : (-(~param411)))) >>> param411))
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h311):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire4;
  input wire [(5'h14):(1'h0)] wire3;
  input wire signed [(5'h13):(1'h0)] wire2;
  input wire signed [(5'h14):(1'h0)] wire1;
  input wire signed [(5'h15):(1'h0)] wire0;
  wire signed [(4'he):(1'h0)] wire403;
  wire signed [(2'h3):(1'h0)] wire402;
  wire signed [(4'he):(1'h0)] wire401;
  wire signed [(5'h10):(1'h0)] wire400;
  wire signed [(5'h13):(1'h0)] wire388;
  wire [(2'h3):(1'h0)] wire387;
  wire signed [(2'h2):(1'h0)] wire386;
  wire signed [(4'ha):(1'h0)] wire384;
  wire signed [(5'h15):(1'h0)] wire378;
  wire [(5'h15):(1'h0)] wire377;
  wire [(3'h4):(1'h0)] wire357;
  wire [(4'hf):(1'h0)] wire356;
  wire signed [(5'h15):(1'h0)] wire355;
  wire signed [(5'h10):(1'h0)] wire354;
  wire signed [(5'h15):(1'h0)] wire353;
  wire [(4'he):(1'h0)] wire171;
  wire signed [(4'hc):(1'h0)] wire351;
  reg signed [(5'h15):(1'h0)] reg410 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg409 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg407 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg405 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg404 = (1'h0);
  reg [(5'h13):(1'h0)] reg399 = (1'h0);
  reg [(5'h14):(1'h0)] reg398 = (1'h0);
  reg [(5'h15):(1'h0)] reg397 = (1'h0);
  reg [(3'h7):(1'h0)] reg396 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg395 = (1'h0);
  reg [(2'h2):(1'h0)] reg394 = (1'h0);
  reg [(5'h14):(1'h0)] reg393 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg392 = (1'h0);
  reg [(4'hd):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg390 = (1'h0);
  reg [(4'hf):(1'h0)] reg389 = (1'h0);
  reg [(5'h11):(1'h0)] reg358 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg359 = (1'h0);
  reg [(3'h4):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg361 = (1'h0);
  reg signed [(4'he):(1'h0)] reg362 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg364 = (1'h0);
  reg [(5'h15):(1'h0)] reg365 = (1'h0);
  reg [(2'h2):(1'h0)] reg366 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg367 = (1'h0);
  reg [(2'h3):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg369 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg370 = (1'h0);
  reg [(5'h12):(1'h0)] reg371 = (1'h0);
  reg [(5'h13):(1'h0)] reg372 = (1'h0);
  reg [(5'h12):(1'h0)] reg373 = (1'h0);
  reg [(5'h14):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg375 = (1'h0);
  reg [(3'h6):(1'h0)] reg376 = (1'h0);
  reg [(3'h4):(1'h0)] reg379 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg380 = (1'h0);
  reg [(2'h3):(1'h0)] reg381 = (1'h0);
  reg [(3'h7):(1'h0)] reg382 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg383 = (1'h0);
  assign y = {wire403,
                 wire402,
                 wire401,
                 wire400,
                 wire388,
                 wire387,
                 wire386,
                 wire384,
                 wire378,
                 wire377,
                 wire357,
                 wire356,
                 wire355,
                 wire354,
                 wire353,
                 wire171,
                 wire351,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg358,
                 reg359,
                 reg360,
                 reg361,
                 reg362,
                 reg363,
                 reg364,
                 reg365,
                 reg366,
                 reg367,
                 reg368,
                 reg369,
                 reg370,
                 reg371,
                 reg372,
                 reg373,
                 reg374,
                 reg375,
                 reg376,
                 reg379,
                 reg380,
                 reg381,
                 reg382,
                 reg383,
                 (1'h0)};
  module5_1 #() modinst172 (wire171, clk, wire0, wire3, wire4, wire2, wire1);
  module173_1 #() modinst352 (wire351, clk, wire171, wire0, wire4, wire3, wire2);
  assign wire353 = {$signed($signed(wire4[(1'h0):(1'h0)])),
                       (((wire4 << wire171[(4'h8):(1'h0)]) ?
                               ((8'hbf) << wire4[(5'h12):(4'ha)]) : $signed(((8'hb9) | wire2))) ?
                           (~&wire3[(4'h9):(3'h5)]) : $unsigned($unsigned($signed(wire3))))};
  assign wire354 = ((({$unsigned((8'haf))} <= {(wire0 ? wire2 : wire353)}) ?
                       $signed((wire353 + ((8'haa) << wire351))) : {$unsigned(wire351)}) || (((wire1[(5'h12):(3'h7)] ?
                               $unsigned((8'hb3)) : $signed(wire353)) ?
                           (wire351[(1'h0):(1'h0)] ?
                               wire171[(1'h0):(1'h0)] : (wire171 ?
                                   wire353 : wire1)) : $signed($signed(wire2))) ?
                       wire353[(5'h10):(2'h2)] : (($unsigned((8'h9d)) ?
                               (7'h42) : wire2) ?
                           $signed(wire0) : (+(wire2 ? (8'haf) : wire4)))));
  assign wire355 = wire0;
  assign wire356 = (8'hb7);
  assign wire357 = (~^$unsigned((-(&wire353))));
  always
    @(posedge clk) begin
      reg358 <= {$unsigned($unsigned((^wire356[(1'h1):(1'h1)])))};
      reg359 <= $unsigned($unsigned(wire353[(4'h8):(4'h8)]));
      reg360 <= {((wire351 ?
                  ((&wire1) ?
                      (wire355 ?
                          reg358 : wire355) : (wire353 * reg359)) : $signed($signed(wire356))) ?
              $signed((|wire1)) : (&($signed((7'h44)) ?
                  (&wire171) : {(8'h9e), wire171}))),
          wire354[(4'he):(4'h8)]};
      reg361 <= wire356;
      reg362 <= $signed({wire355[(4'hc):(1'h1)],
          (~&$unsigned((wire3 ? wire356 : reg361)))});
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned($signed((~^(wire353 ? wire3 : wire1))))))
        begin
          reg363 <= (-$signed({((~|wire353) || {wire3, wire4})}));
          reg364 <= (wire356 <<< wire4);
          reg365 <= ($unsigned(reg360[(2'h3):(1'h0)]) ?
              $signed((($signed(wire1) ?
                  (^wire357) : wire356[(1'h0):(1'h0)]) || wire0)) : $unsigned(reg360));
          reg366 <= (|$signed($signed({reg361, $signed(wire356)})));
        end
      else
        begin
          if ($signed((wire171 ?
              (~&$unsigned($unsigned(reg363))) : wire353[(5'h11):(4'hc)])))
            begin
              reg363 <= wire1[(4'h8):(3'h6)];
              reg364 <= ($unsigned((!$signed($signed(reg362)))) ?
                  wire353 : $signed(wire356[(4'ha):(4'h9)]));
            end
          else
            begin
              reg363 <= wire1[(4'h8):(2'h2)];
              reg364 <= (wire3[(5'h11):(4'h9)] ?
                  {$unsigned($signed((+reg366))),
                      $signed(wire4)} : wire1[(4'hb):(4'h8)]);
            end
          reg365 <= wire171;
          if ((~(($unsigned($signed(reg364)) ?
                  ((reg364 ? reg361 : (8'ha6)) ?
                      (^wire171) : (^~wire4)) : (^~(reg359 || reg364))) ?
              $unsigned(((wire4 ? wire353 : reg360) ?
                  reg366[(1'h1):(1'h1)] : wire4[(4'he):(1'h1)])) : $signed($unsigned((~&wire357))))))
            begin
              reg366 <= wire355;
              reg367 <= ($unsigned((&((reg362 ?
                      reg359 : wire2) - $signed(reg365)))) ?
                  (reg366[(1'h0):(1'h0)] | $signed($unsigned((wire3 ?
                      wire353 : reg360)))) : wire355[(5'h10):(5'h10)]);
              reg368 <= $signed($signed(((^~(wire3 & reg358)) - wire357[(1'h0):(1'h0)])));
            end
          else
            begin
              reg366 <= wire2;
            end
          if ({(($signed($unsigned((8'hb5))) ?
                      wire351[(3'h4):(3'h4)] : $unsigned($signed((7'h43)))) ?
                  $signed(((reg364 ?
                      wire171 : reg365) && (reg359 * wire2))) : {(&$unsigned(wire353))}),
              $unsigned(reg358)})
            begin
              reg369 <= $unsigned(($signed($unsigned(wire1)) ?
                  (($unsigned(reg358) ?
                      (reg358 ?
                          reg364 : wire357) : (~(8'hbc))) & reg368[(1'h0):(1'h0)]) : ($signed(((7'h40) - reg363)) <<< $unsigned($signed(reg358)))));
            end
          else
            begin
              reg369 <= (($signed($signed({wire1, wire171})) ?
                      (~&{reg367[(2'h2):(2'h2)], (&reg367)}) : reg363) ?
                  $unsigned((&$unsigned(reg368[(2'h3):(1'h0)]))) : (~^wire356));
              reg370 <= ((reg366 ~^ wire355[(3'h5):(1'h1)]) | $unsigned($unsigned(wire1[(3'h4):(1'h0)])));
              reg371 <= (wire3[(4'hc):(4'ha)] ?
                  reg364[(4'hb):(3'h7)] : ((reg370[(3'h7):(1'h0)] ?
                          $unsigned((8'ha0)) : $unsigned(reg369)) ?
                      ($signed($unsigned(wire2)) == ((wire4 < wire354) <= wire357[(3'h4):(1'h0)])) : $signed((|wire353))));
              reg372 <= (^~$unsigned($unsigned(({wire1} | {reg368}))));
            end
          reg373 <= (($unsigned(($unsigned(wire353) == $signed(wire353))) ?
                  ((~(wire0 ? (8'h9d) : wire1)) ?
                      $signed({reg361,
                          (8'hb1)}) : (+$signed(wire4))) : {$signed(reg372),
                      ((|reg362) >= wire353)}) ?
              (($signed($unsigned((8'haf))) > {{wire354, wire354},
                  ((8'hb6) << wire355)}) - $unsigned({wire0})) : ({(reg365 ?
                          $signed(reg359) : (|wire2)),
                      wire0} ?
                  {(~^(wire354 && reg368))} : (+(-$unsigned(wire4)))));
        end
      if ({(&{wire356[(4'h8):(3'h6)],
              ((wire3 && wire356) ? $unsigned(wire4) : $signed(wire351))}),
          {{($signed(wire2) ? {wire353} : (reg368 ? reg368 : reg366))}}})
        begin
          reg374 <= $unsigned(wire3[(4'he):(1'h0)]);
        end
      else
        begin
          reg374 <= (-(~^reg359));
        end
      reg375 <= (($signed(reg358[(1'h0):(1'h0)]) ?
              $signed((((8'hbb) >= (8'ha0)) ?
                  {reg372} : (~reg360))) : {$signed(((8'ha0) ?
                      reg360 : wire1))}) ?
          wire3 : $unsigned({$unsigned((8'hba))}));
      reg376 <= $signed(((~^(+$unsigned(wire353))) < (wire0 ?
          $unsigned($unsigned(wire2)) : $signed((^~reg373)))));
    end
  assign wire377 = (8'ha8);
  assign wire378 = {(wire351 ?
                           $signed({reg367[(1'h1):(1'h0)],
                               $unsigned(wire357)}) : ((^$unsigned(wire354)) ?
                               reg373 : (~|wire2)))};
  always
    @(posedge clk) begin
      reg379 <= ($signed(($signed((reg368 >= reg359)) ?
          ((|reg375) ^ $signed(wire353)) : $unsigned(reg372))) && {{($unsigned(reg369) ?
                  $signed((8'hb9)) : reg368),
              $unsigned(reg373[(4'hc):(3'h6)])},
          ({$unsigned(reg364)} ?
              ({reg363, wire2} ?
                  ((8'hb4) ?
                      wire355 : reg370) : (wire353 - reg358)) : reg365)});
      reg380 <= wire3;
      reg381 <= ($unsigned((&reg361)) ?
          $signed({(^$unsigned((7'h42)))}) : (wire356[(4'hd):(3'h4)] ?
              (($unsigned(wire1) == (wire351 >= wire354)) ?
                  reg371 : $signed(wire355[(4'h9):(3'h6)])) : wire355[(1'h0):(1'h0)]));
      reg382 <= $unsigned(((~&reg366[(1'h0):(1'h0)]) && (((reg380 ?
          reg375 : reg369) && (wire378 - reg367)) <<< $unsigned(reg373[(2'h2):(1'h1)]))));
      reg383 <= ($signed(reg376) >>> wire1[(4'hb):(4'h9)]);
    end
  module5_1 #() modinst385 (.wire7(reg359), .clk(clk), .wire10(wire377), .y(wire384), .wire9(reg372), .wire6(wire0), .wire8(reg363));
  assign wire386 = $signed($unsigned(((7'h41) ? reg372 : wire2)));
  assign wire387 = $unsigned((8'hb4));
  assign wire388 = (~({$unsigned(wire384[(4'ha):(4'ha)])} ?
                       (~reg373[(2'h3):(2'h2)]) : $unsigned(wire356[(3'h4):(3'h4)])));
  always
    @(posedge clk) begin
      if ((~(({wire384, reg371[(4'hc):(2'h3)]} >> reg372[(4'h9):(3'h5)]) ?
          ({wire351[(4'hc):(3'h6)],
              (+reg369)} ~^ reg369[(5'h10):(2'h2)]) : $unsigned(($signed(wire0) ^~ (^reg364))))))
        begin
          reg389 <= $signed(((~|(8'haf)) ?
              ((reg360 ? $signed(reg371) : $signed(reg359)) ?
                  wire357[(3'h4):(1'h1)] : reg365[(5'h14):(3'h7)]) : (!(~^$unsigned(wire378)))));
          reg390 <= $unsigned((^wire387[(1'h1):(1'h0)]));
          reg391 <= wire4[(4'hf):(4'ha)];
          reg392 <= ((|wire1[(4'he):(4'he)]) ^~ $signed(wire355));
        end
      else
        begin
          if ((reg389 ?
              {(($signed(reg361) & wire377) <<< wire351[(3'h5):(2'h2)]),
                  {$unsigned($unsigned(reg370)),
                      ($signed((8'hb1)) ?
                          (wire171 | wire388) : (wire355 >>> wire353))}} : reg362))
            begin
              reg389 <= reg364[(5'h11):(5'h10)];
              reg390 <= reg363[(4'hd):(3'h6)];
            end
          else
            begin
              reg389 <= wire1[(1'h0):(1'h0)];
              reg390 <= $signed($unsigned(reg374[(4'h8):(1'h1)]));
              reg391 <= (+((reg392 ?
                      reg389 : ($signed((8'had)) ~^ wire384[(4'h8):(4'h8)])) ?
                  (~|wire354[(4'he):(4'h9)]) : $signed(((-reg381) ?
                      $unsigned(wire353) : wire351[(1'h1):(1'h0)]))));
            end
        end
      if ($signed($unsigned((reg374[(1'h1):(1'h0)] ~^ reg383[(1'h0):(1'h0)]))))
        begin
          reg393 <= $signed(reg382[(3'h4):(3'h4)]);
        end
      else
        begin
          reg393 <= {(+(reg391[(4'h8):(1'h1)] >> (|wire4[(4'h9):(3'h4)])))};
          reg394 <= ($signed($signed(reg392[(3'h5):(2'h3)])) ?
              (8'h9d) : $unsigned(reg369[(4'he):(1'h0)]));
          reg395 <= ((((~((8'ha0) ? reg369 : (8'ha3))) ?
              reg372 : reg381[(2'h2):(1'h1)]) <= reg392) && $signed($signed(($signed(wire377) <= {reg379}))));
          reg396 <= $signed((~^$signed(((reg392 + (8'h9e)) ?
              (reg358 ? reg367 : wire4) : (reg376 >>> (8'hae))))));
          if ({wire355, $signed($signed($signed((~&(8'hb5)))))})
            begin
              reg397 <= (($signed({reg395[(4'hb):(1'h0)]}) ?
                      ((!(8'ha5)) >>> (~|(^reg381))) : reg359) ?
                  reg358 : ({$signed((reg395 <<< reg364)), (!$signed(reg383))} ?
                      reg380 : $unsigned($unsigned((reg395 && (8'hb4))))));
              reg398 <= ((|reg392[(1'h0):(1'h0)]) ?
                  (((wire354 ?
                      (reg361 ?
                          reg382 : reg361) : (^~reg376)) >>> wire387) ^ (((reg369 ?
                          wire386 : reg362) | (-wire378)) ?
                      (^~(8'hac)) : $signed($unsigned((8'hbf))))) : $unsigned((8'ha9)));
            end
          else
            begin
              reg397 <= wire1;
              reg398 <= reg398;
            end
        end
      reg399 <= $unsigned(reg366[(1'h0):(1'h0)]);
    end
  assign wire400 = $signed({(-$unsigned(reg367))});
  assign wire401 = wire356;
  assign wire402 = {$signed(wire354),
                       ({$signed((reg393 < wire386)),
                           wire2[(3'h6):(3'h5)]} < $unsigned($unsigned((wire355 >>> wire3))))};
  assign wire403 = wire171[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg404 <= reg397[(5'h11):(5'h11)];
      reg405 <= reg372[(5'h12):(2'h2)];
      reg406 <= reg364[(5'h10):(4'h9)];
      if (wire171)
        begin
          reg407 <= $unsigned($unsigned(wire1[(4'he):(3'h5)]));
          reg408 <= wire351[(2'h3):(1'h1)];
          reg409 <= reg368;
          reg410 <= $signed(reg364);
        end
      else
        begin
          reg407 <= (^wire4[(5'h10):(3'h4)]);
          if (reg394)
            begin
              reg408 <= (~&(($unsigned($signed(reg363)) > {reg395,
                  (wire171 ? reg399 : reg362)}) ^ $unsigned(((&reg394) ?
                  $unsigned((8'hb7)) : $unsigned(wire1)))));
            end
          else
            begin
              reg408 <= $signed(({wire171[(4'he):(4'hc)]} ?
                  {(8'hb6)} : reg409[(3'h4):(1'h0)]));
            end
          reg409 <= $signed($signed($signed(((reg375 ? reg398 : wire403) ?
              {reg368} : $unsigned((8'had))))));
        end
    end
endmodule

module module173_1  (y, clk, wire174, wire175, wire176, wire177, wire178);
  output wire [(32'h21f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire174;
  input wire signed [(4'h9):(1'h0)] wire175;
  input wire [(5'h14):(1'h0)] wire176;
  input wire [(5'h14):(1'h0)] wire177;
  input wire signed [(5'h13):(1'h0)] wire178;
  wire signed [(4'h9):(1'h0)] wire350;
  wire signed [(4'hc):(1'h0)] wire349;
  wire [(5'h10):(1'h0)] wire333;
  wire [(4'he):(1'h0)] wire273;
  wire signed [(5'h11):(1'h0)] wire228;
  wire [(2'h3):(1'h0)] wire227;
  wire [(2'h3):(1'h0)] wire226;
  wire [(5'h13):(1'h0)] wire212;
  wire [(5'h10):(1'h0)] wire211;
  wire [(3'h4):(1'h0)] wire210;
  wire [(5'h14):(1'h0)] wire209;
  wire signed [(5'h11):(1'h0)] wire179;
  wire [(5'h12):(1'h0)] wire180;
  wire [(4'hc):(1'h0)] wire181;
  wire [(5'h11):(1'h0)] wire182;
  wire signed [(4'ha):(1'h0)] wire207;
  wire [(2'h3):(1'h0)] wire275;
  wire signed [(5'h11):(1'h0)] wire276;
  wire [(2'h3):(1'h0)] wire277;
  wire [(3'h5):(1'h0)] wire331;
  reg [(4'hd):(1'h0)] reg348 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg347 = (1'h0);
  reg [(2'h3):(1'h0)] reg346 = (1'h0);
  reg [(5'h15):(1'h0)] reg345 = (1'h0);
  reg [(4'h9):(1'h0)] reg344 = (1'h0);
  reg [(5'h15):(1'h0)] reg343 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg342 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg341 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg340 = (1'h0);
  reg [(4'hf):(1'h0)] reg339 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg338 = (1'h0);
  reg [(3'h6):(1'h0)] reg337 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg336 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg334 = (1'h0);
  reg [(2'h3):(1'h0)] reg213 = (1'h0);
  reg [(5'h12):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg216 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg217 = (1'h0);
  reg signed [(4'he):(1'h0)] reg218 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg220 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg221 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg222 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg223 = (1'h0);
  reg [(5'h14):(1'h0)] reg224 = (1'h0);
  reg [(4'hb):(1'h0)] reg225 = (1'h0);
  assign y = {wire350,
                 wire349,
                 wire333,
                 wire273,
                 wire228,
                 wire227,
                 wire226,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 wire179,
                 wire180,
                 wire181,
                 wire182,
                 wire207,
                 wire275,
                 wire276,
                 wire277,
                 wire331,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg213,
                 reg214,
                 reg215,
                 reg216,
                 reg217,
                 reg218,
                 reg219,
                 reg220,
                 reg221,
                 reg222,
                 reg223,
                 reg224,
                 reg225,
                 (1'h0)};
  assign wire179 = $unsigned(wire174);
  assign wire180 = (+wire176);
  assign wire181 = (^wire176);
  assign wire182 = (($unsigned(wire176) ? wire179 : $unsigned(wire175)) ?
                       (wire181[(3'h4):(1'h1)] == $unsigned(wire179[(1'h1):(1'h1)])) : (+wire178[(4'hf):(4'hf)]));
  module183_1 #() modinst208 (wire207, clk, wire181, wire174, wire179, wire177, wire182);
  assign wire209 = wire175;
  assign wire210 = $signed(({{$signed(wire180),
                           (^wire180)}} == $signed(wire209)));
  assign wire211 = {(wire181[(3'h5):(1'h0)] ?
                           $signed($signed(wire176)) : wire178[(4'hd):(4'hd)])};
  assign wire212 = ($signed($unsigned(wire181)) ?
                       $unsigned($unsigned((8'hbb))) : {wire207[(4'h8):(2'h2)]});
  always
    @(posedge clk) begin
      reg213 <= (+(wire180[(3'h5):(2'h3)] ?
          wire179[(3'h7):(3'h5)] : ($unsigned((wire182 ?
              wire209 : wire212)) & wire209)));
      reg214 <= ($signed($unsigned((^~((8'hb7) || wire177)))) ?
          (($signed($signed(wire176)) >>> wire211) ?
              (^((+wire180) == $signed(wire182))) : (~^wire211)) : wire211);
      reg215 <= (wire210 ~^ $unsigned((wire182[(4'h8):(3'h7)] & $unsigned(((8'hbb) ~^ wire212)))));
      if (wire179[(3'h6):(3'h5)])
        begin
          if ($unsigned((!wire209[(4'h9):(3'h5)])))
            begin
              reg216 <= (-(~$unsigned(reg214)));
              reg217 <= $signed((8'hab));
              reg218 <= ((~^{$unsigned((-reg213)),
                  (+(wire209 ?
                      wire178 : (8'hb2)))}) & (~&wire211[(4'hd):(4'hd)]));
            end
          else
            begin
              reg216 <= wire182[(4'hf):(2'h3)];
              reg217 <= (8'hb4);
              reg218 <= $unsigned((!(reg218 ^~ ($unsigned(wire210) ?
                  wire175 : (8'ha8)))));
              reg219 <= wire182[(4'hb):(1'h0)];
              reg220 <= wire211;
            end
        end
      else
        begin
          reg216 <= (($signed(($signed(wire211) < reg220)) ?
              $unsigned(((&wire174) || ((7'h44) == (8'ha2)))) : (({reg215,
                          wire209} ?
                      (reg218 | wire176) : reg218[(3'h5):(2'h3)]) ?
                  wire212[(4'hc):(2'h2)] : (&wire207))) != (|(wire207 + ($unsigned(reg217) ?
              $unsigned((8'hae)) : reg219[(3'h5):(2'h3)]))));
          reg217 <= {(^$unsigned(((~wire181) >>> (+reg217))))};
          if (reg214[(2'h2):(1'h0)])
            begin
              reg218 <= ((~|reg219[(2'h2):(1'h0)]) ^ $signed((-($unsigned((8'hb7)) ?
                  (reg218 ? reg219 : wire182) : $signed(reg217)))));
              reg219 <= wire207[(4'h9):(1'h1)];
              reg220 <= (+(wire209[(2'h3):(2'h2)] ~^ wire178[(5'h13):(4'hd)]));
              reg221 <= wire210;
              reg222 <= ({((+$unsigned(wire210)) ?
                          $unsigned((wire174 ?
                              reg217 : (8'haa))) : ($signed(wire209) ?
                              wire182[(2'h3):(1'h1)] : {wire175})),
                      reg218[(4'hb):(4'h9)]} ?
                  (((8'hae) ?
                          {$unsigned((8'hb8)),
                              ((8'hb2) ? reg214 : wire181)} : wire175) ?
                      ($unsigned($signed(wire181)) && ($signed(wire179) ?
                          wire174 : $signed(wire211))) : {((!reg220) << (wire209 || wire178))}) : $unsigned(wire179));
            end
          else
            begin
              reg218 <= (^~((8'had) ?
                  ($unsigned(wire211[(4'hb):(3'h6)]) ?
                      (reg219[(4'h9):(3'h6)] | reg220[(4'hf):(3'h5)]) : (wire174 ?
                          reg220[(5'h10):(2'h3)] : (reg214 ?
                              wire182 : (8'ha2)))) : $unsigned($unsigned((~&(7'h44))))));
              reg219 <= ((!reg214[(3'h4):(1'h1)]) ?
                  reg214[(2'h2):(1'h0)] : ((((wire177 >>> wire210) > wire179) ?
                          wire175[(4'h8):(3'h6)] : (~reg220)) ?
                      (&(^$unsigned(reg219))) : wire179));
              reg220 <= ($signed((((8'hb2) ?
                          reg219[(3'h5):(3'h5)] : $signed(wire174)) ?
                      reg216 : (~^(^reg213)))) ?
                  ((~&((reg220 * wire175) || (8'ha5))) ?
                      {{(wire174 ?
                                  wire174 : (8'had))}} : reg222) : {(($signed(reg220) ?
                          $unsigned(wire181) : reg214) & (reg219[(3'h4):(1'h0)] < (wire181 ?
                          wire181 : (7'h41))))});
              reg221 <= $signed((~&$signed((~&wire209[(5'h12):(1'h1)]))));
              reg222 <= (~|$signed(($unsigned($unsigned(wire181)) ?
                  (^~$unsigned((8'hae))) : ((~^(8'h9c)) ?
                      wire178 : (reg222 ^~ wire182)))));
            end
          reg223 <= ($unsigned((7'h41)) || reg215);
          reg224 <= $unsigned((~^$signed($unsigned($unsigned(reg220)))));
        end
      reg225 <= ((reg219[(4'h9):(3'h7)] ? (wire181 << (8'hb2)) : (8'ha1)) ?
          wire179 : (|wire176[(1'h1):(1'h0)]));
    end
  assign wire226 = $signed(reg224);
  assign wire227 = (wire226 != (^~reg213));
  assign wire228 = wire182[(1'h0):(1'h0)];
  module229_1 #() modinst274 (.wire232(reg224), .wire233(reg218), .clk(clk), .wire230(wire176), .y(wire273), .wire231(reg222));
  assign wire275 = wire209;
  assign wire276 = ($unsigned($unsigned($signed({wire177}))) && $unsigned(reg217[(1'h1):(1'h1)]));
  assign wire277 = ($unsigned((+$unsigned($signed(wire179)))) <= $signed({(8'ha5)}));
  module278_1 #() modinst332 (wire331, clk, reg225, reg220, wire174, reg221, reg214);
  assign wire333 = {$unsigned(((~|reg221) && {reg224[(3'h4):(2'h2)], reg218})),
                       $unsigned(wire209[(5'h12):(4'ha)])};
  always
    @(posedge clk) begin
      reg334 <= $unsigned($signed((wire228[(4'hd):(1'h0)] ?
          $unsigned((wire227 != (8'h9e))) : (^wire177[(4'hc):(3'h7)]))));
      reg335 <= reg217;
      reg336 <= $signed(wire210);
      if ($signed((wire277 <= (^~(wire179 * {reg215})))))
        begin
          reg337 <= $signed(((^wire331) ?
              reg334[(5'h13):(2'h2)] : wire227[(1'h0):(1'h0)]));
          if ($signed((($unsigned(((7'h42) ? wire277 : reg219)) ?
                  (!$unsigned((8'hbc))) : ((&wire333) ?
                      (wire212 ? (8'hac) : wire174) : $signed((8'hb3)))) ?
              reg224 : (~reg334))))
            begin
              reg338 <= (8'ha2);
              reg339 <= wire179[(5'h11):(1'h1)];
              reg340 <= wire177[(4'hc):(2'h3)];
              reg341 <= ((wire182 != {(reg214[(3'h5):(3'h4)] ?
                          (wire179 != reg225) : (|wire176))}) ?
                  $unsigned(((^~$unsigned(wire277)) ?
                      {reg339,
                          (reg219 == wire226)} : $unsigned((~^wire209)))) : (|wire174));
            end
          else
            begin
              reg338 <= reg339;
              reg339 <= reg215[(4'he):(4'h9)];
            end
        end
      else
        begin
          reg337 <= ((|reg218) != (!(reg337 == reg341[(1'h1):(1'h1)])));
          if ((((~&reg216) ?
                  {wire175, reg341} : ($signed($unsigned(wire176)) ?
                      (+reg221) : wire209)) ?
              (8'hb0) : $unsigned(((|(reg221 - reg338)) ?
                  $signed((wire182 ? reg334 : (8'ha0))) : $unsigned(wire179)))))
            begin
              reg338 <= $unsigned(wire174[(3'h7):(1'h0)]);
              reg339 <= {(reg338[(4'h9):(4'h9)] ?
                      $unsigned(((^wire212) && (~&reg216))) : ({(8'haa)} == {(reg341 ?
                              (8'hbf) : reg341),
                          (wire276 ? reg220 : reg221)}))};
            end
          else
            begin
              reg338 <= $signed($unsigned($signed($signed($signed(wire177)))));
              reg339 <= wire275[(2'h2):(1'h0)];
              reg340 <= wire207[(4'h8):(3'h6)];
              reg341 <= (reg220 ?
                  ((!((~wire277) ?
                          (reg334 == wire210) : wire177[(5'h10):(4'he)])) ?
                      (~wire275) : (^~$unsigned(wire226[(1'h0):(1'h0)]))) : (!$unsigned(reg214)));
              reg342 <= $unsigned(($signed(reg213[(1'h1):(1'h0)]) | wire275));
            end
          if (reg225)
            begin
              reg343 <= wire181;
              reg344 <= $signed(($signed({(^~(8'hb1))}) - (($unsigned(wire331) < wire228[(2'h2):(2'h2)]) ?
                  $unsigned((wire176 ?
                      reg334 : wire226)) : $unsigned($unsigned(wire174)))));
              reg345 <= (!wire276);
            end
          else
            begin
              reg343 <= reg214[(3'h5):(1'h1)];
              reg344 <= (reg224[(5'h10):(4'hd)] + $unsigned((~(+((8'ha0) != wire277)))));
            end
          reg346 <= {(($unsigned((reg343 ? reg345 : (7'h40))) ?
                      ({wire228,
                          wire210} != (wire227 && wire179)) : ((^~reg223) & (wire276 > wire180))) ?
                  {{reg215[(3'h7):(2'h3)],
                          $signed(wire276)}} : $signed($signed({reg342})))};
          reg347 <= (8'hbc);
        end
      reg348 <= $unsigned({{$signed($signed(reg346))}});
    end
  assign wire349 = ((^~wire176[(4'hd):(4'h8)]) ?
                       ($signed(reg336) ^~ (&$signed($signed(wire277)))) : reg213[(1'h0):(1'h0)]);
  assign wire350 = (((8'h9c) ?
                           reg345[(5'h15):(4'hd)] : (reg335 & ($signed((8'haf)) > (reg213 ?
                               reg220 : reg225)))) ?
                       reg337[(1'h0):(1'h0)] : ((wire176[(3'h4):(3'h4)] << {$unsigned(reg213),
                           $unsigned(wire276)}) ^~ $unsigned((&$unsigned(reg342)))));
endmodule

module module5_1  (y, clk, wire10, wire9, wire8, wire7, wire6);
  output wire [(32'h3d0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire10;
  input wire signed [(4'hf):(1'h0)] wire9;
  input wire [(4'hd):(1'h0)] wire8;
  input wire [(4'ha):(1'h0)] wire7;
  input wire signed [(5'h12):(1'h0)] wire6;
  wire signed [(4'h9):(1'h0)] wire170;
  wire signed [(5'h14):(1'h0)] wire72;
  wire [(5'h14):(1'h0)] wire12;
  wire [(5'h10):(1'h0)] wire11;
  wire signed [(5'h14):(1'h0)] wire103;
  wire [(4'hf):(1'h0)] wire134;
  wire signed [(5'h13):(1'h0)] wire135;
  wire signed [(4'hb):(1'h0)] wire152;
  wire [(4'h8):(1'h0)] wire168;
  reg [(4'h9):(1'h0)] reg151 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg150 = (1'h0);
  reg [(5'h13):(1'h0)] reg149 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg148 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg146 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg145 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg143 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg142 = (1'h0);
  reg [(3'h6):(1'h0)] reg141 = (1'h0);
  reg [(4'hb):(1'h0)] reg140 = (1'h0);
  reg [(3'h5):(1'h0)] reg139 = (1'h0);
  reg [(3'h5):(1'h0)] reg138 = (1'h0);
  reg [(3'h5):(1'h0)] reg137 = (1'h0);
  reg [(2'h3):(1'h0)] reg136 = (1'h0);
  reg [(5'h13):(1'h0)] reg133 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg132 = (1'h0);
  reg [(3'h7):(1'h0)] reg131 = (1'h0);
  reg [(4'hd):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg128 = (1'h0);
  reg [(4'hf):(1'h0)] reg127 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg125 = (1'h0);
  reg [(5'h11):(1'h0)] reg124 = (1'h0);
  reg [(4'hf):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg122 = (1'h0);
  reg [(5'h14):(1'h0)] reg121 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg120 = (1'h0);
  reg [(4'h8):(1'h0)] reg119 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg117 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg116 = (1'h0);
  reg [(3'h5):(1'h0)] reg115 = (1'h0);
  reg [(4'he):(1'h0)] reg114 = (1'h0);
  reg [(3'h5):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg112 = (1'h0);
  reg [(2'h3):(1'h0)] reg111 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg110 = (1'h0);
  reg [(3'h5):(1'h0)] reg109 = (1'h0);
  reg [(4'hd):(1'h0)] reg108 = (1'h0);
  reg [(5'h10):(1'h0)] reg107 = (1'h0);
  reg [(2'h3):(1'h0)] reg106 = (1'h0);
  reg [(4'hb):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg102 = (1'h0);
  reg [(4'h8):(1'h0)] reg101 = (1'h0);
  reg [(3'h7):(1'h0)] reg100 = (1'h0);
  reg signed [(4'he):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg98 = (1'h0);
  reg [(3'h4):(1'h0)] reg97 = (1'h0);
  reg [(3'h7):(1'h0)] reg96 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg95 = (1'h0);
  reg [(5'h13):(1'h0)] reg94 = (1'h0);
  reg [(4'hb):(1'h0)] reg93 = (1'h0);
  reg [(3'h7):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg91 = (1'h0);
  reg [(5'h11):(1'h0)] reg90 = (1'h0);
  reg [(5'h13):(1'h0)] reg89 = (1'h0);
  reg [(5'h10):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg87 = (1'h0);
  reg signed [(4'he):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg85 = (1'h0);
  reg [(4'hf):(1'h0)] reg84 = (1'h0);
  reg [(4'h9):(1'h0)] reg83 = (1'h0);
  reg signed [(4'he):(1'h0)] reg82 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg81 = (1'h0);
  reg signed [(4'he):(1'h0)] reg80 = (1'h0);
  reg [(5'h15):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg78 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg76 = (1'h0);
  reg [(4'h8):(1'h0)] reg75 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg74 = (1'h0);
  assign y = {wire170,
                 wire72,
                 wire12,
                 wire11,
                 wire103,
                 wire134,
                 wire135,
                 wire152,
                 wire168,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 (1'h0)};
  assign wire11 = wire8[(4'hb):(3'h4)];
  assign wire12 = {wire6[(3'h7):(1'h0)]};
  module13_1 #() modinst73 (.wire15(wire9), .wire17(wire11), .wire18(wire6), .wire14(wire8), .clk(clk), .y(wire72), .wire16(wire12));
  always
    @(posedge clk) begin
      reg74 <= (~(~wire72));
      if ($signed({{(|(!wire10)), reg74[(1'h1):(1'h0)]}, wire6}))
        begin
          reg75 <= $signed({$signed($signed((wire6 ? wire10 : wire6)))});
          if ({wire6, {$signed(reg74)}})
            begin
              reg76 <= (((~$unsigned({wire11,
                  (7'h43)})) + $unsigned(wire12)) ~^ (&(&reg74)));
              reg77 <= {wire7,
                  (($signed((reg76 & wire7)) < wire11) ~^ ((~|(^~wire6)) ?
                      ($unsigned(reg74) ?
                          (wire9 ?
                              (8'hbc) : reg76) : (|wire9)) : (^~((8'ha4) || wire6))))};
            end
          else
            begin
              reg76 <= (((~|{(!reg74)}) ?
                      $signed($signed($unsigned(reg74))) : {(|(~wire10)),
                          ((wire6 <= wire72) ^~ {wire9})}) ?
                  $unsigned(wire8) : (({(reg76 ?
                              (8'hb4) : wire6)} - $signed(reg75[(3'h7):(3'h6)])) ?
                      (^~(+(wire6 ?
                          wire9 : wire7))) : {($unsigned(wire7) >>> reg77[(3'h6):(1'h0)]),
                          wire10}));
              reg77 <= (&(8'ha9));
              reg78 <= $signed(wire8);
            end
          reg79 <= wire7[(4'ha):(1'h0)];
          reg80 <= $signed(reg79);
        end
      else
        begin
          reg75 <= {$signed(reg75)};
          reg76 <= $unsigned((~&wire8));
          reg77 <= $signed({(8'hb3)});
          if ((($unsigned(reg79) | $signed((+wire10))) ?
              $signed((-(reg80 ?
                  ((8'ha5) ?
                      wire12 : wire12) : (~reg80)))) : ((~|reg78[(3'h6):(3'h4)]) * (wire9 ?
                  reg76 : {$signed(wire8)}))))
            begin
              reg78 <= $unsigned(wire12);
              reg79 <= reg78;
              reg80 <= wire7;
              reg81 <= {$unsigned(reg74[(2'h2):(1'h1)])};
            end
          else
            begin
              reg78 <= (({reg77[(1'h1):(1'h1)]} >> (8'ha5)) <= (reg74[(1'h0):(1'h0)] ?
                  (~|$unsigned($unsigned(wire8))) : (((8'had) ?
                          (^reg80) : {(8'h9c), (8'hb9)}) ?
                      wire8[(3'h5):(3'h4)] : {((8'ha1) ? reg79 : wire72),
                          {wire11}})));
              reg79 <= $unsigned($unsigned(wire72[(1'h1):(1'h0)]));
              reg80 <= wire8;
              reg81 <= ($signed(((wire7[(2'h2):(1'h1)] >>> (reg74 ?
                  wire8 : reg78)) >>> (((8'ha1) ? reg75 : wire7) ?
                  (reg80 ?
                      wire7 : reg79) : reg76))) ~^ $signed({($signed((8'hbf)) && wire9)}));
              reg82 <= {(~&(|reg77))};
            end
          reg83 <= ($unsigned($signed(({wire9, (8'ha2)} ?
                  (reg82 ? reg80 : reg80) : $unsigned(reg75)))) ?
              ((wire11[(4'hd):(4'h8)] ?
                      (&wire11[(3'h6):(2'h3)]) : $unsigned($unsigned(wire10))) ?
                  $signed($signed((wire7 ?
                      (8'hbb) : (8'hbc)))) : $unsigned(wire10)) : $signed(reg74));
        end
      if ($signed($signed((((8'hbe) ^ $signed(reg83)) ?
          reg80 : $unsigned((wire10 ? wire6 : reg76))))))
        begin
          if ((-$signed(wire11)))
            begin
              reg84 <= (~|{(~^(^~{reg79, reg78}))});
              reg85 <= (8'hb8);
              reg86 <= reg85[(4'he):(4'hd)];
            end
          else
            begin
              reg84 <= $signed($unsigned(reg86));
              reg85 <= reg86;
              reg86 <= $signed(((~^reg83[(2'h3):(2'h2)]) <<< reg78[(2'h3):(1'h0)]));
              reg87 <= ({{wire7, $unsigned($unsigned(wire10))}} << wire72);
            end
          reg88 <= $signed($signed($unsigned($unsigned((~|reg77)))));
          reg89 <= reg84;
          reg90 <= (8'hb0);
          if ({wire12[(3'h4):(2'h2)], wire11})
            begin
              reg91 <= reg87[(2'h2):(1'h1)];
              reg92 <= (reg75[(4'h8):(1'h0)] ?
                  $signed($signed(wire12[(4'h8):(2'h2)])) : $signed(reg81[(3'h4):(1'h1)]));
              reg93 <= reg77;
              reg94 <= (~&wire12[(4'hc):(3'h7)]);
              reg95 <= $signed(wire12[(5'h11):(3'h5)]);
            end
          else
            begin
              reg91 <= (reg85 ?
                  {(($signed(reg85) & {reg93}) | ((^reg78) >= (reg93 | (8'hbf)))),
                      ({(~reg81),
                          reg94[(1'h1):(1'h1)]} && (~^(wire8 & reg94)))} : {wire72,
                      ($signed((~|reg88)) & $signed(wire8[(4'hc):(3'h7)]))});
              reg92 <= $unsigned((8'ha5));
              reg93 <= (~|((~&$signed(reg95)) || ((wire8[(1'h0):(1'h0)] ?
                      ((8'hb6) ? reg76 : reg82) : (reg86 < reg75)) ?
                  ((wire11 == reg78) ?
                      $unsigned((8'ha9)) : reg86[(3'h7):(3'h7)]) : ((reg87 + (8'ha3)) ?
                      (8'ha3) : (reg80 ? reg79 : (7'h43))))));
              reg94 <= $unsigned($signed(($unsigned($signed(reg86)) ?
                  (|(reg80 ? (8'ha6) : reg92)) : (reg77[(3'h4):(2'h3)] ?
                      {(7'h42)} : $unsigned(reg87)))));
            end
        end
      else
        begin
          reg84 <= reg81;
        end
      reg96 <= $signed(($signed((^~(reg87 < wire10))) >>> {$signed((reg80 ?
              reg80 : reg91))}));
      reg97 <= reg80[(4'he):(4'ha)];
    end
  always
    @(posedge clk) begin
      reg98 <= reg86;
      reg99 <= (reg81[(4'hf):(4'ha)] ^ ({((reg75 ? reg90 : wire12) ?
                  (reg85 ? reg75 : reg75) : $unsigned(reg90)),
              $unsigned($unsigned(reg79))} ?
          $signed(((&reg90) >> ((8'ha7) <<< (8'hb2)))) : $unsigned($signed((reg78 ?
              reg83 : wire72)))));
      if ((~|reg98))
        begin
          reg100 <= (wire10 * ((^~(!(reg91 ? reg89 : reg79))) ?
              $signed(reg89[(4'hf):(3'h6)]) : reg93[(4'ha):(2'h2)]));
          reg101 <= $signed(((($unsigned(wire6) ?
                  (reg75 ? reg85 : (8'hb4)) : reg86) ~^ $signed((-wire10))) ?
              (+(8'ha1)) : ({(~^(8'hb7))} ^ ((wire10 ? wire11 : reg82) ?
                  $signed(reg98) : $unsigned((8'hbd))))));
          reg102 <= $signed($signed((^~($signed(wire6) <= $signed(reg90)))));
        end
      else
        begin
          reg100 <= $signed(((8'hb3) ?
              $unsigned($unsigned($signed((8'h9f)))) : reg88));
          reg101 <= reg84;
        end
    end
  assign wire103 = ($signed({(+(8'hbb)),
                       $signed((wire72 ^ reg75))}) <<< {$unsigned(((reg84 ?
                               (7'h42) : reg85) ?
                           wire72[(4'hc):(1'h1)] : reg82[(4'he):(1'h0)])),
                       $signed((((8'hb1) <= wire72) ?
                           (reg96 == reg77) : reg83))});
  always
    @(posedge clk) begin
      if (reg93[(3'h6):(1'h1)])
        begin
          if ((reg99 ?
              $signed($signed($signed({wire10}))) : (wire11 && (!{$signed(reg98),
                  (reg83 ? reg83 : reg101)}))))
            begin
              reg104 <= ($unsigned({(~|$unsigned((8'hbf)))}) ?
                  (($unsigned($signed(wire11)) ?
                          reg88[(4'hb):(1'h0)] : (8'hb8)) ?
                      $signed($unsigned((wire9 >= wire12))) : (8'hbe)) : reg94[(4'h9):(4'h9)]);
              reg105 <= reg102;
            end
          else
            begin
              reg104 <= $signed($unsigned($unsigned(reg100)));
              reg105 <= ($signed($unsigned(((reg93 >>> wire6) << $unsigned((8'hb3))))) && reg85[(5'h13):(4'hc)]);
            end
          reg106 <= $signed((^wire10));
        end
      else
        begin
          reg104 <= {$unsigned((+($unsigned((8'ha1)) >>> (wire6 >>> reg86))))};
        end
      if (reg106[(2'h2):(1'h0)])
        begin
          if ({{($unsigned($signed(reg79)) < (wire8[(3'h4):(3'h4)] || $unsigned(reg98))),
                  $signed(($unsigned((7'h43)) <= (^~wire10)))},
              reg90})
            begin
              reg107 <= wire103;
              reg108 <= reg92[(2'h3):(1'h0)];
              reg109 <= reg86[(2'h2):(1'h1)];
            end
          else
            begin
              reg107 <= reg94;
              reg108 <= {(wire103 ^ (reg76 ? (|wire9) : reg105)),
                  $signed((~$signed({wire11})))};
              reg109 <= {(8'hb6)};
              reg110 <= reg84;
              reg111 <= $signed(((~^{(+reg101), {wire103, (8'hbb)}}) ?
                  {reg85} : (~reg78)));
            end
          if ({{((reg81 ^ (reg77 | reg91)) ?
                      $signed(wire103[(5'h11):(2'h3)]) : ({reg99} ?
                          (reg91 ? reg94 : wire103) : (reg106 > reg83))),
                  $signed(($signed(reg88) + {(8'h9c), reg110}))}})
            begin
              reg112 <= wire11;
              reg113 <= reg101;
            end
          else
            begin
              reg112 <= $unsigned({$signed(($unsigned(reg83) == (~^reg91)))});
            end
          if ((wire72 >>> $signed({((reg78 << reg96) == {(8'ha0), reg86})})))
            begin
              reg114 <= ((~|(8'hab)) ?
                  reg105[(4'hb):(3'h4)] : (reg92 >> reg100[(1'h0):(1'h0)]));
              reg115 <= (reg79 - $signed((reg111[(2'h2):(1'h1)] ?
                  ($unsigned(reg99) == $unsigned((8'hac))) : reg80[(1'h0):(1'h0)])));
              reg116 <= {$signed(({wire103[(4'h8):(1'h0)]} ^~ $signed(reg90))),
                  ($signed({reg84}) ?
                      ($signed((reg98 ^~ reg85)) - ($signed(reg85) ?
                          (^~reg76) : $unsigned(reg109))) : (8'hb3))};
            end
          else
            begin
              reg114 <= reg116[(3'h6):(1'h1)];
            end
          reg117 <= reg76[(2'h3):(1'h1)];
          reg118 <= (reg99 ?
              reg106 : ({reg91[(1'h0):(1'h0)]} ?
                  {$unsigned((reg95 ? reg92 : reg76))} : (($signed(reg107) ?
                          reg104 : {reg100, (8'hb6)}) ?
                      ((reg115 >>> reg74) > (reg92 ?
                          reg107 : (7'h42))) : reg115)));
        end
      else
        begin
          reg107 <= ($signed($signed((~&$signed(wire103)))) ?
              ((~|(^~(reg87 ^ reg92))) * $unsigned(reg92)) : (~&$unsigned($unsigned((!reg118)))));
          reg108 <= reg102[(4'hc):(2'h3)];
        end
      reg119 <= (reg95 ?
          $unsigned(reg97[(1'h1):(1'h1)]) : {reg83[(4'h8):(3'h6)],
              (+$signed($unsigned(reg80)))});
      reg120 <= (reg116[(3'h4):(3'h4)] * ($unsigned(reg104) ?
          (8'hb5) : reg89[(5'h12):(4'hf)]));
    end
  always
    @(posedge clk) begin
      if (($unsigned((8'hba)) ?
          ((reg82[(3'h7):(3'h4)] ?
              reg108[(1'h1):(1'h1)] : reg94[(5'h10):(3'h7)]) >= ($unsigned($signed(reg120)) <= reg112[(5'h11):(2'h3)])) : reg95[(3'h5):(2'h2)]))
        begin
          if (reg119)
            begin
              reg121 <= $signed(reg74[(1'h0):(1'h0)]);
              reg122 <= ($signed({reg81}) ?
                  reg112[(4'ha):(3'h5)] : reg101[(2'h2):(2'h2)]);
              reg123 <= (reg120 ?
                  ({(reg121[(4'he):(2'h3)] ^~ $unsigned(reg116)),
                          $unsigned((|reg106))} ?
                      wire9[(4'he):(4'h9)] : reg83) : (~|$signed({(~^reg107),
                      $unsigned((8'hae))})));
              reg124 <= {{(reg111 < {(wire11 ? reg82 : reg102)}),
                      $unsigned($unsigned($unsigned(wire103)))}};
            end
          else
            begin
              reg121 <= reg94;
              reg122 <= (((~|(^~{(8'h9e), reg80})) ?
                  ($unsigned(wire72[(1'h1):(1'h0)]) == ((!wire6) >>> $signed(reg94))) : $signed((((8'hb5) << reg81) ?
                      (reg74 != reg99) : (|reg95)))) * wire12);
            end
          reg125 <= reg120;
          reg126 <= (({$signed(reg110[(4'h8):(1'h1)])} ?
                  $unsigned($unsigned((8'ha8))) : (($signed(wire8) ?
                          $unsigned(reg106) : $signed(reg111)) ?
                      {$unsigned(reg122)} : reg99)) ?
              reg111 : ((^(reg91[(2'h2):(2'h2)] ? (~reg80) : reg121)) ?
                  wire7[(1'h0):(1'h0)] : reg82));
          reg127 <= reg80[(4'hd):(1'h1)];
        end
      else
        begin
          reg121 <= (($signed((((7'h41) != reg122) ?
                  reg96[(3'h4):(2'h2)] : $unsigned(reg101))) ?
              {reg89} : (reg97 >> reg75[(3'h4):(1'h0)])) <<< (!$unsigned(((wire8 || reg76) ?
              (reg81 ? reg117 : reg111) : (reg109 == (8'h9c))))));
        end
      reg128 <= (~$signed(reg90));
      reg129 <= {wire72[(5'h12):(4'hc)]};
      if ($unsigned((8'hab)))
        begin
          reg130 <= {(8'h9c),
              {reg118,
                  $unsigned(((~reg97) ?
                      $unsigned(reg129) : (reg82 ? reg77 : (8'h9f))))}};
          reg131 <= $signed($unsigned(reg78));
        end
      else
        begin
          reg130 <= (~^(($signed((~^reg125)) ?
              reg123[(1'h0):(1'h0)] : reg74[(2'h2):(2'h2)]) ~^ reg97[(2'h3):(1'h1)]));
          reg131 <= (reg87[(1'h0):(1'h0)] != (~&(((reg100 | reg89) ?
              (reg111 || (8'haf)) : $unsigned(reg130)) == $unsigned(reg92[(2'h2):(1'h0)]))));
          reg132 <= reg100[(2'h2):(1'h1)];
        end
      reg133 <= $signed((~&reg131[(3'h6):(3'h6)]));
    end
  assign wire134 = ({reg112, reg79} & $signed($unsigned(reg121)));
  assign wire135 = reg85;
  always
    @(posedge clk) begin
      reg136 <= (&reg126);
      if ($signed((($unsigned($signed(wire6)) ?
              $signed({reg114}) : (~^(reg88 << reg99))) ?
          reg115 : (reg118[(2'h3):(2'h2)] ?
              $unsigned((reg121 >= (8'h9e))) : reg74[(1'h1):(1'h0)]))))
        begin
          if ($signed(reg78[(4'ha):(3'h4)]))
            begin
              reg137 <= {reg131[(2'h2):(2'h2)]};
              reg138 <= $unsigned(($unsigned(((reg81 ^ reg128) << $unsigned(reg98))) ?
                  ({reg119[(2'h2):(2'h2)], (reg74 ? reg115 : wire134)} ?
                      ((+reg129) >> {reg85,
                          wire7}) : $unsigned((reg128 ^ (8'ha4)))) : reg101));
              reg139 <= ($signed({reg86[(2'h2):(2'h2)]}) ?
                  ((&(reg104 + (+reg80))) * (~&$unsigned((~&reg79)))) : ((wire72 != (wire134 ?
                      reg114 : (wire9 ?
                          reg126 : reg114))) - (reg124 >> $unsigned((~^reg99)))));
            end
          else
            begin
              reg137 <= $signed((&reg100[(2'h3):(2'h3)]));
              reg138 <= {$unsigned($signed(reg139))};
              reg139 <= $unsigned(reg84);
              reg140 <= ($signed(reg120[(4'h9):(3'h7)]) ?
                  $unsigned({(8'hb9),
                      reg88}) : ((~|reg112[(3'h4):(2'h2)]) << (reg139[(2'h3):(1'h1)] == $signed((wire135 ?
                      (8'hb2) : reg84)))));
            end
        end
      else
        begin
          reg137 <= wire8[(4'h8):(3'h4)];
          reg138 <= ($unsigned(reg130) ?
              {((^~(reg113 ? reg74 : reg123)) ?
                      (+$unsigned(reg131)) : $unsigned($unsigned((8'hb1))))} : $unsigned((8'h9d)));
        end
      if (reg120[(3'h5):(2'h3)])
        begin
          reg141 <= ($signed((reg82 ?
              (-reg140[(3'h4):(1'h0)]) : {reg125,
                  reg126[(2'h2):(2'h2)]})) < (reg108 ^ (wire103 <<< (~&reg124))));
          reg142 <= ({{$signed(reg91[(1'h1):(1'h0)]),
                      ((reg112 && reg90) ? (reg113 == (8'hb3)) : {reg102})},
                  {((reg131 ? reg92 : reg129) >> (^reg118)),
                      $signed((~&reg75))}} ?
              reg89[(5'h10):(5'h10)] : (reg79 << reg80[(2'h2):(2'h2)]));
          reg143 <= ((reg113[(3'h4):(2'h2)] + $signed(reg98)) ?
              (&(-(!(wire103 << reg102)))) : $unsigned($signed(reg107)));
          reg144 <= ((reg105[(3'h4):(3'h4)] ?
                  ({(reg101 ? reg99 : reg90),
                      (reg114 ~^ reg131)} > $unsigned($signed(reg88))) : {(8'hb9),
                      reg137[(1'h0):(1'h0)]}) ?
              ((wire9 ? $unsigned($signed(reg123)) : reg101) < (wire134 ?
                  wire9 : $unsigned(wire72))) : (8'hb6));
        end
      else
        begin
          reg141 <= {(^reg142), ({(!reg123)} <= reg126)};
          if (reg94[(4'h8):(3'h5)])
            begin
              reg142 <= (~|(reg120 || $unsigned(((7'h43) || (reg75 ?
                  wire11 : reg92)))));
            end
          else
            begin
              reg142 <= $signed(reg116[(3'h6):(2'h2)]);
              reg143 <= (reg93 ?
                  $unsigned(($signed(reg112[(4'hc):(1'h1)]) != ((reg124 ?
                      reg91 : reg115) | (8'hbc)))) : reg102);
            end
          if ((8'h9f))
            begin
              reg144 <= ((+(reg93 != $signed((wire7 <= reg129)))) ?
                  $unsigned(($unsigned($unsigned(reg108)) ^ $unsigned((wire8 ?
                      reg89 : (8'hb8))))) : $unsigned((~($signed(reg121) ?
                      (8'ha3) : (+reg86)))));
              reg145 <= ($unsigned(reg112[(3'h4):(2'h2)]) >>> $unsigned(reg115));
              reg146 <= (~(wire7[(2'h2):(2'h2)] ?
                  reg137[(3'h4):(2'h3)] : $unsigned((8'h9f))));
              reg147 <= reg99;
              reg148 <= $signed(reg132[(1'h1):(1'h0)]);
            end
          else
            begin
              reg144 <= (^$signed(reg143));
              reg145 <= reg121;
            end
          reg149 <= reg99[(4'h9):(1'h0)];
          reg150 <= $signed((($signed($unsigned(reg101)) >= $unsigned($unsigned(reg94))) >>> reg127[(4'hb):(4'ha)]));
        end
      reg151 <= $signed((~$unsigned(($unsigned(reg118) ?
          $signed((8'had)) : (reg127 < reg136)))));
    end
  assign wire152 = reg95[(1'h0):(1'h0)];
  module153_1 #() modinst169 (.clk(clk), .wire157(wire11), .wire155(reg76), .wire156(reg117), .y(wire168), .wire158(reg112), .wire154(reg121));
  assign wire170 = reg129[(5'h12):(3'h6)];
endmodule

module module153_1  (y, clk, wire158, wire157, wire156, wire155, wire154);
  output wire [(32'h6c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire158;
  input wire signed [(4'hc):(1'h0)] wire157;
  input wire [(3'h5):(1'h0)] wire156;
  input wire [(3'h4):(1'h0)] wire155;
  input wire signed [(5'h12):(1'h0)] wire154;
  wire [(2'h3):(1'h0)] wire167;
  wire signed [(5'h14):(1'h0)] wire166;
  wire signed [(3'h7):(1'h0)] wire165;
  wire [(5'h13):(1'h0)] wire164;
  wire signed [(5'h10):(1'h0)] wire163;
  wire [(4'he):(1'h0)] wire162;
  wire [(3'h4):(1'h0)] wire161;
  reg [(3'h6):(1'h0)] reg160 = (1'h0);
  reg [(5'h12):(1'h0)] reg159 = (1'h0);
  assign y = {wire167,
                 wire166,
                 wire165,
                 wire164,
                 wire163,
                 wire162,
                 wire161,
                 reg160,
                 reg159,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg159 <= wire158[(3'h5):(1'h0)];
      reg160 <= $unsigned((&(reg159 ~^ $signed($signed(reg159)))));
    end
  assign wire161 = wire156;
  assign wire162 = $signed(wire155[(2'h2):(2'h2)]);
  assign wire163 = $signed($unsigned($unsigned(((reg160 - (8'h9c)) == wire158[(3'h6):(3'h4)]))));
  assign wire164 = ({$unsigned({$signed(wire157)})} ?
                       (((wire157[(1'h0):(1'h0)] ?
                               (wire161 ? wire157 : (7'h44)) : (reg160 ?
                                   wire163 : wire154)) <<< $unsigned({wire161})) ?
                           ($signed($unsigned(wire157)) - reg160[(1'h1):(1'h0)]) : wire154[(5'h11):(3'h7)]) : wire156);
  assign wire165 = wire162[(1'h0):(1'h0)];
  assign wire166 = wire165[(1'h1):(1'h0)];
  assign wire167 = reg159;
endmodule

module module13_1
#(parameter param71 = (^(-({((8'hb6) ? (8'hb6) : (8'hba)), ((8'hb9) >>> (8'had))} ? ({(8'hae), (8'hb8)} ? ((8'ha9) ? (8'hb8) : (7'h42)) : ((8'hba) >> (7'h40))) : ((8'hbb) >>> {(8'hb5), (8'hb9)})))))
(y, clk, wire18, wire17, wire16, wire15, wire14);
  output wire [(32'h23e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire18;
  input wire signed [(4'he):(1'h0)] wire17;
  input wire signed [(5'h14):(1'h0)] wire16;
  input wire signed [(4'hd):(1'h0)] wire15;
  input wire [(2'h2):(1'h0)] wire14;
  wire signed [(5'h12):(1'h0)] wire65;
  wire signed [(4'ha):(1'h0)] wire44;
  wire signed [(5'h11):(1'h0)] wire35;
  wire signed [(4'hd):(1'h0)] wire34;
  wire [(3'h7):(1'h0)] wire33;
  wire [(4'he):(1'h0)] wire32;
  wire [(3'h4):(1'h0)] wire31;
  wire [(4'hc):(1'h0)] wire30;
  wire signed [(4'h9):(1'h0)] wire29;
  wire [(4'hc):(1'h0)] wire28;
  wire [(2'h2):(1'h0)] wire27;
  wire signed [(5'h13):(1'h0)] wire26;
  wire signed [(3'h6):(1'h0)] wire25;
  wire [(4'h9):(1'h0)] wire24;
  wire signed [(5'h15):(1'h0)] wire23;
  wire [(3'h5):(1'h0)] wire22;
  wire [(3'h4):(1'h0)] wire21;
  wire signed [(4'h9):(1'h0)] wire20;
  wire signed [(4'hf):(1'h0)] wire19;
  reg signed [(5'h11):(1'h0)] reg70 = (1'h0);
  reg [(2'h2):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg68 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg66 = (1'h0);
  reg [(4'hd):(1'h0)] reg64 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg63 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg62 = (1'h0);
  reg [(5'h15):(1'h0)] reg61 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg60 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg59 = (1'h0);
  reg [(4'he):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg56 = (1'h0);
  reg [(4'ha):(1'h0)] reg55 = (1'h0);
  reg [(3'h7):(1'h0)] reg54 = (1'h0);
  reg [(5'h15):(1'h0)] reg53 = (1'h0);
  reg [(4'he):(1'h0)] reg52 = (1'h0);
  reg [(2'h3):(1'h0)] reg51 = (1'h0);
  reg [(4'hc):(1'h0)] reg50 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg49 = (1'h0);
  reg [(5'h12):(1'h0)] reg48 = (1'h0);
  reg [(4'hc):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg46 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg45 = (1'h0);
  reg [(3'h5):(1'h0)] reg43 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg42 = (1'h0);
  reg [(3'h7):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg39 = (1'h0);
  reg [(3'h4):(1'h0)] reg38 = (1'h0);
  reg [(5'h12):(1'h0)] reg37 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg36 = (1'h0);
  assign y = {wire65,
                 wire44,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 wire31,
                 wire30,
                 wire29,
                 wire28,
                 wire27,
                 wire26,
                 wire25,
                 wire24,
                 wire23,
                 wire22,
                 wire21,
                 wire20,
                 wire19,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 (1'h0)};
  assign wire19 = (|$signed(wire18));
  assign wire20 = $unsigned(wire18[(2'h2):(1'h1)]);
  assign wire21 = $signed($signed(wire20[(1'h0):(1'h0)]));
  assign wire22 = $signed((wire18 ?
                      (((8'hbd) ?
                          $signed(wire18) : $signed(wire16)) * {(wire16 ?
                              wire21 : wire17)}) : $unsigned({wire18,
                          (wire19 ? wire18 : wire16)})));
  assign wire23 = wire18[(2'h2):(1'h0)];
  assign wire24 = ($unsigned(($signed($unsigned((8'ha9))) ?
                      $signed({wire21,
                          wire20}) : wire15[(4'h9):(2'h3)])) <<< $signed($unsigned($signed(wire20))));
  assign wire25 = ($unsigned(wire21) ^~ wire15);
  assign wire26 = $unsigned($signed(({(wire19 >= wire21),
                      $signed(wire16)} << (~|$signed(wire15)))));
  assign wire27 = wire23[(4'hd):(3'h7)];
  assign wire28 = $unsigned((~|$signed(wire14[(2'h2):(2'h2)])));
  assign wire29 = (7'h44);
  assign wire30 = (wire18[(2'h2):(2'h2)] ~^ wire14);
  assign wire31 = {(wire25[(3'h4):(1'h0)] - {{(wire29 || (8'ha9)),
                              (wire22 ? (7'h42) : wire26)},
                          ($unsigned(wire16) <<< wire24)})};
  assign wire32 = {wire30[(4'hb):(4'hb)], $signed(wire31)};
  assign wire33 = wire21;
  assign wire34 = $unsigned($signed({((~&wire25) ?
                          $signed(wire30) : (wire27 << wire20)),
                      $signed(wire25[(3'h6):(1'h0)])}));
  assign wire35 = {wire22,
                      $unsigned(((!$unsigned((8'had))) ?
                          (^$signed((8'hb2))) : {(~|wire31)}))};
  always
    @(posedge clk) begin
      reg36 <= {(+(wire27 & $unsigned($unsigned(wire33))))};
      if ($unsigned((wire22 ?
          $signed(({(8'hbd), wire30} <<< wire14)) : wire26)))
        begin
          reg37 <= wire21;
        end
      else
        begin
          reg37 <= (wire28[(3'h6):(2'h3)] | (((|(+wire26)) ?
              (wire21 ?
                  wire30[(3'h5):(3'h4)] : (wire31 >> (8'hb7))) : (^~{wire29,
                  (8'ha1)})) <<< {$unsigned({wire17, wire30})}));
          reg38 <= (({$unsigned((^~wire16))} && (!{wire29[(1'h0):(1'h0)]})) + wire27[(1'h1):(1'h0)]);
          reg39 <= $unsigned($unsigned(({((8'ha1) ? reg37 : wire35),
              $signed(wire23)} == (8'ha3))));
          reg40 <= $signed($signed((+wire30[(4'hc):(2'h3)])));
          reg41 <= (8'hb3);
        end
      reg42 <= ($signed((!(wire25 >= wire22[(2'h3):(2'h2)]))) ?
          ((wire20 == wire24[(4'h9):(3'h5)]) >>> reg39[(1'h1):(1'h1)]) : $unsigned(wire16[(3'h5):(2'h3)]));
      reg43 <= ($unsigned($signed((wire24[(3'h5):(1'h1)] ? wire24 : wire32))) ?
          $unsigned((wire18 ?
              (wire27 ? (wire33 != wire15) : $unsigned(wire31)) : {{reg42,
                      reg39}})) : ($signed(((reg38 ?
                  reg36 : wire18) < wire30)) ?
              ($signed((reg39 ?
                  wire26 : wire32)) >= $unsigned($signed(wire27))) : (({wire24,
                      reg37} != (wire23 * (7'h40))) ?
                  ((wire34 ? wire32 : wire32) ?
                      (~^reg37) : $unsigned(reg39)) : wire33[(1'h1):(1'h0)])));
    end
  assign wire44 = (!$unsigned($signed(({wire23} != (wire19 ?
                      wire34 : reg38)))));
  always
    @(posedge clk) begin
      if (wire16[(4'ha):(3'h6)])
        begin
          if ((^{$signed((!(!wire33)))}))
            begin
              reg45 <= (~(((^(8'hac)) < {(reg38 < wire31)}) || (($signed(wire18) ?
                      wire16 : {reg40}) ?
                  wire29[(3'h5):(3'h4)] : $unsigned(((8'hb7) ?
                      (8'haa) : (8'hbb))))));
              reg46 <= ((wire14 ?
                  {(+((8'hbc) - (8'ha2))),
                      ((|(8'hbf)) - {reg36})} : ($signed((!wire30)) ?
                      wire34[(1'h0):(1'h0)] : reg37[(2'h3):(1'h0)])) >>> reg39[(3'h6):(3'h6)]);
            end
          else
            begin
              reg45 <= $signed((wire19 ? (8'hbb) : reg46[(3'h4):(2'h3)]));
              reg46 <= wire24;
            end
          if ((($signed(((~reg36) >>> wire31)) - $unsigned((^$unsigned(wire16)))) ?
              wire20 : $unsigned({(wire25[(2'h3):(2'h3)] + reg46[(1'h0):(1'h0)])})))
            begin
              reg47 <= (wire19 | (^(((wire20 | wire31) ?
                  {(8'ha4)} : $signed(reg43)) <<< wire19[(4'ha):(1'h0)])));
              reg48 <= $signed(wire16[(2'h2):(1'h1)]);
            end
          else
            begin
              reg47 <= {$unsigned($unsigned(($unsigned(wire27) <= $unsigned(reg36)))),
                  $unsigned((wire32 ?
                      $unsigned((wire17 ? wire22 : (8'hbb))) : (-(~^wire21))))};
              reg48 <= $unsigned($signed(wire21));
              reg49 <= (&wire28[(1'h1):(1'h1)]);
            end
        end
      else
        begin
          reg45 <= $signed($signed({$unsigned(((7'h40) - wire28))}));
          if ($signed($unsigned(($unsigned($unsigned(reg40)) ?
              reg48 : $signed((-(8'ha0)))))))
            begin
              reg46 <= wire22[(2'h2):(2'h2)];
              reg47 <= $signed({(({wire15} ?
                      (8'hb5) : reg43[(3'h4):(2'h3)]) << reg37)});
              reg48 <= ($signed({($signed(wire26) ?
                          (reg41 >> (8'hb4)) : $unsigned(wire19)),
                      $unsigned((!reg43))}) ?
                  (wire23[(3'h5):(3'h5)] ?
                      $signed((^~(+wire29))) : {$unsigned({reg38, wire19}),
                          $unsigned($unsigned(wire24))}) : wire14[(1'h1):(1'h1)]);
              reg49 <= $unsigned((wire26 > (((&wire34) <= reg46) | {$signed(reg47),
                  wire28[(4'h8):(3'h7)]})));
              reg50 <= ($signed({$unsigned((wire21 | wire23)), wire30}) ?
                  reg45 : $signed($unsigned(wire16)));
            end
          else
            begin
              reg46 <= (+$unsigned(reg46));
              reg47 <= (reg42[(2'h2):(2'h2)] ?
                  $unsigned((~|(wire35 || reg45[(1'h1):(1'h1)]))) : ((wire32[(4'he):(2'h3)] <<< (wire16 ?
                          wire27[(1'h0):(1'h0)] : (wire28 <<< reg45))) ?
                      {$unsigned((reg42 ^~ wire33)),
                          $signed((+(8'hab)))} : $unsigned({(~^reg37),
                          $signed(wire17)})));
            end
          reg51 <= wire35[(4'hd):(1'h0)];
          reg52 <= $unsigned($unsigned(reg37[(4'hd):(2'h3)]));
          if ((7'h40))
            begin
              reg53 <= ($signed(((8'hac) ?
                      (wire24 ?
                          (reg36 ?
                              reg36 : wire22) : (wire20 != reg40)) : {(reg42 & wire17),
                          (&wire28)})) ?
                  wire24[(2'h2):(1'h1)] : reg51[(1'h1):(1'h0)]);
              reg54 <= (8'hb4);
              reg55 <= reg38;
              reg56 <= $unsigned((!$unsigned(wire16)));
            end
          else
            begin
              reg53 <= wire35[(4'ha):(4'ha)];
              reg54 <= (($signed({$unsigned(reg48),
                  $unsigned(reg50)}) < $unsigned((~|reg36[(4'h8):(4'h8)]))) >= ({$signed(wire44),
                      $signed(((8'hb0) > wire19))} ?
                  $unsigned((wire32 ?
                      (wire26 ?
                          reg55 : wire17) : $unsigned(reg46))) : $unsigned(((reg51 >>> reg37) ?
                      reg46[(2'h3):(1'h0)] : (^reg36)))));
              reg55 <= ($unsigned((~&reg54[(2'h2):(1'h1)])) != (~&(wire30 ?
                  $signed(reg49) : (~$signed(wire35)))));
            end
        end
      if (((~&((!(~&reg36)) ? (wire35 * $unsigned(reg37)) : $signed(reg54))) ?
          reg49 : wire28[(1'h0):(1'h0)]))
        begin
          reg57 <= ((|(((8'hbb) ?
                  $unsigned((8'hbd)) : $unsigned((8'hb2))) <<< ((reg45 ?
                  reg48 : wire21) << $signed(reg41)))) ?
              $unsigned((($signed(wire29) != wire34) ?
                  ((8'ha1) ?
                      (+wire35) : $unsigned(wire25)) : $unsigned($signed(reg53)))) : $signed(wire30[(3'h7):(3'h4)]));
        end
      else
        begin
          reg57 <= wire19;
          if ((^~$unsigned(reg38)))
            begin
              reg58 <= wire29[(3'h5):(1'h1)];
              reg59 <= ((^~wire25[(1'h1):(1'h0)]) ^~ ((|wire29) ?
                  $unsigned({$signed(wire20)}) : $unsigned($unsigned((wire16 ?
                      wire27 : reg50)))));
              reg60 <= {reg55, wire19[(4'hb):(1'h0)]};
              reg61 <= $signed({$signed(($signed(wire35) && (wire25 ?
                      reg58 : reg50))),
                  $unsigned(wire27)});
              reg62 <= wire22;
            end
          else
            begin
              reg58 <= (|wire31[(2'h3):(1'h0)]);
              reg59 <= ((&($signed($unsigned(reg42)) ?
                  ((reg51 ? reg54 : wire25) & reg39) : (reg39[(4'hb):(3'h7)] ?
                      reg38[(1'h0):(1'h0)] : $signed(wire23)))) < $signed($signed(($unsigned(wire23) ?
                  wire22 : $unsigned(reg55)))));
              reg60 <= wire35[(2'h2):(1'h1)];
              reg61 <= reg51[(2'h2):(1'h1)];
            end
        end
      reg63 <= reg54[(2'h2):(1'h1)];
      reg64 <= (+$unsigned($unsigned(wire14[(1'h1):(1'h1)])));
    end
  assign wire65 = reg41;
  always
    @(posedge clk) begin
      reg66 <= {$signed($unsigned({$signed(reg49), wire17}))};
      if ((((-{(7'h41)}) ?
          $signed($signed((wire23 <<< reg38))) : (($unsigned(reg64) ?
              wire18 : (~wire23)) ~^ (wire65 ?
              (wire20 ?
                  reg39 : wire14) : $signed(reg59)))) | reg52[(4'ha):(3'h5)]))
        begin
          reg67 <= {$signed((^($signed(wire23) ?
                  wire19 : reg62[(3'h7):(3'h4)]))),
              ((reg62 ?
                  wire16[(5'h10):(3'h7)] : $signed((wire65 | reg61))) > ((wire19[(3'h6):(3'h4)] + $unsigned(wire17)) != (~|wire20[(2'h2):(2'h2)])))};
          reg68 <= (^$signed(($signed($signed((8'hb4))) ?
              (|wire26[(4'h8):(4'h8)]) : reg67[(1'h0):(1'h0)])));
          reg69 <= (~^{reg66[(1'h0):(1'h0)]});
          if ($signed({($unsigned((reg56 == (8'ha6))) || $unsigned((^~reg55)))}))
            begin
              reg70 <= wire24;
            end
          else
            begin
              reg70 <= $unsigned($unsigned((|reg61)));
            end
        end
      else
        begin
          reg67 <= (~|$signed(wire30));
          if ((reg48[(4'hf):(4'ha)] ?
              (reg63 > wire33) : (({reg36[(2'h3):(2'h2)]} ?
                  (^reg69[(2'h2):(2'h2)]) : reg55[(4'h9):(1'h0)]) >> $unsigned(reg47))))
            begin
              reg68 <= ($signed(reg38[(3'h4):(2'h3)]) != ((+((&reg62) || $signed(wire15))) ?
                  (~|$unsigned(wire26)) : (~|reg49)));
              reg69 <= (8'h9e);
            end
          else
            begin
              reg68 <= reg69;
            end
          reg70 <= reg42[(2'h3):(2'h3)];
        end
    end
endmodule

module module278_1
#(parameter param329 = (~|{(&((-(8'hb0)) ? ((7'h40) ? (8'hab) : (8'h9d)) : {(7'h43), (8'h9f)}))}), 
parameter param330 = {((+(7'h43)) & ({{param329}, (^~(8'had))} >>> ((|param329) ^ {param329, param329})))})
(y, clk, wire283, wire282, wire281, wire280, wire279);
  output wire [(32'h1f4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire283;
  input wire [(4'hc):(1'h0)] wire282;
  input wire signed [(4'he):(1'h0)] wire281;
  input wire [(3'h6):(1'h0)] wire280;
  input wire signed [(5'h12):(1'h0)] wire279;
  wire [(4'ha):(1'h0)] wire324;
  wire [(4'h8):(1'h0)] wire312;
  wire [(4'hb):(1'h0)] wire311;
  wire signed [(5'h10):(1'h0)] wire307;
  wire [(4'h8):(1'h0)] wire306;
  wire [(5'h10):(1'h0)] wire305;
  wire signed [(4'hc):(1'h0)] wire304;
  wire signed [(4'h9):(1'h0)] wire296;
  wire [(3'h6):(1'h0)] wire284;
  reg signed [(5'h12):(1'h0)] reg328 = (1'h0);
  reg [(4'ha):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg326 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg325 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg323 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg321 = (1'h0);
  reg [(4'he):(1'h0)] reg320 = (1'h0);
  reg [(5'h10):(1'h0)] reg319 = (1'h0);
  reg [(2'h3):(1'h0)] reg318 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg317 = (1'h0);
  reg [(5'h12):(1'h0)] reg316 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg315 = (1'h0);
  reg [(3'h4):(1'h0)] reg314 = (1'h0);
  reg [(4'h9):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg310 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg309 = (1'h0);
  reg [(5'h13):(1'h0)] reg308 = (1'h0);
  reg [(5'h14):(1'h0)] reg303 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg302 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg301 = (1'h0);
  reg [(4'hd):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg299 = (1'h0);
  reg [(4'h9):(1'h0)] reg298 = (1'h0);
  reg [(5'h10):(1'h0)] reg297 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg295 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg294 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg293 = (1'h0);
  reg signed [(4'he):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg291 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg290 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg288 = (1'h0);
  reg [(5'h15):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg286 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg285 = (1'h0);
  assign y = {wire324,
                 wire312,
                 wire311,
                 wire307,
                 wire306,
                 wire305,
                 wire304,
                 wire296,
                 wire284,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg310,
                 reg309,
                 reg308,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 (1'h0)};
  assign wire284 = wire279[(3'h4):(3'h4)];
  always
    @(posedge clk) begin
      reg285 <= $unsigned($signed(((8'ha7) ?
          {$unsigned(wire281)} : wire281[(4'he):(3'h7)])));
      reg286 <= (wire281[(1'h1):(1'h0)] < {(wire281[(2'h2):(1'h0)] ?
              ($unsigned(reg285) ?
                  wire284[(3'h4):(1'h1)] : wire284) : $unsigned(((8'ha3) != (8'ha2)))),
          {{(~&wire282), {wire283, wire283}},
              (wire283 ? wire279 : (~wire284))}});
    end
  always
    @(posedge clk) begin
      reg287 <= {(((&(wire281 ? reg286 : wire284)) ?
              reg286[(4'hd):(4'ha)] : $signed($unsigned(wire284))) * $unsigned(reg285[(2'h2):(1'h0)])),
          wire281};
      reg288 <= $unsigned(((~|(reg285[(2'h3):(1'h0)] ?
          {wire283, wire280} : reg286[(5'h10):(1'h1)])) ^~ wire283));
      if ($signed((7'h44)))
        begin
          reg289 <= wire280;
          reg290 <= ($signed($unsigned({((8'haa) ?
                  wire280 : wire284)})) < ($unsigned(reg289) ?
              wire279 : (~&(!$signed(reg286)))));
          reg291 <= reg286;
          reg292 <= reg287[(4'hd):(4'h9)];
          reg293 <= ($unsigned(reg286) ?
              $unsigned(({(|wire279), $signed(wire284)} ^ ((~&wire280) ?
                  $unsigned(wire284) : $unsigned(reg290)))) : reg288);
        end
      else
        begin
          if ({$signed(($signed((reg288 ? reg291 : reg285)) ^ ({reg292} ?
                  $unsigned(wire280) : (reg285 ? reg293 : reg287)))),
              (((~&(-reg291)) ?
                  {$unsigned(reg286),
                      reg292} : {$signed((8'ha0))}) & $unsigned(reg287[(2'h2):(1'h0)]))})
            begin
              reg289 <= $signed(reg288);
              reg290 <= (^($signed(reg288[(4'h9):(2'h2)]) < (($unsigned(wire284) >> $unsigned(reg287)) ~^ reg293)));
            end
          else
            begin
              reg289 <= reg287[(5'h12):(4'hb)];
              reg290 <= {wire284,
                  ((&reg287) != $unsigned(($unsigned(reg289) * {reg289})))};
            end
          reg291 <= $signed(((8'hb8) & $signed(((wire283 ?
              wire282 : reg290) && reg285))));
          reg292 <= ((!wire282) ?
              ({$signed({reg291,
                      (7'h41)})} ~^ wire279[(4'hf):(3'h4)]) : (reg286 ?
                  $unsigned((8'ha4)) : $signed($unsigned({reg292}))));
          if (((wire280[(3'h4):(1'h1)] < (reg288 ?
                  $unsigned($unsigned(reg289)) : ((-wire281) ?
                      ((8'h9f) ? reg289 : reg292) : (~&wire282)))) ?
              (-(~^((~&wire279) != $unsigned(reg292)))) : (8'hb9)))
            begin
              reg293 <= ((reg290 ?
                  ($unsigned((~wire281)) || ({(7'h43)} | (wire283 ?
                      reg290 : reg291))) : ((~|(!(8'ha2))) ?
                      (((8'ha1) ?
                          wire284 : (8'ha8)) >> (reg289 <= reg290)) : ($unsigned(wire281) ?
                          {reg287,
                              reg286} : (reg285 >>> (8'hb5))))) - $signed((wire282[(2'h2):(1'h1)] | {{reg291},
                  $signed((8'h9c))})));
            end
          else
            begin
              reg293 <= reg286[(4'hf):(4'he)];
            end
        end
      reg294 <= {{(^~$unsigned({(7'h41)}))}};
      reg295 <= $unsigned((wire280 & ((wire279 ?
              (wire281 << wire283) : ((8'had) ? wire280 : reg286)) ?
          ({(8'hb5)} ? reg294 : (+reg294)) : (|reg286))));
    end
  assign wire296 = wire283[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg297 <= {{(~&reg286[(1'h1):(1'h1)]), (8'ha4)}};
      reg298 <= (^$signed(wire281[(4'h9):(3'h5)]));
      if ($unsigned(reg286))
        begin
          reg299 <= wire284[(3'h4):(2'h3)];
          reg300 <= wire284[(1'h0):(1'h0)];
          reg301 <= ((reg300[(3'h4):(1'h1)] ?
                  $signed(((~^wire279) <= reg297[(5'h10):(3'h6)])) : (~^(reg297 <<< reg286))) ?
              {((^(reg289 << wire284)) <<< $signed((!wire284)))} : (wire284[(2'h2):(1'h1)] < (-((^reg295) || reg291[(3'h7):(2'h2)]))));
        end
      else
        begin
          reg299 <= reg299[(1'h0):(1'h0)];
          reg300 <= reg297[(2'h2):(2'h2)];
          if ({(~reg301[(1'h1):(1'h1)])})
            begin
              reg301 <= ($signed((&{(reg294 ?
                      (8'h9d) : wire280)})) > $signed(({$unsigned(wire279)} >>> ((~wire279) ?
                  reg299 : ((7'h42) ? reg299 : wire283)))));
              reg302 <= (~^wire283);
              reg303 <= $unsigned($unsigned($signed({$unsigned(reg298)})));
            end
          else
            begin
              reg301 <= $unsigned($signed((((reg293 ? reg288 : reg300) ?
                      wire280 : (reg299 * reg300)) ?
                  ((~reg290) ?
                      $unsigned(wire280) : (wire284 ?
                          reg297 : reg299)) : (reg288 ?
                      $unsigned(reg295) : (^~reg295)))));
            end
        end
    end
  assign wire304 = $unsigned($signed($signed($signed($unsigned((8'haf))))));
  assign wire305 = (~&$unsigned({(reg301 ?
                           {reg287, wire280} : {reg299, reg300})}));
  assign wire306 = ((~$unsigned((^reg292))) ?
                       ($signed($signed(wire283[(1'h1):(1'h0)])) << ((&{(8'ha5)}) ?
                           $unsigned((reg297 ?
                               reg285 : (8'h9d))) : (8'hb1))) : reg292[(1'h0):(1'h0)]);
  assign wire307 = (8'hb7);
  always
    @(posedge clk) begin
      reg308 <= {(reg302 & $signed(((reg303 ? reg288 : reg303) ?
              {reg297} : $unsigned(reg288))))};
      reg309 <= (^reg302);
      reg310 <= wire283[(1'h0):(1'h0)];
    end
  assign wire311 = ({$unsigned($signed($unsigned(reg297)))} ?
                       {(&reg286)} : $unsigned({wire307[(4'hd):(4'ha)]}));
  assign wire312 = $unsigned($signed(wire305[(4'hc):(3'h7)]));
  always
    @(posedge clk) begin
      reg313 <= (((wire296[(3'h4):(1'h0)] * ((!reg301) ?
              reg298 : $signed(reg297))) ?
          reg290[(3'h4):(1'h1)] : reg309[(2'h2):(1'h0)]) ^ ((|$signed((reg301 ?
              wire283 : reg294))) ?
          reg309 : (8'hb2)));
      if ($unsigned((reg298[(1'h0):(1'h0)] | (^~(8'h9c)))))
        begin
          reg314 <= reg299;
          reg315 <= $unsigned($signed(($unsigned(reg308) ?
              wire312 : (reg297 ? wire304 : ((7'h40) ? reg314 : reg294)))));
          if ($signed(((((reg303 + (8'ha7)) < $unsigned(reg313)) ^~ reg309[(2'h2):(2'h2)]) > $signed(wire306[(1'h1):(1'h0)]))))
            begin
              reg316 <= (~&$unsigned($signed($unsigned(wire305))));
              reg317 <= reg289;
              reg318 <= $unsigned(((((wire281 >= (7'h42)) ?
                  reg315 : {reg293,
                      reg290}) ~^ $signed(reg292[(4'h9):(4'h8)])) >= $signed((reg293[(3'h4):(3'h4)] ?
                  $signed(reg303) : $unsigned(reg291)))));
            end
          else
            begin
              reg316 <= $signed($signed((-wire283[(1'h0):(1'h0)])));
              reg317 <= ({{$unsigned({reg290, wire304})}} | (wire279 ?
                  $unsigned(reg292[(3'h5):(3'h5)]) : ($signed($unsigned(reg285)) == $unsigned(((8'hb7) && reg301)))));
              reg318 <= {(-($unsigned((reg316 ~^ reg289)) ?
                      (reg314[(1'h0):(1'h0)] ?
                          (reg309 ? reg294 : reg294) : {wire307,
                              wire307}) : (!(8'h9c))))};
              reg319 <= (|(reg303 > (^~(~^(reg293 ? wire284 : (8'hb0))))));
              reg320 <= (~&(~&($unsigned($signed((8'hbe))) ?
                  ($signed((8'hb7)) ?
                      {wire279,
                          reg315} : (+reg317)) : (((8'h9c) && reg298) | reg309[(2'h3):(1'h1)]))));
            end
          reg321 <= wire283[(1'h1):(1'h0)];
          reg322 <= reg290;
        end
      else
        begin
          if ({$unsigned(wire296),
              {$signed(((reg286 >>> reg322) ?
                      ((8'ha9) ? reg293 : wire283) : reg318))}})
            begin
              reg314 <= $unsigned(($unsigned($unsigned((~|reg309))) >> (((&reg308) || (reg319 < (8'hbd))) ?
                  reg314[(2'h3):(1'h0)] : ($unsigned(wire283) ^~ reg308[(5'h13):(2'h2)]))));
              reg315 <= reg298;
              reg316 <= $unsigned($unsigned(reg321));
              reg317 <= (|($unsigned({{reg291, wire306}, $unsigned(wire280)}) ?
                  ($unsigned($signed(reg287)) ?
                      wire283[(2'h3):(1'h0)] : reg314[(3'h4):(2'h2)]) : $unsigned((&(&wire312)))));
              reg318 <= reg316[(1'h0):(1'h0)];
            end
          else
            begin
              reg314 <= ($signed((reg318 + reg308[(5'h12):(4'h8)])) ^~ (^~reg294[(2'h3):(1'h0)]));
              reg315 <= $unsigned((($unsigned(reg290[(2'h2):(1'h1)]) ?
                  (8'h9f) : (~&$unsigned(wire306))) | reg300[(1'h1):(1'h1)]));
              reg316 <= $signed(((^($unsigned(wire312) && reg295)) ?
                  $signed($unsigned((|(8'hb7)))) : (((reg313 <<< reg287) | (reg320 ?
                          reg315 : wire306)) ?
                      $unsigned($signed((8'hb6))) : ((reg322 ?
                              (8'h9c) : reg320) ?
                          reg290 : $unsigned((8'ha3))))));
            end
          reg319 <= reg308[(4'hc):(4'hb)];
        end
      reg323 <= (((($signed((7'h44)) ?
                  reg319[(4'hb):(3'h4)] : $unsigned(wire312)) ?
              reg308 : $unsigned($unsigned(wire306))) ?
          $unsigned(reg301[(2'h2):(2'h2)]) : $signed({$signed(reg302)})) << reg301[(1'h0):(1'h0)]);
    end
  assign wire324 = $signed(($signed(wire296[(3'h7):(3'h5)]) ?
                       reg313[(3'h7):(1'h0)] : reg298));
  always
    @(posedge clk) begin
      reg325 <= reg287[(1'h0):(1'h0)];
      reg326 <= (|($signed((^~$signed(reg315))) | {(&wire306),
          (^(reg301 ^~ wire312))}));
      reg327 <= $signed(reg301[(3'h5):(3'h4)]);
      reg328 <= ((wire312[(4'h8):(1'h1)] >>> (^~reg310)) <= {reg322,
          (({reg317} * reg320) ? $signed($unsigned((8'hb2))) : wire324)});
    end
endmodule

module module229_1
#(parameter param271 = (-(((((8'hbb) ? (8'hb2) : (8'ha4)) && {(8'ha0)}) ? (!((8'h9c) ? (8'hae) : (8'haa))) : (((8'hbb) && (8'ha7)) ? {(8'hb0)} : ((8'hab) & (8'hbd)))) >= ((8'ha0) == ((8'hb8) ? ((8'hb2) & (8'haa)) : (8'ha4))))), 
parameter param272 = (!(^param271)))
(y, clk, wire233, wire232, wire231, wire230);
  output wire [(32'h1c0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire233;
  input wire [(2'h2):(1'h0)] wire232;
  input wire signed [(2'h2):(1'h0)] wire231;
  input wire [(5'h14):(1'h0)] wire230;
  wire signed [(4'h8):(1'h0)] wire257;
  wire signed [(4'hc):(1'h0)] wire256;
  wire [(2'h3):(1'h0)] wire239;
  wire [(3'h4):(1'h0)] wire238;
  wire signed [(5'h15):(1'h0)] wire237;
  wire signed [(4'hf):(1'h0)] wire236;
  wire [(4'h9):(1'h0)] wire235;
  wire signed [(4'h9):(1'h0)] wire234;
  reg [(5'h10):(1'h0)] reg270 = (1'h0);
  reg [(3'h5):(1'h0)] reg269 = (1'h0);
  reg [(3'h5):(1'h0)] reg268 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg267 = (1'h0);
  reg [(5'h14):(1'h0)] reg266 = (1'h0);
  reg [(5'h11):(1'h0)] reg265 = (1'h0);
  reg [(4'ha):(1'h0)] reg264 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg263 = (1'h0);
  reg [(4'hc):(1'h0)] reg262 = (1'h0);
  reg [(4'hf):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg258 = (1'h0);
  reg [(4'hc):(1'h0)] reg255 = (1'h0);
  reg [(5'h11):(1'h0)] reg254 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg253 = (1'h0);
  reg [(4'hb):(1'h0)] reg252 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg251 = (1'h0);
  reg [(4'he):(1'h0)] reg250 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg249 = (1'h0);
  reg [(5'h13):(1'h0)] reg248 = (1'h0);
  reg [(5'h15):(1'h0)] reg247 = (1'h0);
  reg [(2'h2):(1'h0)] reg246 = (1'h0);
  reg [(5'h13):(1'h0)] reg245 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg243 = (1'h0);
  reg [(3'h4):(1'h0)] reg242 = (1'h0);
  reg [(3'h7):(1'h0)] reg241 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg240 = (1'h0);
  assign y = {wire257,
                 wire256,
                 wire239,
                 wire238,
                 wire237,
                 wire236,
                 wire235,
                 wire234,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 (1'h0)};
  assign wire234 = ({wire232[(2'h2):(1'h1)]} ?
                       ($signed($unsigned(((8'hbc) ?
                           wire232 : wire230))) < $signed({$unsigned(wire232)})) : $unsigned($unsigned($signed(((8'hb3) ?
                           wire230 : wire231)))));
  assign wire235 = (wire232 & $signed(wire231));
  assign wire236 = (|(~wire234[(4'h8):(2'h2)]));
  assign wire237 = $signed($unsigned(($signed((^wire236)) ~^ $unsigned($unsigned((8'hb4))))));
  assign wire238 = $signed(wire231);
  assign wire239 = (&{{wire231[(2'h2):(1'h0)]}});
  always
    @(posedge clk) begin
      if ($signed(((^~wire237[(5'h10):(4'h8)]) ?
          (8'ha2) : ($unsigned($signed((8'ha3))) ?
              wire230[(1'h1):(1'h0)] : (wire232 ?
                  (^~wire237) : (wire233 ? wire232 : wire231))))))
        begin
          reg240 <= ({$unsigned(($unsigned((8'h9d)) - (wire235 ?
                      wire239 : wire239))),
                  wire239[(1'h1):(1'h0)]} ?
              {((wire236 ? (~|wire231) : $unsigned(wire232)) ?
                      ((~&wire231) & wire236) : ((wire231 ?
                          (8'hb0) : wire233) && $unsigned((8'hbd)))),
                  (+$unsigned((wire234 < (8'hba))))} : ((8'ha0) & $signed({(8'hb4)})));
          reg241 <= $unsigned({$unsigned(wire234),
              (wire235[(3'h7):(2'h3)] >= wire237)});
          if ((wire234[(3'h7):(1'h1)] || (&(8'hbc))))
            begin
              reg242 <= $signed((($unsigned(reg241) > ($unsigned(wire230) ~^ (wire231 > wire230))) ?
                  (~^wire238) : reg240));
              reg243 <= $signed(((wire234[(3'h7):(2'h3)] ?
                      {(wire232 ? wire230 : wire239),
                          $signed(wire232)} : reg240[(2'h2):(1'h0)]) ?
                  {(7'h44)} : $signed(({reg242} >= {reg240, wire233}))));
              reg244 <= (~&$unsigned($unsigned($unsigned(wire238))));
              reg245 <= ($signed((~&$signed((&wire233)))) ^~ wire234[(3'h4):(1'h1)]);
              reg246 <= wire233[(1'h1):(1'h0)];
            end
          else
            begin
              reg242 <= reg241;
              reg243 <= (~&((~|(-$unsigned(reg243))) ?
                  (^(~^$signed(reg245))) : ($signed(wire230) ?
                      ((reg241 != wire234) ?
                          wire233[(2'h2):(1'h0)] : (wire233 ?
                              (8'hbb) : reg240)) : ((~|(8'ha4)) & $signed(reg243)))));
            end
        end
      else
        begin
          reg240 <= ((wire234[(4'h8):(3'h4)] < wire238) ^~ (-(^~{(~^wire235)})));
          reg241 <= {reg244,
              {(wire233[(2'h2):(2'h2)] ?
                      (^~$signed(wire235)) : ((reg241 && reg246) ?
                          reg245[(4'hf):(4'hb)] : (wire234 ^ reg240)))}};
          if ((^($signed((+$signed(wire239))) != ((|(8'ha7)) && ((wire233 ?
                  reg246 : wire235) ?
              (wire231 <= (8'h9c)) : (wire230 >> wire234))))))
            begin
              reg242 <= $signed((wire238 ?
                  wire234[(1'h1):(1'h1)] : $signed(reg243)));
              reg243 <= (((+reg246) <= $unsigned(((~wire236) && (wire236 >> (8'hac))))) || (($signed(reg242[(2'h2):(1'h0)]) ?
                      wire237 : $unsigned((wire230 | wire233))) ?
                  $unsigned(wire233[(1'h0):(1'h0)]) : $unsigned($unsigned((wire237 ?
                      wire238 : reg245)))));
              reg244 <= (|$signed((($unsigned(wire235) ?
                  {wire233, reg244} : (~|reg246)) | (wire237 ?
                  (8'hb6) : (wire239 == (7'h41))))));
            end
          else
            begin
              reg242 <= (~(7'h41));
              reg243 <= reg241;
            end
          reg245 <= $signed($signed((+($unsigned((8'ha9)) ?
              wire239 : ((8'haa) ? wire234 : wire235)))));
        end
      if ((+(8'ha4)))
        begin
          if ({((^((^wire235) ? (8'ha2) : reg245)) <= (|{reg240})),
              (|(((wire238 ? wire237 : (8'ha7)) ?
                  wire238[(3'h4):(2'h2)] : reg242) > (+wire233[(1'h0):(1'h0)])))})
            begin
              reg247 <= (-((((wire232 * wire238) > (!wire233)) * wire237) ?
                  wire232[(1'h0):(1'h0)] : ((reg244 ? (~^wire231) : (-reg242)) ?
                      {(wire235 <= wire231)} : (~^reg242))));
              reg248 <= {(~&$unsigned(reg242[(1'h0):(1'h0)])),
                  ($unsigned($unsigned((~&(7'h40)))) ?
                      (~&$signed(reg240[(1'h1):(1'h1)])) : ((+(-reg242)) ?
                          reg246[(1'h1):(1'h0)] : ((wire239 ?
                              reg245 : wire231) && wire230[(5'h10):(2'h3)])))};
              reg249 <= $unsigned((-wire232));
            end
          else
            begin
              reg247 <= (~|($unsigned(($signed(wire236) - {reg249,
                  (7'h40)})) >>> (($signed(reg241) ?
                  $signed(wire233) : (&reg248)) + $unsigned(wire237[(3'h6):(1'h1)]))));
            end
        end
      else
        begin
          reg247 <= (8'hbc);
          if ($unsigned((wire237 ?
              $signed($signed((~(7'h43)))) : (({reg249} >> (|wire233)) ?
                  (wire234 ?
                      $unsigned((8'ha3)) : $signed(reg247)) : reg243[(5'h13):(3'h4)]))))
            begin
              reg248 <= (~|wire235[(3'h4):(3'h4)]);
              reg249 <= wire239;
              reg250 <= wire233;
              reg251 <= reg243;
            end
          else
            begin
              reg248 <= $signed(wire236);
              reg249 <= reg245[(4'hb):(1'h0)];
            end
          reg252 <= reg246;
          reg253 <= (^~{({(^wire237)} * ($signed(wire234) ?
                  $signed(reg240) : (reg242 << reg244)))});
          reg254 <= $unsigned((|(reg243 >>> (~^reg243[(4'h9):(3'h6)]))));
        end
      reg255 <= ($signed((wire231[(1'h0):(1'h0)] ?
          (~^reg250[(4'h8):(3'h4)]) : $unsigned((reg247 ?
              (8'hb8) : wire235)))) > (&reg250));
    end
  assign wire256 = ($unsigned($signed((&reg252))) << (reg246 ?
                       reg249[(3'h5):(1'h1)] : (reg249[(3'h5):(1'h1)] != (|$signed(reg242)))));
  assign wire257 = $unsigned(((((reg253 ?
                           wire230 : wire230) * $unsigned((8'hba))) ?
                       wire231 : (~&$unsigned(reg246))) >= reg253[(2'h2):(2'h2)]));
  always
    @(posedge clk) begin
      if (reg249[(3'h4):(2'h2)])
        begin
          reg258 <= ($unsigned(({(!wire256)} >> reg243[(4'ha):(2'h3)])) ?
              $unsigned($unsigned(((~&(7'h43)) ?
                  ((8'hb6) > reg246) : ((8'haa) ?
                      reg252 : (8'hbb))))) : {$unsigned({{reg251, reg254},
                      $signed(reg241)})});
          reg259 <= ((8'hb1) ?
              {(!$unsigned($unsigned(wire233))),
                  wire233[(3'h6):(2'h3)]} : (wire234 <<< {((wire235 ?
                      reg252 : reg249) - wire234[(4'h8):(4'h8)]),
                  (((8'hb2) ? wire238 : reg243) && reg252)}));
          if ((&{(~&$unsigned($unsigned(reg244))), reg240[(1'h0):(1'h0)]}))
            begin
              reg260 <= $unsigned(($signed(wire233) ?
                  (-$signed(reg249[(1'h1):(1'h1)])) : $unsigned(reg250[(3'h6):(1'h1)])));
            end
          else
            begin
              reg260 <= (^($signed($signed((wire239 != reg243))) <= {(~|(-reg243)),
                  reg252[(2'h3):(2'h2)]}));
              reg261 <= wire236[(4'hd):(4'ha)];
              reg262 <= reg261;
              reg263 <= {wire257[(2'h3):(2'h3)], reg255};
            end
          if (($unsigned(reg250) & (~|($unsigned(reg259) ?
              (^(wire234 <<< wire236)) : wire236[(4'ha):(2'h3)]))))
            begin
              reg264 <= $signed((&{((reg251 ? wire237 : reg240) ?
                      (^wire236) : $unsigned(wire256))}));
              reg265 <= $unsigned(($unsigned(wire238[(2'h2):(1'h1)]) ^~ {$unsigned(reg246),
                  $unsigned(reg242)}));
              reg266 <= $signed($unsigned(($signed($signed(reg265)) != ($unsigned(reg253) ?
                  wire257 : $unsigned(wire235)))));
              reg267 <= $unsigned({({reg265[(2'h2):(2'h2)]} >>> (reg261[(3'h5):(1'h1)] ?
                      reg266 : {reg241, (8'hb2)}))});
            end
          else
            begin
              reg264 <= ($signed(($unsigned((-(8'hb0))) ?
                      $unsigned($unsigned(reg260)) : $signed((wire230 ?
                          reg264 : wire257)))) ?
                  {reg249[(2'h3):(2'h2)],
                      $signed($unsigned({(8'hbf), reg252}))} : (~reg242));
              reg265 <= (~&(wire236 ?
                  $unsigned(wire230) : ((8'ha8) < reg264[(1'h0):(1'h0)])));
              reg266 <= (!($signed($signed(((7'h40) <<< wire231))) ?
                  (~(+(+wire234))) : $unsigned(reg265)));
            end
        end
      else
        begin
          if ({$unsigned({$signed(reg242[(3'h4):(2'h2)]), $signed(wire235)})})
            begin
              reg258 <= (8'hac);
            end
          else
            begin
              reg258 <= (8'hb1);
              reg259 <= ($signed(reg254) ?
                  $signed(($unsigned((wire232 <= wire232)) == ((reg249 == reg247) <<< {reg261}))) : $unsigned(reg264));
              reg260 <= reg249;
            end
        end
      reg268 <= wire238[(1'h1):(1'h1)];
      reg269 <= ($signed(($unsigned((reg260 <<< wire239)) ?
          ($unsigned(reg254) ?
              reg266[(4'hc):(4'ha)] : $signed((8'hae))) : reg244)) ^~ ((((wire237 ?
                  wire257 : reg251) ?
              $unsigned((7'h43)) : wire230) ?
          $unsigned(wire234) : reg261) & $signed(({reg261} < (reg252 || reg245)))));
      reg270 <= (~(8'hb1));
    end
endmodule

module module183_1
#(parameter param205 = {(((((8'hb6) - (8'hac)) ? (!(8'h9c)) : ((8'h9d) ? (7'h40) : (8'hb8))) || (((8'ha0) ? (7'h40) : (7'h41)) ? {(8'hac)} : (|(8'hb8)))) ? ((~&((8'hb9) ? (8'hbb) : (8'haf))) ? ((&(8'hba)) ? (8'h9e) : ((8'hbd) ? (7'h41) : (8'hb3))) : (+(8'hae))) : ((8'hbb) ? {((8'hb9) ? (8'hb2) : (8'ha5)), ((8'h9e) <= (7'h42))} : ((&(8'hbb)) << (8'hb7))))}, 
parameter param206 = ({param205, ((param205 & (param205 ? param205 : param205)) ? param205 : (param205 | param205))} ? (param205 ? (!((param205 ? param205 : param205) << (^param205))) : param205) : ((((param205 ? param205 : param205) ? (param205 * param205) : (param205 ? (8'hbf) : param205)) == ((param205 >= (8'ha9)) ? (&param205) : (7'h43))) == {(param205 ? (~&(8'ha8)) : (param205 ^~ param205)), (param205 ? (param205 ? param205 : param205) : (param205 ? param205 : (8'hbf)))})))
(y, clk, wire188, wire187, wire186, wire185, wire184);
  output wire [(32'hc2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire188;
  input wire [(4'he):(1'h0)] wire187;
  input wire signed [(5'h11):(1'h0)] wire186;
  input wire [(5'h14):(1'h0)] wire185;
  input wire [(4'hc):(1'h0)] wire184;
  wire signed [(3'h6):(1'h0)] wire204;
  wire signed [(4'he):(1'h0)] wire197;
  wire signed [(5'h12):(1'h0)] wire196;
  wire signed [(4'h8):(1'h0)] wire195;
  wire [(4'ha):(1'h0)] wire194;
  wire [(4'he):(1'h0)] wire193;
  wire [(4'hc):(1'h0)] wire192;
  wire signed [(4'hc):(1'h0)] wire191;
  wire signed [(5'h10):(1'h0)] wire190;
  wire signed [(5'h13):(1'h0)] wire189;
  reg [(4'h8):(1'h0)] reg203 = (1'h0);
  reg [(4'h8):(1'h0)] reg202 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg201 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg200 = (1'h0);
  reg [(2'h2):(1'h0)] reg199 = (1'h0);
  reg [(5'h14):(1'h0)] reg198 = (1'h0);
  assign y = {wire204,
                 wire197,
                 wire196,
                 wire195,
                 wire194,
                 wire193,
                 wire192,
                 wire191,
                 wire190,
                 wire189,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 (1'h0)};
  assign wire189 = (^wire184);
  assign wire190 = $unsigned(((($signed(wire186) ?
                           {wire185} : (wire185 < wire185)) ~^ $unsigned((7'h41))) ?
                       (wire184[(3'h6):(1'h0)] >>> $unsigned(((8'h9d) < wire186))) : ($signed(wire184[(3'h7):(1'h0)]) << (((8'hbb) ?
                               wire187 : (8'ha4)) ?
                           (wire184 ? wire184 : wire188) : wire189))));
  assign wire191 = $signed((~&(~^(8'hb2))));
  assign wire192 = ((^$unsigned(wire189[(1'h1):(1'h0)])) ?
                       (-wire190) : (+$signed($signed((8'ha2)))));
  assign wire193 = ($unsigned(wire185[(3'h7):(2'h3)]) ?
                       (^~(&wire186[(4'he):(4'ha)])) : {$unsigned({$signed((8'ha2))}),
                           $signed({$unsigned(wire190)})});
  assign wire194 = wire191[(2'h2):(1'h1)];
  assign wire195 = wire186;
  assign wire196 = $signed(wire190[(4'hb):(4'hb)]);
  assign wire197 = (wire192 & ($unsigned($signed(wire187[(1'h0):(1'h0)])) ?
                       $unsigned({$unsigned(wire188),
                           (~^wire195)}) : (~|$signed(wire188))));
  always
    @(posedge clk) begin
      reg198 <= wire195[(2'h3):(1'h0)];
      if (({$signed(wire192)} ? wire194 : wire187))
        begin
          reg199 <= $signed($unsigned(wire191[(3'h6):(1'h0)]));
          reg200 <= ({((~^$signed(wire188)) ?
                      $signed((^wire186)) : $unsigned((~&wire190))),
                  wire186[(3'h6):(1'h0)]} ?
              {(wire195 == $signed(wire193)),
                  $signed($signed((8'ha5)))} : $signed((($unsigned(wire193) ?
                      reg199 : reg198) ?
                  wire190 : ((~^(8'haa)) && ((7'h43) == wire187)))));
          reg201 <= wire185;
          reg202 <= wire189[(1'h0):(1'h0)];
          reg203 <= (~^($unsigned((~^reg202)) >= wire190[(3'h4):(3'h4)]));
        end
      else
        begin
          reg199 <= wire195[(3'h6):(2'h3)];
          reg200 <= wire197[(1'h0):(1'h0)];
          reg201 <= ((^(+{(reg202 ? reg201 : (8'ha0))})) != reg202);
          reg202 <= (~({$signed((wire192 ~^ wire188))} ?
              ({(^reg202), $signed(wire191)} ?
                  ((wire190 ? wire188 : wire190) ?
                      $unsigned(wire192) : $signed(reg202)) : (~|{wire193,
                      reg199})) : ((wire193[(3'h4):(2'h3)] ?
                  $signed(wire196) : $signed((8'ha0))) + $signed(wire196[(4'hf):(4'h9)]))));
        end
    end
  assign wire204 = ($unsigned(wire192) * reg199);
endmodule