(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param639 = (~^(8'hbf)))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h42):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire3;
  input wire [(4'hf):(1'h0)] wire2;
  input wire signed [(5'h15):(1'h0)] wire1;
  input wire signed [(5'h10):(1'h0)] wire0;
  wire signed [(3'h5):(1'h0)] wire638;
  wire [(2'h2):(1'h0)] wire636;
  wire [(5'h15):(1'h0)] wire8;
  wire [(3'h4):(1'h0)] wire7;
  wire [(4'h9):(1'h0)] wire4;
  reg signed [(4'hf):(1'h0)] reg6 = (1'h0);
  reg [(4'h9):(1'h0)] reg5 = (1'h0);
  assign y = {wire638, wire636, wire8, wire7, wire4, reg6, reg5, (1'h0)};
  assign wire4 = $unsigned(wire0);
  always
    @(posedge clk) begin
      reg5 <= $unsigned(wire0);
    end
  always
    @(posedge clk) begin
      reg6 <= $signed((wire3[(5'h15):(4'h9)] ?
          ((~^(-reg5)) >> ((&(8'h9f)) ?
              (7'h44) : (wire2 ? wire2 : (8'hbd)))) : (|(|wire2))));
    end
  assign wire7 = ((!(8'hb4)) ? reg6[(3'h5):(1'h1)] : wire4[(2'h2):(1'h0)]);
  assign wire8 = (~^$unsigned(($unsigned(wire3) * $unsigned($signed(wire0)))));
  module9 #() modinst637 (wire636, clk, wire2, wire1, wire0, wire8);
  assign wire638 = wire4;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module9
#(parameter param634 = ({(7'h43)} <<< {(~^(^~(~^(8'hb6))))}), 
parameter param635 = {((param634 ? param634 : param634) ^ (^(^~param634)))})
(y, clk, wire10, wire11, wire12, wire13);
  output wire [(32'h3cd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire10;
  input wire [(5'h12):(1'h0)] wire11;
  input wire signed [(4'hf):(1'h0)] wire12;
  input wire signed [(5'h15):(1'h0)] wire13;
  wire [(5'h12):(1'h0)] wire632;
  wire [(4'hc):(1'h0)] wire631;
  wire [(4'hb):(1'h0)] wire630;
  wire signed [(3'h4):(1'h0)] wire629;
  wire signed [(3'h5):(1'h0)] wire497;
  wire [(5'h13):(1'h0)] wire346;
  wire signed [(5'h15):(1'h0)] wire14;
  wire signed [(5'h14):(1'h0)] wire122;
  wire [(4'hd):(1'h0)] wire124;
  wire signed [(5'h10):(1'h0)] wire162;
  wire signed [(4'hc):(1'h0)] wire271;
  wire signed [(5'h14):(1'h0)] wire603;
  reg signed [(3'h4):(1'h0)] reg160 = (1'h0);
  reg [(4'h9):(1'h0)] reg157 = (1'h0);
  reg signed [(4'he):(1'h0)] reg155 = (1'h0);
  reg [(5'h10):(1'h0)] reg154 = (1'h0);
  reg [(3'h4):(1'h0)] reg152 = (1'h0);
  reg [(4'hd):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg148 = (1'h0);
  reg [(4'h8):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg144 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg143 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg137 = (1'h0);
  reg [(5'h12):(1'h0)] reg136 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg134 = (1'h0);
  reg [(4'he):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg129 = (1'h0);
  reg [(4'h9):(1'h0)] reg128 = (1'h0);
  reg [(4'hf):(1'h0)] reg499 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg606 = (1'h0);
  reg [(3'h6):(1'h0)] reg607 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg609 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg610 = (1'h0);
  reg [(4'hf):(1'h0)] reg613 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg614 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg615 = (1'h0);
  reg [(5'h14):(1'h0)] reg616 = (1'h0);
  reg [(5'h12):(1'h0)] reg617 = (1'h0);
  reg [(3'h6):(1'h0)] reg619 = (1'h0);
  reg [(3'h7):(1'h0)] reg620 = (1'h0);
  reg [(5'h15):(1'h0)] reg623 = (1'h0);
  reg [(4'hb):(1'h0)] reg625 = (1'h0);
  reg [(2'h2):(1'h0)] reg626 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg628 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar627 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg624 = (1'h0);
  reg [(4'h8):(1'h0)] forvar622 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg621 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg618 = (1'h0);
  reg [(5'h11):(1'h0)] reg612 = (1'h0);
  reg [(2'h3):(1'h0)] forvar606 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar612 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg611 = (1'h0);
  reg [(5'h12):(1'h0)] reg608 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg605 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg501 = (1'h0);
  reg [(4'hb):(1'h0)] forvar500 = (1'h0);
  reg [(3'h7):(1'h0)] reg161 = (1'h0);
  reg [(3'h4):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg156 = (1'h0);
  reg [(4'h9):(1'h0)] forvar153 = (1'h0);
  reg [(4'he):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg149 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg147 = (1'h0);
  reg [(4'h8):(1'h0)] forvar145 = (1'h0);
  reg [(3'h5):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg139 = (1'h0);
  reg [(2'h2):(1'h0)] forvar138 = (1'h0);
  reg [(5'h12):(1'h0)] reg133 = (1'h0);
  reg [(4'he):(1'h0)] forvar132 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg131 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg127 = (1'h0);
  reg [(5'h12):(1'h0)] forvar126 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar125 = (1'h0);
  assign y = {wire632,
                 wire631,
                 wire630,
                 wire629,
                 wire497,
                 wire346,
                 wire14,
                 wire122,
                 wire124,
                 wire162,
                 wire271,
                 wire603,
                 reg160,
                 reg157,
                 reg155,
                 reg154,
                 reg152,
                 reg151,
                 reg148,
                 reg146,
                 reg144,
                 reg143,
                 reg141,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg130,
                 reg129,
                 reg128,
                 reg499,
                 reg606,
                 reg607,
                 reg609,
                 reg610,
                 reg613,
                 reg614,
                 reg615,
                 reg616,
                 reg617,
                 reg619,
                 reg620,
                 reg623,
                 reg625,
                 reg626,
                 reg628,
                 forvar627,
                 reg624,
                 forvar622,
                 reg621,
                 reg618,
                 reg612,
                 forvar606,
                 forvar612,
                 reg611,
                 reg608,
                 reg605,
                 reg501,
                 forvar500,
                 reg161,
                 reg159,
                 reg158,
                 reg156,
                 forvar153,
                 reg150,
                 reg149,
                 reg147,
                 forvar145,
                 reg142,
                 reg140,
                 reg139,
                 forvar138,
                 reg133,
                 forvar132,
                 reg131,
                 reg127,
                 forvar126,
                 forvar125,
                 (1'h0)};
  assign wire14 = wire12;
  assign wire124 = wire13;
  always
    @(posedge clk) begin
      for (forvar125 = (1'h0); (forvar125 < (2'h3)); forvar125 = (forvar125 + (1'h1)))
        begin
          for (forvar126 = (1'h0); (forvar126 < (2'h3)); forvar126 = (forvar126 + (1'h1)))
            begin
              reg127 = (7'h40);
              reg128 <= {$unsigned((~^(wire12 ? wire122 : $unsigned(wire10)))),
                  (wire13[(4'h9):(4'h8)] ?
                      ($unsigned(wire11[(4'he):(4'he)]) <= ((reg127 ?
                          wire13 : wire11) != $signed(wire14))) : wire11)};
              reg129 <= ($unsigned((((reg127 ? forvar125 : wire11) ?
                      {wire10, reg127} : (wire12 ? wire13 : wire124)) ?
                  ($signed(wire12) ?
                      reg128 : $unsigned(wire124)) : $unsigned((8'hbd)))) ~^ ((!(&reg128)) ?
                  ((+$signed(wire14)) - ($signed((8'hb6)) < (wire12 ?
                      wire122 : reg128))) : wire11));
              reg130 <= ($signed(($unsigned($signed(wire124)) ?
                  $unsigned({wire124}) : ((forvar125 * wire11) ?
                      reg127 : $signed(reg129)))) <= (&$unsigned(($signed((8'hb5)) == reg129))));
              reg131 = ($signed((forvar126 ?
                  $unsigned($unsigned(wire14)) : $unsigned(wire124[(3'h4):(3'h4)]))) - ($unsigned(((reg129 ?
                          reg127 : wire12) ?
                      reg129 : $signed(reg129))) ?
                  $unsigned(({wire13,
                      wire11} <<< wire13[(4'h8):(2'h3)])) : $unsigned($unsigned($unsigned(reg128)))));
            end
          for (forvar132 = (1'h0); (forvar132 < (1'h0)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 = (forvar132 ? wire124[(4'ha):(3'h4)] : (~^reg127));
              reg134 <= wire11;
              reg135 <= $unsigned(wire10);
              reg136 <= wire14;
              reg137 <= wire14;
            end
          for (forvar138 = (1'h0); (forvar138 < (2'h2)); forvar138 = (forvar138 + (1'h1)))
            begin
              reg139 = ($unsigned($signed(wire122[(5'h10):(4'hc)])) ^~ {(|{wire14})});
              reg140 = forvar138;
            end
        end
      if (wire122[(4'hb):(4'ha)])
        begin
          reg141 <= $unsigned($signed((reg137 ? (7'h40) : (7'h44))));
        end
      else
        begin
          if ($unsigned((forvar125[(1'h1):(1'h1)] <<< forvar126)))
            begin
              reg142 = {(~|(|$signed($unsigned(reg141)))),
                  reg133[(4'h9):(2'h3)]};
            end
          else
            begin
              reg142 = (~|$unsigned($signed((+reg142))));
              reg143 <= $unsigned({$signed(wire10)});
              reg144 <= ((&(((wire124 ? reg134 : reg135) > reg137) ?
                      $signed($unsigned((8'hba))) : reg133)) ?
                  (forvar126[(4'hf):(1'h1)] ?
                      {reg134[(4'h9):(4'h9)],
                          ($unsigned(reg134) != forvar138[(1'h1):(1'h0)])} : (((~&reg137) ?
                          reg131 : wire13[(3'h4):(1'h0)]) ~^ ((wire124 ?
                          wire11 : reg128) <<< (reg142 ?
                          (8'hb2) : (8'ha8))))) : $signed($signed($signed(reg141[(3'h5):(3'h4)]))));
            end
          for (forvar145 = (1'h0); (forvar145 < (2'h3)); forvar145 = (forvar145 + (1'h1)))
            begin
              reg146 <= wire14[(4'hb):(1'h0)];
              reg147 = $signed($unsigned($signed($unsigned(wire122))));
            end
          if (((({reg143, (+reg133)} >> {reg146}) && {(^~wire12),
              $unsigned($unsigned(reg143))}) < (~^$unsigned((|(!reg129))))))
            begin
              reg148 <= {(wire11 ?
                      reg127[(3'h7):(3'h5)] : $unsigned(reg139[(2'h2):(1'h0)])),
                  (~|$signed((reg143[(4'hd):(4'h9)] ?
                      (reg135 ^ wire14) : (reg141 < reg137))))};
              reg149 = reg142[(3'h4):(2'h2)];
              reg150 = (reg142[(2'h3):(2'h3)] ^ $signed(wire13));
              reg151 <= ((reg139 >= $unsigned($unsigned($signed(reg144)))) ?
                  (~($signed($unsigned(reg142)) | forvar132)) : reg134);
              reg152 <= {(~^reg147), {reg144[(3'h5):(2'h2)], wire13}};
            end
          else
            begin
              reg148 <= reg140;
              reg149 = (wire122[(5'h13):(4'he)] ?
                  $unsigned($unsigned(($unsigned(forvar125) & (reg133 ?
                      wire122 : (8'hb1))))) : (forvar132 ?
                      (reg130 - $signed({forvar132,
                          reg148})) : $unsigned($signed({reg135}))));
            end
        end
      for (forvar153 = (1'h0); (forvar153 < (2'h3)); forvar153 = (forvar153 + (1'h1)))
        begin
          if ((-{forvar153}))
            begin
              reg154 <= ((wire12 ~^ $signed($signed({reg129}))) ?
                  ($unsigned(((wire124 ? forvar153 : wire11) ?
                          $signed(reg140) : (^reg134))) ?
                      ((+(reg142 <<< reg133)) != reg127[(3'h4):(2'h3)]) : (reg130[(4'h8):(1'h1)] > $unsigned($unsigned(forvar138)))) : ($signed($signed({wire11,
                          reg152})) ?
                      reg134 : ((reg131 ^ reg135[(1'h1):(1'h1)]) ?
                          (reg131 ?
                              $unsigned(forvar145) : (reg137 <= reg150)) : (^~(!reg139)))));
              reg155 <= $unsigned(((reg144 >>> {$signed(reg136)}) != ((&(wire14 || reg134)) ^~ $unsigned((reg136 ?
                  reg140 : reg131)))));
              reg156 = ((wire10[(4'ha):(4'h8)] ? wire14 : forvar138) ?
                  wire124 : {$unsigned(reg155), reg143});
            end
          else
            begin
              reg154 <= reg129;
              reg156 = (7'h44);
              reg157 <= $unsigned($signed(($unsigned(reg130[(4'ha):(4'h9)]) ~^ ($signed(reg148) * reg133[(5'h12):(4'h8)]))));
              reg158 = ($unsigned(reg134) ^ $unsigned((^~reg139)));
            end
          reg159 = (forvar126[(4'hd):(1'h1)] >>> $unsigned((((forvar153 ?
                      reg152 : reg137) ?
                  reg150 : $unsigned(reg140)) ?
              (7'h42) : forvar126)));
          reg160 <= $signed($signed($unsigned(forvar138)));
          reg161 = {({((^~(8'hb2)) && {reg128})} - reg137[(4'ha):(3'h4)])};
        end
    end
  assign wire162 = (($unsigned((8'hbf)) ?
                       {reg130[(4'h8):(4'h8)]} : reg152[(2'h2):(1'h1)]) >>> wire11);
   module273 #() modinst347 (wire346, clk, wire10, reg137, wire122, reg130);
  always
    @(posedge clk) begin
      reg499 <= $unsigned(($unsigned($unsigned($unsigned(reg134))) ?
          {reg144, wire11[(3'h6):(2'h2)]} : wire13));
      for (forvar500 = (1'h0); (forvar500 < (2'h3)); forvar500 = (forvar500 + (1'h1)))
        begin
          reg501 = ($unsigned(reg141) != $signed(wire346[(4'ha):(3'h5)]));
        end
    end
  module502 #() modinst604 (wire603, clk, reg129, wire122, reg136, reg143, reg144);
  always
    @(posedge clk) begin
      if (reg143)
        begin
          reg605 = ((($signed((wire271 ?
                  wire271 : (8'h9e))) & (wire162[(4'h8):(2'h3)] >> (wire346 != wire124))) * reg144[(2'h2):(1'h0)]) ?
              wire13[(3'h7):(2'h2)] : $unsigned({reg137,
                  reg136[(3'h5):(2'h2)]}));
          if ((reg141[(3'h5):(1'h0)] - $signed($unsigned(reg605))))
            begin
              reg606 <= (reg143 << ($signed($unsigned((reg152 ?
                      reg136 : reg144))) ?
                  (~&reg130) : wire271));
              reg607 <= reg499[(4'hc):(3'h6)];
              reg608 = wire162[(3'h4):(1'h0)];
              reg609 <= (({{(reg157 >>> (8'ha0))}} ^~ ($unsigned($unsigned(reg136)) ?
                      $unsigned((reg136 ?
                          wire603 : reg136)) : reg135[(3'h7):(3'h5)])) ?
                  ($unsigned(({wire10, reg148} ?
                      {reg608,
                          reg151} : reg136[(3'h4):(1'h0)])) && $signed(({reg157,
                      wire162} + (8'ha7)))) : ((~|(-(~|wire122))) && (wire603 ?
                      (8'ha3) : reg155)));
            end
          else
            begin
              reg606 <= reg129[(5'h13):(5'h11)];
              reg608 = $signed(reg134);
              reg609 <= (reg151 ~^ ((((reg499 ? reg143 : reg151) && wire10) ?
                  {$unsigned(wire10), reg155} : (((8'ha5) ?
                      reg137 : reg128) | wire603[(3'h4):(3'h4)])) >>> ($unsigned(wire13[(5'h14):(1'h0)]) ?
                  $unsigned(reg129[(2'h3):(1'h1)]) : reg141)));
              reg610 <= $signed(wire603);
              reg611 = {($signed((|reg610)) ?
                      $unsigned((8'hb4)) : (+((reg160 ?
                          wire162 : (8'hbb)) + reg137))),
                  {reg605, $signed((reg144[(5'h11):(4'ha)] ~^ reg146))}};
            end
          for (forvar612 = (1'h0); (forvar612 < (2'h2)); forvar612 = (forvar612 + (1'h1)))
            begin
              reg613 <= ($signed((^~wire271)) ?
                  {($signed($unsigned(wire11)) > $unsigned($unsigned(reg143)))} : $signed(reg134));
              reg614 <= $unsigned(wire162[(4'ha):(3'h6)]);
            end
        end
      else
        begin
          reg605 = ($signed($unsigned((~|(^wire271)))) && reg141);
          for (forvar606 = (1'h0); (forvar606 < (1'h0)); forvar606 = (forvar606 + (1'h1)))
            begin
              reg608 = {$signed(wire12),
                  $signed($signed($signed($unsigned(reg128))))};
              reg611 = ($signed($signed(($unsigned(reg609) - wire346))) + (-((8'hb4) + reg607)));
              reg612 = wire603;
              reg613 <= forvar606;
            end
          reg614 <= ((((~|(reg129 ? reg611 : reg134)) == {$signed(reg152),
                  ((8'hab) ? wire10 : reg608)}) ?
              $unsigned($unsigned(reg148[(2'h3):(1'h1)])) : ($signed($unsigned((8'hb5))) ?
                  (!(~forvar612)) : reg610[(1'h0):(1'h0)])) << reg144[(3'h6):(2'h2)]);
          reg615 <= (wire10 <= $unsigned($signed($unsigned((wire124 ?
              wire162 : reg605)))));
          if (reg157)
            begin
              reg616 <= {(reg613 ?
                      wire11 : $signed($unsigned({(8'hab), reg136}))),
                  reg137};
              reg617 <= $unsigned($unsigned($signed($unsigned((8'ha3)))));
              reg618 = (-reg152);
              reg619 <= ($unsigned({$signed((reg608 ?
                      wire346 : reg144))}) ~^ $unsigned({({wire14} ?
                      (~|reg613) : (reg614 ? reg157 : (8'h9d))),
                  ($unsigned(reg616) + (~|reg141))}));
            end
          else
            begin
              reg616 <= $unsigned({reg136, reg144});
              reg618 = reg155;
              reg619 <= $unsigned(reg609[(4'h9):(1'h0)]);
              reg620 <= $unsigned((~&reg128[(2'h2):(1'h1)]));
            end
        end
    end
  always
    @(posedge clk) begin
      reg621 = wire14[(2'h3):(1'h0)];
      for (forvar622 = (1'h0); (forvar622 < (3'h4)); forvar622 = (forvar622 + (1'h1)))
        begin
          if ((!(~^reg148[(3'h5):(1'h1)])))
            begin
              reg623 <= $unsigned((($signed(reg137) >> ({reg155, reg621} ?
                      $unsigned(reg155) : reg607)) ?
                  ($unsigned((~&(8'hb6))) ?
                      forvar622[(3'h5):(1'h1)] : (-$signed(reg607))) : (^~wire346[(5'h12):(1'h1)])));
              reg624 = ((~$unsigned(((~reg141) ?
                  reg151 : $unsigned(wire603)))) * {(8'hb1)});
              reg625 <= forvar622;
            end
          else
            begin
              reg624 = reg128[(3'h4):(2'h3)];
              reg625 <= ((~|reg614) & (reg615 ?
                  (((-reg130) ^~ reg607) || ($unsigned(reg141) ^ $unsigned(reg134))) : $unsigned({(reg154 ?
                          wire497 : reg141)})));
              reg626 <= {($signed($signed((wire346 | wire12))) != {$unsigned($unsigned(reg620)),
                      ($unsigned(reg617) ?
                          $signed(reg606) : (reg141 ? (7'h43) : reg619))})};
            end
          for (forvar627 = (1'h0); (forvar627 < (3'h4)); forvar627 = (forvar627 + (1'h1)))
            begin
              reg628 = {(&reg152)};
            end
        end
    end
  assign wire629 = (!$unsigned((!$unsigned(reg137))));
  assign wire630 = {reg616, (|(~$signed((8'h9c))))};
  assign wire631 = wire12[(4'ha):(3'h6)];
  module502 #() modinst633 (.wire507(reg616), .wire505(reg148), .clk(clk), .wire503(reg617), .wire506(reg152), .wire504(reg625), .y(wire632));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module502
#(parameter param602 = {((&{(+(8'hbb))}) ? ((((8'hb5) ^ (8'ha9)) >>> ((8'haa) ? (8'ha9) : (8'ha9))) ~^ (!((8'h9c) << (8'hb0)))) : (~|((!(7'h40)) ~^ {(8'hba), (8'hb9)}))), (!((((8'hbc) ? (8'h9d) : (7'h43)) ? ((7'h43) ? (8'hb0) : (8'hbe)) : (!(8'hbe))) ? {((7'h42) ? (8'ha6) : (8'ha6))} : (^~((8'hbd) ? (8'hac) : (8'haa)))))})
(y, clk, wire507, wire506, wire505, wire504, wire503);
  output wire [(32'h488):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire507;
  input wire [(2'h3):(1'h0)] wire506;
  input wire signed [(5'h12):(1'h0)] wire505;
  input wire signed [(4'hb):(1'h0)] wire504;
  input wire [(5'h12):(1'h0)] wire503;
  wire [(4'h8):(1'h0)] wire574;
  wire [(2'h2):(1'h0)] wire542;
  wire [(4'ha):(1'h0)] wire541;
  reg signed [(5'h10):(1'h0)] reg601 = (1'h0);
  reg [(5'h12):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg597 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg596 = (1'h0);
  reg [(3'h6):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg593 = (1'h0);
  reg [(2'h3):(1'h0)] reg589 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg587 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg586 = (1'h0);
  reg [(5'h15):(1'h0)] reg584 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg576 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg579 = (1'h0);
  reg [(3'h7):(1'h0)] reg578 = (1'h0);
  reg [(3'h5):(1'h0)] reg577 = (1'h0);
  reg [(4'he):(1'h0)] reg567 = (1'h0);
  reg [(5'h15):(1'h0)] reg565 = (1'h0);
  reg [(5'h13):(1'h0)] reg562 = (1'h0);
  reg [(4'h9):(1'h0)] reg553 = (1'h0);
  reg [(4'he):(1'h0)] reg551 = (1'h0);
  reg [(5'h12):(1'h0)] reg550 = (1'h0);
  reg [(4'hf):(1'h0)] reg549 = (1'h0);
  reg [(2'h3):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg545 = (1'h0);
  reg [(3'h7):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg540 = (1'h0);
  reg [(4'hb):(1'h0)] reg535 = (1'h0);
  reg [(3'h7):(1'h0)] reg534 = (1'h0);
  reg [(4'hf):(1'h0)] reg533 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg531 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg522 = (1'h0);
  reg [(4'hb):(1'h0)] reg520 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg518 = (1'h0);
  reg [(5'h12):(1'h0)] reg515 = (1'h0);
  reg [(5'h14):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg510 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg599 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg598 = (1'h0);
  reg [(3'h5):(1'h0)] forvar594 = (1'h0);
  reg [(5'h15):(1'h0)] reg592 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg591 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg590 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar588 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg585 = (1'h0);
  reg [(5'h10):(1'h0)] reg583 = (1'h0);
  reg [(5'h14):(1'h0)] reg582 = (1'h0);
  reg [(5'h15):(1'h0)] reg581 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg580 = (1'h0);
  reg [(5'h11):(1'h0)] forvar576 = (1'h0);
  reg [(3'h6):(1'h0)] reg575 = (1'h0);
  reg [(3'h4):(1'h0)] reg573 = (1'h0);
  reg [(3'h7):(1'h0)] reg572 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg571 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg569 = (1'h0);
  reg [(3'h6):(1'h0)] forvar568 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar566 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg564 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar561 = (1'h0);
  reg [(5'h14):(1'h0)] reg560 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg559 = (1'h0);
  reg [(2'h2):(1'h0)] reg558 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg557 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar556 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar555 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg554 = (1'h0);
  reg [(4'h8):(1'h0)] reg552 = (1'h0);
  reg [(5'h12):(1'h0)] reg548 = (1'h0);
  reg [(4'hb):(1'h0)] reg547 = (1'h0);
  reg [(3'h7):(1'h0)] reg543 = (1'h0);
  reg [(3'h7):(1'h0)] forvar539 = (1'h0);
  reg [(2'h2):(1'h0)] reg538 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg537 = (1'h0);
  reg [(3'h6):(1'h0)] reg536 = (1'h0);
  reg [(3'h7):(1'h0)] forvar532 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg530 = (1'h0);
  reg [(4'he):(1'h0)] reg529 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg528 = (1'h0);
  reg [(4'ha):(1'h0)] reg526 = (1'h0);
  reg [(4'hb):(1'h0)] reg525 = (1'h0);
  reg [(5'h11):(1'h0)] reg524 = (1'h0);
  reg [(5'h14):(1'h0)] reg523 = (1'h0);
  reg [(5'h12):(1'h0)] reg521 = (1'h0);
  reg [(4'h8):(1'h0)] reg519 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg517 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg511 = (1'h0);
  reg [(4'he):(1'h0)] forvar510 = (1'h0);
  reg [(4'hf):(1'h0)] reg516 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg514 = (1'h0);
  reg [(5'h15):(1'h0)] reg512 = (1'h0);
  reg [(4'ha):(1'h0)] forvar511 = (1'h0);
  reg [(5'h13):(1'h0)] reg508 = (1'h0);
  assign y = {wire574,
                 wire542,
                 wire541,
                 reg601,
                 reg600,
                 reg597,
                 reg596,
                 reg595,
                 reg593,
                 reg589,
                 reg587,
                 reg586,
                 reg584,
                 reg576,
                 reg579,
                 reg578,
                 reg577,
                 reg567,
                 reg565,
                 reg562,
                 reg553,
                 reg551,
                 reg550,
                 reg549,
                 reg546,
                 reg545,
                 reg544,
                 reg540,
                 reg535,
                 reg534,
                 reg533,
                 reg531,
                 reg527,
                 reg522,
                 reg520,
                 reg518,
                 reg515,
                 reg513,
                 reg510,
                 reg509,
                 reg599,
                 reg598,
                 forvar594,
                 reg592,
                 reg591,
                 reg590,
                 forvar588,
                 reg585,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 forvar576,
                 reg575,
                 reg573,
                 reg572,
                 reg571,
                 reg570,
                 reg569,
                 forvar568,
                 forvar566,
                 reg564,
                 reg563,
                 forvar561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 forvar556,
                 forvar555,
                 reg554,
                 reg552,
                 reg548,
                 reg547,
                 reg543,
                 forvar539,
                 reg538,
                 reg537,
                 reg536,
                 forvar532,
                 reg530,
                 reg529,
                 reg528,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg521,
                 reg519,
                 reg517,
                 reg511,
                 forvar510,
                 reg516,
                 reg514,
                 reg512,
                 forvar511,
                 reg508,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg508 = $signed(($unsigned(((wire503 <= wire505) ?
          $unsigned(wire507) : (wire504 ?
              wire504 : wire503))) >>> $unsigned(wire504[(4'ha):(2'h3)])));
      if (reg508)
        begin
          reg509 <= $signed($unsigned((($unsigned(wire507) || $signed(wire504)) ?
              $unsigned($unsigned(wire503)) : (~$signed(wire505)))));
          reg510 <= ((8'ha0) ?
              reg508 : {($unsigned($signed(wire507)) || ($signed(wire504) ?
                      (wire504 ? wire506 : (8'hbd)) : $signed((8'ha7)))),
                  (reg508 ?
                      {wire506, wire506[(2'h3):(2'h3)]} : $unsigned((reg508 ?
                          reg509 : wire507)))});
          for (forvar511 = (1'h0); (forvar511 < (1'h1)); forvar511 = (forvar511 + (1'h1)))
            begin
              reg512 = $unsigned(($signed({reg508[(3'h4):(2'h3)]}) ?
                  (|(wire505 == wire503[(4'he):(3'h7)])) : forvar511));
              reg513 <= ((+wire507[(4'hd):(3'h5)]) <<< {{wire507, forvar511},
                  forvar511});
              reg514 = ($signed(wire507) ?
                  $signed((~^$signed((wire503 ^ forvar511)))) : wire504[(4'hb):(4'hb)]);
              reg515 <= ({wire505,
                  $unsigned((reg512 ?
                      ((7'h41) ?
                          forvar511 : forvar511) : reg514))} ^ ((({wire504,
                          forvar511} ?
                      wire503[(4'hd):(4'hb)] : $unsigned(reg508)) ?
                  $unsigned((wire506 | (8'hb2))) : (8'hbf)) >> $signed(($signed(reg509) >= $unsigned((8'hb5))))));
            end
          reg516 = wire504;
        end
      else
        begin
          reg509 <= {reg510, $signed($unsigned(((^reg516) >= reg508)))};
          for (forvar510 = (1'h0); (forvar510 < (1'h0)); forvar510 = (forvar510 + (1'h1)))
            begin
              reg511 = (|$unsigned($signed($signed((reg509 >>> wire505)))));
              reg513 <= (reg514 >> reg512);
              reg515 <= $unsigned(forvar511);
              reg516 = $unsigned(forvar510);
              reg517 = wire503[(2'h2):(1'h0)];
            end
          if (($signed($signed(wire504)) ?
              reg509[(3'h5):(1'h0)] : reg513[(2'h3):(1'h0)]))
            begin
              reg518 <= $unsigned(((reg508 ?
                      ($unsigned(reg516) ? wire507 : (~&reg513)) : forvar511) ?
                  (!(reg517 ?
                      $unsigned(reg510) : (reg508 ?
                          reg511 : reg515))) : (reg510[(4'h9):(3'h5)] ?
                      $signed(reg511[(4'hf):(4'he)]) : {$unsigned(wire505)})));
              reg519 = wire507[(4'he):(4'hb)];
              reg520 <= reg511[(5'h11):(4'hd)];
              reg521 = (!reg511);
            end
          else
            begin
              reg518 <= {reg518,
                  ($unsigned($signed((reg512 ?
                      wire507 : reg514))) || forvar510)};
              reg520 <= $unsigned((^~reg519));
              reg521 = $unsigned($unsigned($signed($signed(reg510))));
              reg522 <= $unsigned((~|reg516[(2'h2):(2'h2)]));
            end
          reg523 = $unsigned($signed($unsigned((reg518 || reg519))));
          if ((reg512 >> $signed($unsigned(wire504))))
            begin
              reg524 = ($unsigned($unsigned((~^reg518))) <= reg510);
              reg525 = (reg512[(3'h6):(3'h6)] ^ $unsigned(reg515));
              reg526 = ($unsigned(((8'hb1) ?
                      $signed((reg516 ?
                          reg518 : reg510)) : (~(reg517 - reg524)))) ?
                  reg517[(3'h5):(1'h0)] : $unsigned(wire506[(1'h1):(1'h1)]));
            end
          else
            begin
              reg527 <= reg516[(4'h9):(2'h3)];
              reg528 = (~&$unsigned(reg517));
              reg529 = ((~&($unsigned(reg512) ~^ (wire507[(5'h11):(1'h0)] >>> (reg524 ^ reg508)))) ?
                  ((~forvar510[(3'h7):(1'h0)]) >>> (&$unsigned($signed(wire504)))) : reg517);
              reg530 = $signed(forvar511);
              reg531 <= (+(reg526[(1'h0):(1'h0)] ^~ wire505));
            end
        end
      for (forvar532 = (1'h0); (forvar532 < (1'h0)); forvar532 = (forvar532 + (1'h1)))
        begin
          reg533 <= (+{((-$unsigned(reg508)) ?
                  reg522 : reg521[(4'hc):(1'h0)])});
          if ($unsigned((~(~&$unsigned($signed(forvar510))))))
            begin
              reg534 <= ({(~{$unsigned(wire504)}),
                      ((reg513 <= reg514) - ({reg524} - (~&reg524)))} ?
                  $signed(reg527[(3'h5):(3'h5)]) : (!$unsigned(($signed(reg518) ?
                      $signed(wire503) : (~&wire507)))));
              reg535 <= $unsigned(forvar532);
            end
          else
            begin
              reg536 = {{reg525}, reg520};
              reg537 = (((-reg512) == (~&reg522)) || {wire506});
            end
          reg538 = {(reg514 == $signed(((reg529 ?
                  reg515 : reg526) >> $signed(reg527))))};
        end
      for (forvar539 = (1'h0); (forvar539 < (1'h0)); forvar539 = (forvar539 + (1'h1)))
        begin
          reg540 <= (~|{reg528,
              ({$unsigned(reg521), {(8'hac)}} ?
                  reg533[(4'hd):(4'h9)] : (~|(reg538 ^ reg533)))});
        end
    end
  assign wire541 = $unsigned(reg531);
  assign wire542 = $unsigned(wire504[(4'h9):(3'h5)]);
  always
    @(posedge clk) begin
      if ($signed($unsigned($signed(({wire542, reg540} ?
          reg513[(3'h4):(2'h3)] : reg513)))))
        begin
          if ($signed($unsigned({(reg534[(1'h1):(1'h1)] ?
                  (!reg535) : $unsigned(wire503))})))
            begin
              reg543 = $signed($signed({($unsigned(reg534) < $unsigned(reg533)),
                  $unsigned($unsigned(wire503))}));
              reg544 <= (!({$unsigned((wire504 - reg520))} + $unsigned(((wire505 >>> reg518) ?
                  wire506 : (reg531 - wire507)))));
              reg545 <= ($unsigned($unsigned(($unsigned((8'ha5)) ?
                      (!(8'hb4)) : $signed(reg533)))) ?
                  reg510 : (reg518[(1'h1):(1'h1)] + reg518));
            end
          else
            begin
              reg544 <= $unsigned((^wire504));
              reg545 <= reg533;
              reg546 <= wire506;
            end
        end
      else
        begin
          reg544 <= ($unsigned($signed($signed($unsigned(wire503)))) >> (&reg535));
          reg547 = reg527[(3'h7):(3'h7)];
          if ($unsigned((!{(reg522[(3'h5):(2'h2)] - (wire542 | reg510))})))
            begin
              reg548 = wire542;
              reg549 <= $unsigned(($unsigned($signed(reg544)) ~^ (|reg527)));
              reg550 <= $unsigned(({reg544,
                      ($signed(wire505) ?
                          $signed(wire541) : ((8'h9e) & wire507))} ?
                  {$signed((reg544 ? (8'had) : reg527)),
                      $unsigned((-reg540))} : reg509));
              reg551 <= {$unsigned(reg535[(4'hb):(2'h2)])};
              reg552 = reg513;
            end
          else
            begin
              reg548 = $signed(wire506);
              reg549 <= $unsigned(reg543[(3'h4):(1'h1)]);
              reg550 <= $unsigned((~^wire506));
              reg551 <= $unsigned($unsigned(($unsigned((reg534 || reg549)) == reg551)));
              reg553 <= $unsigned(reg533[(4'h9):(1'h0)]);
            end
          reg554 = reg551;
        end
    end
  always
    @(posedge clk) begin
      for (forvar555 = (1'h0); (forvar555 < (3'h4)); forvar555 = (forvar555 + (1'h1)))
        begin
          for (forvar556 = (1'h0); (forvar556 < (3'h4)); forvar556 = (forvar556 + (1'h1)))
            begin
              reg557 = reg546;
              reg558 = (8'ha2);
              reg559 = $unsigned(forvar555);
              reg560 = {reg513, (reg553 ? wire505[(5'h10):(3'h7)] : reg515)};
            end
          for (forvar561 = (1'h0); (forvar561 < (3'h4)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 <= reg515;
              reg563 = reg545;
              reg564 = reg531[(1'h1):(1'h0)];
              reg565 <= (reg549[(2'h2):(1'h0)] <= (|($signed($signed((8'h9c))) ~^ $signed({reg557}))));
            end
          for (forvar566 = (1'h0); (forvar566 < (3'h4)); forvar566 = (forvar566 + (1'h1)))
            begin
              reg567 <= reg546;
            end
          for (forvar568 = (1'h0); (forvar568 < (2'h3)); forvar568 = (forvar568 + (1'h1)))
            begin
              reg569 = $unsigned((wire542 >= ($signed({reg518}) ?
                  $unsigned((^reg531)) : (reg509 ?
                      $unsigned(reg546) : $unsigned(wire504)))));
              reg570 = (reg509 ?
                  $unsigned($unsigned($signed($unsigned(forvar556)))) : wire503[(1'h1):(1'h0)]);
              reg571 = $signed($signed((8'hb7)));
              reg572 = wire506[(1'h0):(1'h0)];
            end
        end
      reg573 = {($unsigned(((&reg544) ? reg546 : {wire507, (8'hac)})) ?
              reg534 : (wire507 + $signed($signed(reg550))))};
    end
  assign wire574 = (|$unsigned($signed(reg544)));
  always
    @(posedge clk) begin
      if ((~^reg545[(4'hf):(4'hd)]))
        begin
          reg575 = reg549;
          for (forvar576 = (1'h0); (forvar576 < (1'h0)); forvar576 = (forvar576 + (1'h1)))
            begin
              reg577 <= $unsigned(reg567);
              reg578 <= (~^reg551);
            end
          reg579 <= $unsigned({reg540, $signed(wire542[(2'h2):(1'h1)])});
        end
      else
        begin
          reg575 = $unsigned($unsigned(reg534[(3'h7):(3'h7)]));
          reg576 <= $unsigned((~^$signed((wire503 >= (reg522 ?
              wire505 : (8'ha2))))));
          reg577 <= $unsigned(reg520);
          reg580 = (reg531 ?
              reg510 : (-((reg546 < {reg513, wire542}) ?
                  (|$signed(reg567)) : (-(reg518 ? reg567 : reg546)))));
          if (({(^~reg546)} ?
              {$signed($unsigned((reg551 ? reg518 : reg580))),
                  (($unsigned(forvar576) ?
                          $unsigned(reg546) : {reg576, reg515}) ?
                      reg522 : reg544)} : (!$unsigned(({wire574,
                  reg565} & $signed(wire542))))))
            begin
              reg581 = $signed({(~&wire542),
                  $unsigned($signed((reg550 ? reg531 : (8'hbb))))});
              reg582 = $signed($signed(((8'h9d) ?
                  ({wire506, wire542} ?
                      wire574 : $unsigned((8'hb4))) : (~^((8'hbc) ?
                      wire507 : (8'hba))))));
              reg583 = reg562;
            end
          else
            begin
              reg584 <= $signed(reg565[(4'h8):(1'h0)]);
              reg585 = (reg553[(1'h1):(1'h1)] && (reg578 ?
                  reg580[(1'h0):(1'h0)] : (8'ha3)));
            end
        end
    end
  always
    @(posedge clk) begin
      reg586 <= reg551[(3'h7):(2'h2)];
      reg587 <= ((~^{reg567}) ?
          reg544[(2'h3):(2'h3)] : (~|(($unsigned(reg522) ?
                  (reg533 ? reg562 : reg579) : (reg551 ? reg544 : reg531)) ?
              ($signed(wire504) ?
                  $signed(reg586) : ((8'hb6) || reg533)) : reg545[(4'h8):(2'h3)])));
      for (forvar588 = (1'h0); (forvar588 < (1'h1)); forvar588 = (forvar588 + (1'h1)))
        begin
          if (reg544[(1'h0):(1'h0)])
            begin
              reg589 <= (((reg522 <= (^$signed(wire503))) && ($unsigned(((7'h43) + reg586)) ?
                  ($unsigned(reg567) - (reg544 | wire574)) : $unsigned((8'ha8)))) != (+($unsigned({reg578}) > reg520[(4'ha):(4'h8)])));
            end
          else
            begin
              reg590 = (-(|$unsigned($unsigned($unsigned(reg518)))));
              reg591 = $unsigned((($signed($unsigned(reg589)) ?
                      $unsigned((reg587 * wire541)) : ($signed(wire542) ?
                          (wire504 != reg531) : $unsigned((8'had)))) ?
                  (~&reg533[(1'h1):(1'h0)]) : $unsigned((reg546 < (~reg587)))));
              reg592 = (reg544[(1'h0):(1'h0)] ?
                  (reg510[(2'h2):(2'h2)] <= (($signed(reg579) > reg584) * (reg531 ?
                      (~^reg578) : (reg544 & reg515)))) : ({$unsigned((reg515 ?
                              (8'h9f) : reg513))} ?
                      $signed((wire505[(4'he):(4'hb)] ?
                          $unsigned(wire506) : (+wire505))) : reg510));
              reg593 <= reg565[(3'h6):(1'h0)];
            end
          for (forvar594 = (1'h0); (forvar594 < (2'h3)); forvar594 = (forvar594 + (1'h1)))
            begin
              reg595 <= $unsigned(($unsigned((wire542 ?
                      $unsigned(reg545) : {(8'ha8)})) ?
                  (((reg576 << reg591) ?
                          (reg587 ? (7'h43) : reg565) : $unsigned(reg550)) ?
                      $unsigned((reg576 ?
                          (8'h9e) : reg510)) : reg527[(4'hc):(4'hb)]) : ($unsigned(reg520[(1'h1):(1'h1)]) <= $unsigned($unsigned(wire541)))));
            end
          if (((reg510 ?
              ((reg593 & (^(8'ha9))) != $signed(reg553)) : {$signed(reg509[(3'h6):(1'h0)])}) > ((reg595[(1'h1):(1'h1)] ?
                  $signed(reg578[(1'h1):(1'h1)]) : ((reg515 ?
                          wire541 : reg533) ?
                      {wire574, reg551} : $signed(reg590))) ?
              (($unsigned(reg577) <<< (~reg567)) ?
                  reg544 : (^~reg527)) : {$signed({(8'h9f), reg562}),
                  $unsigned($unsigned((8'hac)))})))
            begin
              reg596 <= $unsigned($signed(((^~reg509) ?
                  $unsigned($unsigned(reg584)) : $unsigned($unsigned(reg577)))));
              reg597 <= wire506[(1'h0):(1'h0)];
            end
          else
            begin
              reg598 = (8'hbf);
              reg599 = (7'h42);
              reg600 <= reg565[(4'h8):(2'h3)];
            end
        end
      reg601 <= reg599;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module273
#(parameter param344 = (8'ha5), 
parameter param345 = ({(8'ha0), ({(8'h9c), (7'h44)} <<< (|{param344, param344}))} ? (&param344) : {{(~{param344}), ((param344 * param344) ? param344 : (param344 || param344))}, param344}))
(y, clk, wire277, wire276, wire275, wire274);
  output wire [(32'h358):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire277;
  input wire [(3'h7):(1'h0)] wire276;
  input wire [(4'h8):(1'h0)] wire275;
  input wire [(4'he):(1'h0)] wire274;
  wire [(4'hb):(1'h0)] wire308;
  wire signed [(5'h10):(1'h0)] wire303;
  wire [(4'hd):(1'h0)] wire302;
  wire [(5'h10):(1'h0)] wire301;
  wire [(5'h13):(1'h0)] wire300;
  wire signed [(5'h12):(1'h0)] wire299;
  wire signed [(4'hf):(1'h0)] wire298;
  wire [(5'h14):(1'h0)] wire297;
  wire [(5'h11):(1'h0)] wire278;
  reg signed [(4'hf):(1'h0)] reg343 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg340 = (1'h0);
  reg [(3'h4):(1'h0)] reg339 = (1'h0);
  reg [(4'ha):(1'h0)] reg337 = (1'h0);
  reg [(3'h6):(1'h0)] reg336 = (1'h0);
  reg [(4'ha):(1'h0)] reg334 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg332 = (1'h0);
  reg [(3'h7):(1'h0)] reg331 = (1'h0);
  reg [(4'ha):(1'h0)] reg330 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg326 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg324 = (1'h0);
  reg [(4'h9):(1'h0)] reg323 = (1'h0);
  reg [(3'h4):(1'h0)] reg322 = (1'h0);
  reg [(5'h12):(1'h0)] reg321 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg319 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg314 = (1'h0);
  reg [(5'h12):(1'h0)] reg307 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg305 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg296 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg295 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg294 = (1'h0);
  reg [(4'h9):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg288 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg287 = (1'h0);
  reg [(5'h15):(1'h0)] reg286 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg285 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg284 = (1'h0);
  reg [(4'h9):(1'h0)] reg282 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg281 = (1'h0);
  reg [(4'h9):(1'h0)] reg280 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg342 = (1'h0);
  reg [(4'hc):(1'h0)] reg341 = (1'h0);
  reg [(3'h6):(1'h0)] reg338 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg335 = (1'h0);
  reg [(4'ha):(1'h0)] reg333 = (1'h0);
  reg [(4'h9):(1'h0)] reg329 = (1'h0);
  reg [(4'hb):(1'h0)] reg328 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg327 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg325 = (1'h0);
  reg [(4'hf):(1'h0)] reg320 = (1'h0);
  reg [(4'hc):(1'h0)] forvar317 = (1'h0);
  reg [(2'h2):(1'h0)] forvar311 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar309 = (1'h0);
  reg [(4'hb):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg317 = (1'h0);
  reg signed [(4'he):(1'h0)] reg316 = (1'h0);
  reg signed [(4'he):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg312 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg311 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar310 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg309 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg306 = (1'h0);
  reg [(4'ha):(1'h0)] reg292 = (1'h0);
  reg [(4'h9):(1'h0)] reg293 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar292 = (1'h0);
  reg [(5'h12):(1'h0)] forvar290 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg289 = (1'h0);
  reg [(5'h10):(1'h0)] reg283 = (1'h0);
  reg [(4'hd):(1'h0)] forvar279 = (1'h0);
  assign y = {wire308,
                 wire303,
                 wire302,
                 wire301,
                 wire300,
                 wire299,
                 wire298,
                 wire297,
                 wire278,
                 reg343,
                 reg340,
                 reg339,
                 reg337,
                 reg336,
                 reg334,
                 reg332,
                 reg331,
                 reg330,
                 reg326,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg319,
                 reg314,
                 reg307,
                 reg305,
                 reg304,
                 reg296,
                 reg295,
                 reg294,
                 reg291,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg282,
                 reg281,
                 reg280,
                 reg342,
                 reg341,
                 reg338,
                 reg335,
                 reg333,
                 reg329,
                 reg328,
                 reg327,
                 reg325,
                 reg320,
                 forvar317,
                 forvar311,
                 reg310,
                 forvar309,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg313,
                 reg312,
                 reg311,
                 forvar310,
                 reg309,
                 reg306,
                 reg292,
                 reg293,
                 forvar292,
                 forvar290,
                 reg289,
                 reg283,
                 forvar279,
                 (1'h0)};
  assign wire278 = (wire275[(2'h2):(2'h2)] - (^~$unsigned(((8'ha6) ?
                       (wire274 ? wire277 : wire275) : $unsigned((8'hbf))))));
  always
    @(posedge clk) begin
      for (forvar279 = (1'h0); (forvar279 < (1'h0)); forvar279 = (forvar279 + (1'h1)))
        begin
          if ((wire275 ?
              ($unsigned((&wire275)) ?
                  wire276[(3'h4):(1'h0)] : (^$unsigned(forvar279))) : wire278))
            begin
              reg280 <= wire278;
            end
          else
            begin
              reg280 <= (-($signed($unsigned($signed((8'hbb)))) ?
                  $signed(({wire277, wire274} >= {wire277,
                      wire278})) : wire277));
              reg281 <= $unsigned(($unsigned($signed((reg280 ~^ wire274))) ^~ {(wire275 ?
                      forvar279[(4'hb):(4'h9)] : (reg280 * reg280)),
                  {(wire277 ? (8'h9f) : wire277)}}));
              reg282 <= reg281;
              reg283 = $unsigned((~&wire274[(2'h2):(2'h2)]));
            end
          reg284 <= $unsigned(((+((~^reg280) <= (reg281 ? wire276 : reg282))) ?
              {$unsigned($signed(wire278)), {wire278}} : (+(+(8'ha5)))));
          reg285 <= (wire275 ?
              $unsigned((&reg282)) : (((wire276[(2'h2):(2'h2)] ?
                  $unsigned(wire274) : $unsigned(reg282)) >> reg283[(4'h8):(4'h8)]) ^ (~^forvar279)));
          if ((((!(wire278[(3'h7):(1'h1)] ~^ $unsigned(wire274))) * (wire276 ?
                  ((wire275 >> (8'ha6)) ?
                      $unsigned(reg283) : wire276[(3'h6):(3'h4)]) : $unsigned((wire274 ?
                      wire274 : wire274)))) ?
              (^forvar279) : wire275[(4'h8):(3'h4)]))
            begin
              reg286 <= $signed($signed(reg281));
              reg287 <= (($unsigned($signed((wire275 ? reg282 : reg281))) ?
                  $unsigned({(wire276 | (7'h43)),
                      $signed(reg284)}) : $unsigned({(forvar279 >>> reg283),
                      $unsigned(wire277)})) ~^ $unsigned((reg280 ?
                  {$unsigned(wire276)} : wire274)));
              reg288 <= wire278;
              reg289 = {(wire278 - (~^forvar279)), reg283[(3'h6):(3'h4)]};
            end
          else
            begin
              reg286 <= reg282;
              reg289 = ($unsigned(($unsigned(wire278[(2'h3):(2'h3)]) == wire274)) == $signed(reg285[(3'h4):(2'h2)]));
            end
        end
      for (forvar290 = (1'h0); (forvar290 < (1'h1)); forvar290 = (forvar290 + (1'h1)))
        begin
          reg291 <= $unsigned($unsigned(($unsigned({forvar290}) ?
              $signed((8'ha8)) : (forvar279 ? (8'hae) : reg285))));
        end
      if ((!$unsigned((+$unsigned(reg281)))))
        begin
          for (forvar292 = (1'h0); (forvar292 < (2'h3)); forvar292 = (forvar292 + (1'h1)))
            begin
              reg293 = (~&{{{(wire276 ? (8'haf) : reg282),
                          (forvar290 ? forvar292 : reg281)}},
                  (~^forvar279[(3'h5):(1'h1)])});
            end
        end
      else
        begin
          if ($unsigned(wire275[(3'h6):(3'h4)]))
            begin
              reg292 = reg281[(1'h0):(1'h0)];
            end
          else
            begin
              reg294 <= $signed((&(!$unsigned($unsigned((8'hab))))));
              reg295 <= ($signed((8'hab)) && reg286[(5'h13):(2'h3)]);
            end
          reg296 <= ($signed(forvar292) >> reg284);
        end
    end
  assign wire297 = (($signed(reg294) || $signed({wire278})) ?
                       (&$unsigned(wire278)) : $signed(reg291));
  assign wire298 = reg287[(1'h0):(1'h0)];
  assign wire299 = ((wire275 <<< wire298) ?
                       {{$unsigned($unsigned(reg282))}, (+reg282)} : (({wire298,
                           $unsigned(wire298)} - $signed($signed(reg285))) <<< reg281[(2'h3):(2'h2)]));
  assign wire300 = $signed(wire298);
  assign wire301 = (7'h44);
  assign wire302 = (~|(~|wire297[(5'h10):(3'h4)]));
  assign wire303 = reg287;
  always
    @(posedge clk) begin
      reg304 <= reg296;
      reg305 <= (wire301 ? $unsigned(reg282) : wire274);
      reg306 = $unsigned((reg296 ?
          (~$unsigned(reg280)) : $signed($unsigned((reg305 ~^ reg305)))));
      reg307 <= (~^$signed($unsigned((-$signed(reg282)))));
    end
  assign wire308 = $unsigned($unsigned((8'ha5)));
  always
    @(posedge clk) begin
      if (reg304)
        begin
          reg309 = $signed(reg282[(3'h6):(2'h2)]);
          for (forvar310 = (1'h0); (forvar310 < (2'h3)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 = wire301[(4'h9):(2'h3)];
              reg312 = $unsigned((-($signed($unsigned(reg288)) ?
                  {(!reg287)} : reg296)));
            end
          if (reg307)
            begin
              reg313 = (^~$unsigned((8'hab)));
              reg314 <= $unsigned((-reg291[(3'h4):(2'h2)]));
              reg315 = $unsigned(($unsigned({$signed(wire275)}) ?
                  reg294 : (((&wire308) ?
                          {reg284, wire303} : {reg313, reg287}) ?
                      (^~(reg280 ? reg309 : wire301)) : reg294)));
              reg316 = (wire276[(1'h1):(1'h0)] ?
                  $unsigned((^~wire299)) : ((reg305 ?
                          $unsigned(wire277) : reg291) ?
                      (^~((reg281 ? reg295 : (8'ha2)) ?
                          (reg311 ?
                              (8'ha3) : wire301) : wire277[(1'h1):(1'h1)])) : (wire302 == (|$signed((8'ha3))))));
            end
          else
            begin
              reg313 = $unsigned({$unsigned(($signed(reg286) ?
                      reg285 : (wire303 ? wire297 : reg281)))});
              reg315 = ($signed($unsigned(($signed(wire300) | (reg312 ?
                      reg313 : reg281)))) ?
                  $unsigned((~(&wire302[(4'hb):(2'h2)]))) : ($signed((!(reg284 ?
                      wire302 : wire275))) >> reg285));
              reg316 = reg291;
              reg317 = wire301[(3'h4):(1'h0)];
              reg318 = reg294[(3'h4):(3'h4)];
            end
        end
      else
        begin
          for (forvar309 = (1'h0); (forvar309 < (2'h3)); forvar309 = (forvar309 + (1'h1)))
            begin
              reg310 = (($signed((8'hbb)) > (^wire297)) ?
                  $unsigned($signed(reg314[(3'h6):(1'h1)])) : (-forvar310[(3'h4):(1'h1)]));
            end
          for (forvar311 = (1'h0); (forvar311 < (1'h1)); forvar311 = (forvar311 + (1'h1)))
            begin
              reg314 <= (wire308 | reg313[(4'h8):(3'h6)]);
              reg315 = (wire301 ?
                  $signed($unsigned((^(wire308 * reg291)))) : (($signed((&wire274)) ?
                          reg284 : reg313) ?
                      reg311 : (reg288 ~^ (~{reg309, wire301}))));
            end
          reg316 = {$unsigned(reg313), (~^(|$signed({reg304})))};
          for (forvar317 = (1'h0); (forvar317 < (2'h2)); forvar317 = (forvar317 + (1'h1)))
            begin
              reg319 <= reg288[(3'h6):(1'h0)];
              reg320 = (~&(~^(8'hb1)));
            end
          reg321 <= {wire299};
        end
      reg322 <= wire301[(4'hf):(4'he)];
      if ((^~wire275))
        begin
          if ($unsigned($signed($unsigned($unsigned($unsigned((8'h9e)))))))
            begin
              reg323 <= ($signed(reg284) != ($unsigned($unsigned($signed(forvar310))) == (($unsigned(wire277) ?
                      $signed(wire303) : (reg313 ^~ (8'hb4))) ?
                  $unsigned((~&forvar310)) : forvar309)));
              reg324 <= $signed((^reg309));
              reg325 = reg319[(4'h8):(3'h5)];
            end
          else
            begin
              reg325 = (reg312 ?
                  $signed(reg311) : ((|reg284) ~^ $signed({(reg288 >> forvar311)})));
              reg326 <= ($unsigned(reg287) ^ {(($signed(reg282) > (wire308 >= (8'hbe))) ?
                      {(reg317 <= reg319), wire303} : wire275),
                  $unsigned(reg324[(3'h4):(2'h2)])});
            end
          if (wire301)
            begin
              reg327 = $unsigned($unsigned($signed($unsigned(wire298[(4'h8):(3'h4)]))));
              reg328 = $signed(($signed($unsigned(reg311[(1'h0):(1'h0)])) > reg322));
              reg329 = $unsigned((8'hba));
              reg330 <= ($signed((!forvar311)) + $unsigned((~|((-reg314) + (|reg282)))));
              reg331 <= $unsigned(reg315);
            end
          else
            begin
              reg330 <= reg296;
              reg331 <= ({$signed($unsigned((-forvar311)))} ?
                  $unsigned({$signed((wire301 - reg328)),
                      ((reg315 && reg321) ?
                          reg282[(1'h0):(1'h0)] : reg327[(2'h2):(2'h2)])}) : (8'hbc));
              reg332 <= $unsigned(forvar311[(1'h0):(1'h0)]);
              reg333 = reg315;
              reg334 <= reg330[(3'h7):(3'h4)];
            end
        end
      else
        begin
          if ({($signed($unsigned(reg321[(4'hd):(4'hd)])) ?
                  (reg291 ? reg310 : reg329) : $unsigned({reg312[(3'h7):(1'h0)],
                      $unsigned((8'ha2))}))})
            begin
              reg325 = $signed($signed((|((reg294 ~^ reg294) ?
                  $unsigned(reg287) : reg309[(3'h4):(1'h1)]))));
              reg326 <= reg328;
            end
          else
            begin
              reg325 = (wire274[(3'h4):(1'h0)] ?
                  {reg284, reg288} : reg282[(3'h4):(2'h3)]);
              reg327 = $signed(reg334);
              reg330 <= forvar309;
              reg331 <= ((^~reg330) ?
                  $signed((reg330[(2'h2):(1'h1)] ?
                      (|$unsigned(reg319)) : wire299)) : ($unsigned(((wire275 != (8'ha4)) >>> $signed(wire303))) ^~ $signed(($unsigned(reg314) ?
                      (reg329 || wire302) : $signed((8'hac))))));
            end
          reg333 = $unsigned((-(~&forvar317)));
          if (((({(-reg294), {wire274}} ?
              (reg313[(3'h5):(1'h1)] >= reg309) : $signed(wire276)) >>> $unsigned({(wire303 ^~ reg327)})) && $unsigned((wire297 ?
              (reg316[(4'h9):(1'h1)] ?
                  (reg284 && wire298) : forvar317) : (-reg295[(2'h2):(1'h0)])))))
            begin
              reg334 <= reg280[(2'h2):(1'h0)];
              reg335 = (reg323 ?
                  forvar310 : $unsigned(($unsigned(wire274) ~^ $unsigned(reg291[(1'h0):(1'h0)]))));
              reg336 <= reg305[(1'h1):(1'h1)];
              reg337 <= (reg286[(1'h0):(1'h0)] ?
                  (wire301[(1'h1):(1'h1)] & $signed((|reg324[(4'h8):(1'h1)]))) : ($unsigned(((reg322 ?
                      reg280 : reg336) ^~ (reg312 | (8'had)))) >= reg334));
            end
          else
            begin
              reg334 <= $unsigned(reg291[(3'h6):(1'h1)]);
              reg336 <= ($unsigned($unsigned($signed(reg319))) ^ reg329);
              reg338 = reg296[(3'h5):(1'h1)];
              reg339 <= (reg326 <<< $unsigned((reg304[(2'h2):(1'h1)] > reg281)));
            end
          reg340 <= $unsigned(wire276);
          reg341 = ($unsigned((reg338 ?
                  {reg331, (8'hbb)} : $unsigned($signed(wire297)))) ?
              $unsigned({$unsigned(wire275),
                  (!{reg296})}) : ((reg287[(1'h0):(1'h0)] ?
                      {$unsigned(reg285),
                          $unsigned(reg284)} : $signed((8'haf))) ?
                  reg338[(1'h1):(1'h0)] : (wire297 ?
                      (~^$signed(reg332)) : wire299)));
        end
      reg342 = reg287;
      reg343 <= $signed($signed(reg342[(2'h3):(2'h3)]));
    end
endmodule
