(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param394 = (^~((!((8'haa) ? (~(8'hb6)) : ((8'hb6) ? (7'h43) : (8'hb1)))) ? {(((8'ha1) ? (8'hb4) : (8'h9c)) ? ((8'ha7) ^~ (8'ha2)) : ((8'had) ? (7'h40) : (8'hb4)))} : (-(^(8'ha4))))), 
parameter param395 = (((param394 ? param394 : ((param394 ? param394 : param394) - (8'ha4))) ? (|(~param394)) : param394) ? {(~&param394), ((~(param394 ? param394 : param394)) ~^ param394)} : (~&({(param394 ? param394 : (7'h43)), (&param394)} + (param394 * param394)))))
(y, clk, wire152, wire151, wire150, wire149, wire148);
  output wire [(32'hb8f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire152;
  input wire signed [(5'h12):(1'h0)] wire151;
  input wire [(3'h5):(1'h0)] wire150;
  input wire [(4'hb):(1'h0)] wire149;
  input wire [(4'hd):(1'h0)] wire148;
  wire signed [(5'h10):(1'h0)] wire393;
  wire [(2'h2):(1'h0)] wire392;
  wire signed [(2'h2):(1'h0)] wire391;
  wire [(5'h15):(1'h0)] wire390;
  wire [(3'h6):(1'h0)] wire389;
  wire [(3'h5):(1'h0)] wire153;
  reg signed [(4'hb):(1'h0)] reg387 = (1'h0);
  reg [(5'h13):(1'h0)] reg386 = (1'h0);
  reg [(5'h11):(1'h0)] reg385 = (1'h0);
  reg [(4'hd):(1'h0)] reg383 = (1'h0);
  reg [(5'h11):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg380 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg377 = (1'h0);
  reg [(3'h6):(1'h0)] reg376 = (1'h0);
  reg [(5'h14):(1'h0)] reg375 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg373 = (1'h0);
  reg [(4'h8):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg370 = (1'h0);
  reg [(4'hb):(1'h0)] reg367 = (1'h0);
  reg [(2'h2):(1'h0)] reg364 = (1'h0);
  reg [(4'hf):(1'h0)] reg362 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg361 = (1'h0);
  reg [(4'he):(1'h0)] reg360 = (1'h0);
  reg [(3'h6):(1'h0)] reg358 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg355 = (1'h0);
  reg [(4'h9):(1'h0)] reg354 = (1'h0);
  reg [(4'hb):(1'h0)] reg352 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg351 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg349 = (1'h0);
  reg [(4'he):(1'h0)] reg348 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg347 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg346 = (1'h0);
  reg [(4'h8):(1'h0)] reg345 = (1'h0);
  reg [(5'h10):(1'h0)] reg343 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg341 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg340 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg338 = (1'h0);
  reg [(4'hb):(1'h0)] reg337 = (1'h0);
  reg [(5'h13):(1'h0)] reg335 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg333 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg332 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg330 = (1'h0);
  reg [(5'h13):(1'h0)] reg329 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg328 = (1'h0);
  reg [(2'h3):(1'h0)] reg325 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg320 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg318 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg317 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg308 = (1'h0);
  reg [(5'h11):(1'h0)] reg307 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg306 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg305 = (1'h0);
  reg [(4'hf):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg302 = (1'h0);
  reg [(4'ha):(1'h0)] reg295 = (1'h0);
  reg [(5'h14):(1'h0)] reg294 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg293 = (1'h0);
  reg [(4'ha):(1'h0)] reg292 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg291 = (1'h0);
  reg [(2'h3):(1'h0)] reg286 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg283 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg279 = (1'h0);
  reg [(4'hd):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg276 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg275 = (1'h0);
  reg [(4'he):(1'h0)] reg274 = (1'h0);
  reg [(4'hd):(1'h0)] reg273 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg266 = (1'h0);
  reg [(3'h6):(1'h0)] reg265 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg262 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg260 = (1'h0);
  reg [(4'hc):(1'h0)] reg258 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg255 = (1'h0);
  reg [(3'h7):(1'h0)] reg254 = (1'h0);
  reg [(4'ha):(1'h0)] reg253 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg246 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg240 = (1'h0);
  reg [(2'h2):(1'h0)] reg252 = (1'h0);
  reg signed [(4'he):(1'h0)] reg249 = (1'h0);
  reg [(3'h4):(1'h0)] reg248 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg247 = (1'h0);
  reg [(5'h14):(1'h0)] reg244 = (1'h0);
  reg [(4'hc):(1'h0)] reg241 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg239 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg238 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg233 = (1'h0);
  reg [(2'h3):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg230 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg229 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg228 = (1'h0);
  reg [(3'h5):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg226 = (1'h0);
  reg [(3'h5):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg220 = (1'h0);
  reg [(4'ha):(1'h0)] reg216 = (1'h0);
  reg [(5'h12):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg213 = (1'h0);
  reg [(5'h10):(1'h0)] reg212 = (1'h0);
  reg [(4'ha):(1'h0)] reg211 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg210 = (1'h0);
  reg [(5'h11):(1'h0)] reg204 = (1'h0);
  reg [(4'hb):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg196 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg194 = (1'h0);
  reg [(3'h6):(1'h0)] reg192 = (1'h0);
  reg [(3'h7):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg188 = (1'h0);
  reg [(5'h12):(1'h0)] reg187 = (1'h0);
  reg [(5'h11):(1'h0)] reg186 = (1'h0);
  reg [(5'h12):(1'h0)] reg185 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg174 = (1'h0);
  reg [(4'hb):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg171 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg168 = (1'h0);
  reg [(5'h12):(1'h0)] reg167 = (1'h0);
  reg [(5'h12):(1'h0)] reg165 = (1'h0);
  reg [(4'hf):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg161 = (1'h0);
  reg [(4'ha):(1'h0)] reg160 = (1'h0);
  reg [(4'h9):(1'h0)] reg159 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg158 = (1'h0);
  reg [(4'he):(1'h0)] reg156 = (1'h0);
  reg [(3'h6):(1'h0)] reg155 = (1'h0);
  reg [(2'h2):(1'h0)] reg384 = (1'h0);
  reg [(4'hb):(1'h0)] reg378 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg388 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar384 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg381 = (1'h0);
  reg [(3'h4):(1'h0)] forvar378 = (1'h0);
  reg [(4'hb):(1'h0)] reg374 = (1'h0);
  reg [(3'h5):(1'h0)] reg372 = (1'h0);
  reg [(2'h2):(1'h0)] reg369 = (1'h0);
  reg [(5'h15):(1'h0)] forvar355 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg368 = (1'h0);
  reg [(4'hc):(1'h0)] reg366 = (1'h0);
  reg [(2'h3):(1'h0)] reg365 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg363 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg359 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg357 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg356 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar353 = (1'h0);
  reg signed [(4'he):(1'h0)] reg350 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg344 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg342 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg339 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg336 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar333 = (1'h0);
  reg [(4'he):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg331 = (1'h0);
  reg [(5'h14):(1'h0)] reg327 = (1'h0);
  reg [(2'h2):(1'h0)] reg326 = (1'h0);
  reg [(4'hb):(1'h0)] reg324 = (1'h0);
  reg [(5'h13):(1'h0)] reg323 = (1'h0);
  reg [(4'hb):(1'h0)] reg322 = (1'h0);
  reg [(4'h8):(1'h0)] forvar321 = (1'h0);
  reg [(4'ha):(1'h0)] reg319 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg316 = (1'h0);
  reg [(4'h9):(1'h0)] forvar313 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg312 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg311 = (1'h0);
  reg [(4'hd):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg309 = (1'h0);
  reg signed [(4'he):(1'h0)] reg303 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar287 = (1'h0);
  reg [(5'h12):(1'h0)] reg301 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg299 = (1'h0);
  reg [(4'hb):(1'h0)] reg298 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar297 = (1'h0);
  reg [(4'ha):(1'h0)] reg296 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg290 = (1'h0);
  reg [(5'h11):(1'h0)] reg289 = (1'h0);
  reg [(5'h10):(1'h0)] reg288 = (1'h0);
  reg [(4'he):(1'h0)] reg287 = (1'h0);
  reg [(5'h13):(1'h0)] reg285 = (1'h0);
  reg [(3'h7):(1'h0)] reg284 = (1'h0);
  reg [(4'h8):(1'h0)] reg282 = (1'h0);
  reg [(5'h11):(1'h0)] forvar260 = (1'h0);
  reg [(5'h12):(1'h0)] reg281 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg280 = (1'h0);
  reg [(4'ha):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg272 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg271 = (1'h0);
  reg [(3'h7):(1'h0)] reg269 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg268 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg267 = (1'h0);
  reg [(4'h9):(1'h0)] reg264 = (1'h0);
  reg [(3'h5):(1'h0)] reg261 = (1'h0);
  reg [(4'h9):(1'h0)] reg259 = (1'h0);
  reg [(5'h15):(1'h0)] reg257 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg250 = (1'h0);
  reg [(4'hc):(1'h0)] forvar242 = (1'h0);
  reg [(5'h15):(1'h0)] reg234 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg251 = (1'h0);
  reg [(5'h10):(1'h0)] forvar250 = (1'h0);
  reg [(3'h4):(1'h0)] forvar246 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg245 = (1'h0);
  reg [(4'h9):(1'h0)] reg243 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar240 = (1'h0);
  reg [(5'h10):(1'h0)] reg237 = (1'h0);
  reg [(3'h5):(1'h0)] reg236 = (1'h0);
  reg [(5'h13):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar234 = (1'h0);
  reg [(5'h11):(1'h0)] reg231 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg225 = (1'h0);
  reg [(5'h14):(1'h0)] reg223 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg222 = (1'h0);
  reg [(3'h6):(1'h0)] reg219 = (1'h0);
  reg [(4'he):(1'h0)] reg218 = (1'h0);
  reg [(2'h2):(1'h0)] reg217 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar214 = (1'h0);
  reg [(2'h3):(1'h0)] reg209 = (1'h0);
  reg [(5'h11):(1'h0)] reg208 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar207 = (1'h0);
  reg [(5'h10):(1'h0)] reg206 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg205 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg202 = (1'h0);
  reg [(4'h9):(1'h0)] reg201 = (1'h0);
  reg [(3'h5):(1'h0)] forvar194 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg197 = (1'h0);
  reg [(5'h10):(1'h0)] reg195 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg193 = (1'h0);
  reg [(5'h13):(1'h0)] reg190 = (1'h0);
  reg [(4'hf):(1'h0)] reg189 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar180 = (1'h0);
  reg [(5'h10):(1'h0)] forvar178 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg176 = (1'h0);
  reg [(3'h7):(1'h0)] reg175 = (1'h0);
  reg [(4'hc):(1'h0)] forvar173 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg166 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg170 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg169 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar166 = (1'h0);
  reg [(4'hb):(1'h0)] reg163 = (1'h0);
  reg [(4'hc):(1'h0)] reg162 = (1'h0);
  reg [(4'h8):(1'h0)] reg157 = (1'h0);
  reg [(4'ha):(1'h0)] reg154 = (1'h0);
  assign y = {reg258,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg246,
                 reg240,
                 reg252,
                 reg249,
                 reg248,
                 reg247,
                 reg244,
                 reg241,
                 reg239,
                 reg238,
                 reg233,
                 reg232,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg224,
                 reg221,
                 reg220,
                 reg216,
                 reg215,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg204,
                 reg200,
                 reg199,
                 reg198,
                 reg196,
                 reg194,
                 reg192,
                 reg191,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg182,
                 reg179,
                 reg174,
                 reg172,
                 reg171,
                 reg168,
                 reg167,
                 reg165,
                 reg164,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg156,
                 reg155,
                 reg384,
                 reg378,
                 reg388,
                 forvar384,
                 reg381,
                 forvar378,
                 reg374,
                 reg372,
                 reg369,
                 forvar355,
                 reg368,
                 reg366,
                 reg365,
                 reg363,
                 reg359,
                 reg357,
                 reg356,
                 forvar353,
                 reg350,
                 reg344,
                 reg342,
                 reg339,
                 reg336,
                 forvar333,
                 reg334,
                 reg331,
                 reg327,
                 reg326,
                 reg324,
                 reg323,
                 reg322,
                 forvar321,
                 reg319,
                 reg316,
                 forvar313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg303,
                 reg297,
                 forvar287,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 forvar297,
                 reg296,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg285,
                 reg284,
                 reg282,
                 forvar260,
                 reg281,
                 reg280,
                 reg277,
                 reg272,
                 reg271,
                 reg269,
                 reg268,
                 reg267,
                 reg264,
                 reg261,
                 reg259,
                 reg257,
                 reg250,
                 forvar242,
                 reg234,
                 reg251,
                 forvar250,
                 forvar246,
                 reg245,
                 reg243,
                 reg242,
                 forvar240,
                 reg237,
                 reg236,
                 reg235,
                 forvar234,
                 reg231,
                 reg225,
                 reg223,
                 reg222,
                 reg219,
                 reg218,
                 reg217,
                 forvar214,
                 reg209,
                 reg208,
                 forvar207,
                 reg206,
                 reg205,
                 reg203,
                 reg202,
                 reg201,
                 forvar194,
                 reg197,
                 reg195,
                 reg193,
                 reg190,
                 reg189,
                 reg184,
                 reg183,
                 reg181,
                 forvar180,
                 forvar178,
                 reg177,
                 reg176,
                 reg175,
                 forvar173,
                 reg166,
                 reg170,
                 reg169,
                 forvar166,
                 reg163,
                 reg162,
                 reg157,
                 reg154,
                 (1'h0)};
  assign wire153 = ({wire150[(1'h0):(1'h0)]} && wire149);
  always
    @(posedge clk) begin
      if (($unsigned((8'haf)) ^~ $unsigned($unsigned((~&$signed(wire152))))))
        begin
          reg154 = (!$signed($signed({{wire151, wire151},
              ((8'ha1) || (8'ha1))})));
          if ($signed((8'hb5)))
            begin
              reg155 <= ($unsigned($signed(wire148)) < ($signed(wire152) && $unsigned((~wire149))));
              reg156 <= $signed(wire149);
            end
          else
            begin
              reg157 = (reg156[(2'h2):(1'h0)] << $unsigned({{(~&(8'hb8))},
                  wire153[(1'h0):(1'h0)]}));
              reg158 <= (|{(~&$unsigned(reg157)),
                  (-$signed($unsigned(wire149)))});
              reg159 <= reg156[(4'h8):(3'h5)];
              reg160 <= {(8'hbe)};
            end
          if (wire150)
            begin
              reg161 <= {wire153[(2'h2):(1'h0)],
                  {((((8'hbf) && wire152) ?
                              $signed((8'ha7)) : reg159[(2'h3):(1'h0)]) ?
                          $unsigned((-reg154)) : $signed($unsigned(reg159)))}};
            end
          else
            begin
              reg161 <= reg156;
              reg162 = wire151;
              reg163 = (^~(reg156[(3'h4):(2'h3)] == ({((8'hb3) ?
                          reg154 : reg154),
                      $unsigned(reg161)} ?
                  $signed((wire152 ?
                      (8'had) : reg162)) : {((8'ha6) + reg159)})));
              reg164 <= (8'hb5);
              reg165 <= reg158;
            end
          for (forvar166 = (1'h0); (forvar166 < (1'h0)); forvar166 = (forvar166 + (1'h1)))
            begin
              reg167 <= {$unsigned(reg165),
                  (~(~|($unsigned(wire149) ?
                      (wire148 < (8'haa)) : (reg156 ^ reg159))))};
              reg168 <= {{{(~^(reg155 >= (8'hac))), (8'ha1)}}};
              reg169 = ((8'hb2) & wire153[(2'h3):(2'h2)]);
            end
          reg170 = $signed({{$unsigned((!reg156)), reg158[(4'h9):(3'h5)]}});
        end
      else
        begin
          if (reg156[(2'h3):(2'h2)])
            begin
              reg155 <= ((|(((wire149 ?
                      reg163 : reg156) - (8'hb0)) + (7'h40))) ?
                  $unsigned(wire152[(4'hf):(4'h8)]) : $signed({{(forvar166 > reg154)},
                      (wire148 + (reg154 ? forvar166 : reg167))}));
              reg156 <= reg157;
              reg158 <= (reg156[(1'h0):(1'h0)] ?
                  ((&{$unsigned(reg156)}) ?
                      ($unsigned($unsigned(wire153)) <<< reg163) : (($unsigned(wire153) << $unsigned(reg170)) ?
                          ({reg162} | reg160[(4'h8):(3'h5)]) : ((8'hb6) ?
                              {reg168, reg158} : $signed(reg162)))) : reg164);
              reg159 <= (-reg160[(3'h5):(2'h2)]);
            end
          else
            begin
              reg154 = $unsigned((-wire152[(5'h13):(4'hd)]));
              reg157 = reg164;
              reg158 <= reg155;
              reg159 <= $signed($signed($unsigned(((reg163 ?
                  reg168 : wire151) ^~ (reg168 + reg160)))));
              reg160 <= $unsigned(reg168[(2'h2):(2'h2)]);
            end
          if (reg156)
            begin
              reg161 <= (|$unsigned({{(wire148 ? (8'hb4) : wire152), reg158},
                  $signed(wire153)}));
            end
          else
            begin
              reg162 = $signed($signed(reg157));
              reg163 = (!(reg161 ?
                  $signed($signed($unsigned(reg159))) : reg161));
            end
          if (wire151[(4'hf):(4'h9)])
            begin
              reg166 = reg154;
              reg167 <= wire148;
              reg168 <= reg162;
            end
          else
            begin
              reg166 = $signed({(reg158[(2'h3):(1'h1)] ?
                      reg163[(1'h1):(1'h1)] : {(reg163 + reg170)})});
              reg169 = ($unsigned(({$unsigned((8'ha4)),
                  {reg163}} & $unsigned($signed(wire149)))) << (~&($unsigned($unsigned(reg169)) ?
                  $unsigned(reg157[(3'h6):(3'h5)]) : $signed($unsigned(forvar166)))));
              reg170 = ({$unsigned($signed((wire150 ? wire149 : reg158))),
                      $unsigned(((reg162 ? wire152 : reg168) ?
                          wire150 : $signed(reg168)))} ?
                  reg161[(4'he):(4'ha)] : reg161);
              reg171 <= reg164[(3'h6):(3'h4)];
            end
          reg172 <= (($signed(((8'hba) ?
                  (wire151 ? reg168 : reg155) : ((8'hbf) ? reg166 : reg165))) ?
              {$unsigned((reg158 ? (8'ha0) : reg158))} : (reg160 ?
                  $signed($unsigned(wire151)) : $unsigned(wire153[(1'h0):(1'h0)]))) - ((^~($signed(wire150) ?
              (reg155 ? reg167 : reg154) : (reg164 ?
                  (8'hab) : reg169))) >= (^reg159)));
          for (forvar173 = (1'h0); (forvar173 < (2'h2)); forvar173 = (forvar173 + (1'h1)))
            begin
              reg174 <= (wire150[(1'h1):(1'h0)] || (~^$signed(((~^reg161) >>> (-reg160)))));
              reg175 = wire150;
              reg176 = $signed(reg171[(4'ha):(1'h0)]);
              reg177 = ((~^(8'hb2)) ?
                  (reg162 ?
                      $unsigned(wire153[(2'h2):(1'h0)]) : reg161) : (|({$signed(reg170)} >= {reg167})));
            end
        end
      for (forvar178 = (1'h0); (forvar178 < (2'h3)); forvar178 = (forvar178 + (1'h1)))
        begin
          reg179 <= reg162[(4'hb):(1'h1)];
          for (forvar180 = (1'h0); (forvar180 < (1'h1)); forvar180 = (forvar180 + (1'h1)))
            begin
              reg181 = ($unsigned(forvar166) ?
                  wire151 : (($signed(((8'ha5) == forvar173)) | (~reg157[(2'h3):(1'h1)])) - $signed($signed(((8'hb6) ?
                      (8'ha8) : reg159)))));
              reg182 <= {($unsigned(({reg162, reg176} ?
                      ((8'ha2) | reg160) : reg156)) >> (^{reg163,
                      $unsigned(reg166)}))};
            end
          if ($signed({(+($unsigned(reg172) ?
                  (reg174 ? reg154 : (8'hb4)) : (&(8'hac)))),
              $signed($unsigned({reg170}))}))
            begin
              reg183 = $unsigned(reg158);
              reg184 = ((8'hbc) ?
                  $unsigned($signed($signed({wire152}))) : $unsigned((-reg174[(2'h2):(1'h1)])));
            end
          else
            begin
              reg185 <= (wire152 <<< ({((reg181 * forvar173) || reg170)} ?
                  $unsigned(({reg165,
                      reg175} * wire153[(3'h4):(3'h4)])) : (8'ha3)));
              reg186 <= (~|$unsigned(((&(reg156 ?
                  (8'ha9) : reg168)) | reg169[(3'h6):(3'h6)])));
              reg187 <= (forvar178[(4'he):(4'h9)] != wire151[(1'h1):(1'h0)]);
              reg188 <= $unsigned(reg163[(4'h8):(3'h6)]);
            end
          if ((~&($signed(((reg181 + reg187) ?
              (forvar173 <<< (8'ha9)) : (reg188 ~^ forvar166))) <<< (^reg187[(3'h5):(1'h0)]))))
            begin
              reg189 = $unsigned((reg177[(1'h1):(1'h1)] ?
                  (reg181 ?
                      {$unsigned(forvar173)} : ((reg176 ?
                          (8'hbe) : wire151) >> reg157)) : reg171));
              reg190 = (($signed($signed($signed(reg162))) ^~ {(8'h9e)}) ^~ forvar166[(1'h0):(1'h0)]);
            end
          else
            begin
              reg189 = {{$unsigned(reg163),
                      $signed(($signed(reg170) ^~ reg170))},
                  ($unsigned({(reg156 ?
                          (8'h9c) : (8'hb3))}) ~^ ((~(|reg175)) ^~ (~&(reg177 ?
                      (7'h43) : reg170))))};
              reg190 = (~^{$unsigned($unsigned((wire149 <= reg184)))});
              reg191 <= ((^~(&$unsigned($unsigned(reg182)))) <<< ((^((wire149 ?
                      reg161 : forvar178) >> wire148)) ?
                  reg174 : forvar178[(1'h1):(1'h0)]));
              reg192 <= {({reg163, {reg184, {reg156, reg164}}} ?
                      (((wire149 ? reg162 : reg165) ?
                              (reg175 ? (8'ha0) : reg177) : (|reg172)) ?
                          reg166[(2'h2):(2'h2)] : $signed(reg157[(3'h6):(2'h3)])) : reg171[(4'hd):(2'h2)])};
            end
          reg193 = $unsigned(reg172[(3'h4):(2'h3)]);
        end
      if ({reg163[(4'h9):(2'h2)],
          $signed(((~reg163) ?
              ($unsigned(reg159) ?
                  ((8'h9c) ? reg161 : (8'hb2)) : (^reg183)) : reg166))})
        begin
          if (reg165[(1'h1):(1'h1)])
            begin
              reg194 <= (^~reg186[(1'h1):(1'h0)]);
              reg195 = $signed(reg189[(4'he):(4'hc)]);
              reg196 <= forvar178[(3'h4):(1'h0)];
              reg197 = (($signed((|reg183)) ?
                  $unsigned(reg166[(4'hd):(1'h1)]) : $signed(($unsigned(reg155) ?
                      {reg169} : reg175))) >>> ($unsigned((&(reg162 - reg185))) ?
                  $unsigned(wire151) : (reg177 << $signed($signed(reg196)))));
              reg198 <= reg156[(4'ha):(4'h8)];
            end
          else
            begin
              reg195 = $unsigned(((-($unsigned(reg187) ^ (~|wire151))) > (reg186 << {{reg196,
                      reg182},
                  (8'hbd)})));
              reg196 <= {$unsigned((~|$unsigned(reg195[(2'h2):(1'h0)])))};
            end
        end
      else
        begin
          for (forvar194 = (1'h0); (forvar194 < (2'h2)); forvar194 = (forvar194 + (1'h1)))
            begin
              reg196 <= ($unsigned((reg171[(2'h3):(1'h1)] ^~ ($unsigned(reg171) ?
                  (|reg156) : forvar180))) * (|((~^(reg193 >> wire149)) == (^~{(8'ha2),
                  (8'ha3)}))));
              reg197 = (+(reg187[(3'h4):(2'h3)] ^~ (+reg189[(4'hb):(1'h1)])));
            end
          if ($signed((wire149 ?
              ($unsigned(reg167[(4'hf):(4'h9)]) ?
                  ((reg185 <= reg168) ?
                      $signed(reg179) : reg176[(2'h2):(2'h2)]) : $signed($signed(reg179))) : ($unsigned($unsigned(reg162)) <<< $unsigned({reg156,
                  reg191})))))
            begin
              reg198 <= (&($signed({$signed(reg155)}) ?
                  {reg182[(3'h7):(3'h4)],
                      $signed(((7'h42) ?
                          reg169 : forvar166))} : reg158[(3'h6):(3'h6)]));
              reg199 <= reg175[(3'h7):(3'h5)];
              reg200 <= $signed({$unsigned(((reg181 * reg172) != $signed(wire149))),
                  $signed($signed(reg187[(1'h0):(1'h0)]))});
              reg201 = ($signed((~((reg197 == reg195) ?
                      $signed(reg198) : (wire150 ? reg181 : reg159)))) ?
                  {($signed($unsigned(reg177)) ?
                          $unsigned({reg171}) : forvar173),
                      reg196[(4'ha):(1'h1)]} : ((^reg163) * (((reg165 ?
                          wire153 : reg179) ?
                      reg162[(2'h2):(2'h2)] : $signed(reg156)) && $unsigned(reg159))));
            end
          else
            begin
              reg201 = {({reg193} ? $signed(reg191) : reg184[(1'h1):(1'h1)])};
              reg202 = (&forvar178[(3'h6):(3'h4)]);
              reg203 = ({(~(~|(reg172 ? reg198 : (8'hab))))} ?
                  (7'h41) : (~&(reg182 ^ (8'hab))));
            end
          if ($signed($unsigned($signed(($unsigned(reg184) >= $signed(forvar180))))))
            begin
              reg204 <= ($signed((reg184[(2'h2):(1'h1)] ?
                      wire150 : $unsigned(reg201[(3'h5):(2'h2)]))) ?
                  $unsigned(reg199[(4'h9):(4'h8)]) : $signed((((reg160 ?
                              reg159 : (8'hb4)) ?
                          (reg181 ? reg202 : reg187) : $unsigned(reg193)) ?
                      $unsigned((reg156 << forvar173)) : wire152[(5'h12):(4'hb)])));
              reg205 = $unsigned((reg203[(3'h6):(1'h0)] != ((^(reg163 ?
                      reg196 : reg186)) ?
                  ((reg167 || reg181) * (reg179 <<< reg157)) : $unsigned($unsigned((7'h41))))));
              reg206 = $unsigned((reg157 || $signed($signed($signed(reg197)))));
            end
          else
            begin
              reg204 <= reg154[(4'ha):(3'h5)];
            end
          for (forvar207 = (1'h0); (forvar207 < (3'h4)); forvar207 = (forvar207 + (1'h1)))
            begin
              reg208 = reg161[(5'h11):(5'h10)];
              reg209 = ((reg183[(4'ha):(2'h2)] ^ (&$signed(reg203[(4'hb):(4'ha)]))) - reg192);
              reg210 <= {(({$unsigned(reg156), $unsigned(reg176)} ?
                          $unsigned($signed(reg177)) : $unsigned((|reg198))) ?
                      ($unsigned((reg169 & wire150)) ?
                          $unsigned($unsigned(reg169)) : {reg205[(2'h3):(2'h2)]}) : ($unsigned((reg176 ?
                          reg182 : reg187)) > reg197[(4'h9):(1'h1)]))};
              reg211 <= ($unsigned((~|$signed(reg172[(3'h5):(1'h1)]))) ?
                  $unsigned((reg162 ^ (&{reg164,
                      (8'ha3)}))) : reg176[(1'h1):(1'h0)]);
              reg212 <= reg199;
            end
          reg213 <= reg169[(1'h0):(1'h0)];
        end
      for (forvar214 = (1'h0); (forvar214 < (2'h3)); forvar214 = (forvar214 + (1'h1)))
        begin
          reg215 <= (^~(8'ha2));
          reg216 <= reg211[(2'h2):(1'h1)];
          if ((~((~$unsigned((reg185 == (8'ha6)))) && reg181)))
            begin
              reg217 = $unsigned($signed(wire149));
            end
          else
            begin
              reg217 = ($signed(reg187) ?
                  (8'hba) : $unsigned(reg204[(4'h9):(3'h4)]));
              reg218 = reg195;
              reg219 = reg156;
              reg220 <= (!reg162);
              reg221 <= (($unsigned(((8'hae) >> $signed(reg185))) ~^ (forvar173[(3'h7):(3'h6)] ^ $unsigned((wire149 ?
                  reg166 : (8'h9e))))) > ($signed(reg161) ?
                  {((-reg161) < (forvar214 & reg216)),
                      $signed(reg211)} : (~|$unsigned($unsigned(wire149)))));
            end
          if ($unsigned($unsigned(($unsigned((reg208 <<< reg155)) | ({forvar173} ~^ {wire153,
              reg192})))))
            begin
              reg222 = forvar173[(4'hb):(3'h5)];
              reg223 = reg186[(4'hb):(3'h5)];
            end
          else
            begin
              reg222 = reg223;
              reg224 <= (reg165[(4'hd):(4'ha)] ^~ reg163[(4'hb):(4'ha)]);
              reg225 = $unsigned(((^(8'h9f)) ~^ reg177[(2'h2):(1'h1)]));
              reg226 <= reg188;
            end
          if (((8'hb5) ?
              {{$unsigned(((8'hab) >>> reg225))}} : ($signed($signed((^~wire153))) ^~ ($unsigned($unsigned(forvar166)) && reg196))))
            begin
              reg227 <= ({wire148[(4'h8):(2'h2)],
                  (($unsigned(reg167) <<< reg191) ^ $unsigned((7'h42)))} != $unsigned((((forvar178 ~^ reg161) < (reg223 >>> reg182)) ?
                  (^(reg199 | reg200)) : $signed({reg190, reg195}))));
              reg228 <= $signed({$unsigned((reg196[(3'h4):(3'h4)] ?
                      $unsigned(reg186) : $signed(forvar173))),
                  reg155[(2'h3):(2'h2)]});
              reg229 <= $signed(reg221);
              reg230 <= $unsigned($unsigned(reg202[(3'h7):(3'h7)]));
              reg231 = (8'ha6);
            end
          else
            begin
              reg227 <= reg193;
              reg231 = (|(reg222 & $unsigned((+((8'hb2) ? reg224 : reg204)))));
              reg232 <= reg189;
              reg233 <= {((&$unsigned(reg219[(3'h4):(3'h4)])) >> $unsigned($signed(reg158))),
                  $signed(reg232[(1'h1):(1'h0)])};
            end
        end
      if (((~&$signed((-(~|reg225)))) ?
          ($signed(reg166) ?
              (reg154[(1'h0):(1'h0)] == ({(8'h9f),
                  reg210} <= (reg193 >>> (8'h9c)))) : (reg219 ?
                  (((8'haf) ?
                      reg176 : (8'ha2)) <= $signed((8'haa))) : (~|{reg205,
                      reg232}))) : $signed((~|($unsigned(reg167) ?
              (reg210 ? reg210 : wire152) : reg222)))))
        begin
          for (forvar234 = (1'h0); (forvar234 < (3'h4)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 = ({$unsigned(($unsigned((8'hb0)) ?
                      wire149 : (~|reg217)))} >> $signed($unsigned(($unsigned((7'h44)) || reg204[(3'h7):(3'h4)]))));
              reg236 = (+reg159);
              reg237 = $unsigned(($unsigned((reg169[(4'h9):(1'h0)] ^~ (reg211 ^~ forvar178))) ?
                  reg228[(1'h0):(1'h0)] : ((~|reg194) ?
                      $unsigned((reg199 ? (7'h44) : reg202)) : (8'had))));
              reg238 <= ((!$unsigned((reg163 ?
                  $unsigned(reg172) : (reg221 && reg184)))) <<< $signed(reg157));
              reg239 <= reg222;
            end
          for (forvar240 = (1'h0); (forvar240 < (1'h1)); forvar240 = (forvar240 + (1'h1)))
            begin
              reg241 <= $unsigned((&reg237[(2'h2):(1'h1)]));
              reg242 = ((forvar178 >= $unsigned($unsigned((~&reg204)))) ?
                  $unsigned((+reg212)) : (reg175[(1'h0):(1'h0)] ?
                      reg227[(1'h0):(1'h0)] : (forvar240 ?
                          $signed(reg155) : reg199)));
              reg243 = ((~$signed($signed((8'ha5)))) ?
                  (+$unsigned(({reg183, reg159} ?
                      (reg236 ?
                          reg184 : (8'ha7)) : (!(8'ha9))))) : $unsigned($unsigned(reg209[(1'h0):(1'h0)])));
              reg244 <= $signed({$unsigned((-$unsigned(reg176)))});
              reg245 = $unsigned((8'hbe));
            end
          for (forvar246 = (1'h0); (forvar246 < (3'h4)); forvar246 = (forvar246 + (1'h1)))
            begin
              reg247 <= ((reg194 <= reg237[(4'ha):(3'h6)]) == (((~&(reg198 >> reg167)) + reg213) ?
                  $signed(reg219) : wire152));
              reg248 <= ($signed(wire151[(5'h12):(4'hf)]) ~^ reg211);
              reg249 <= reg232;
            end
          for (forvar250 = (1'h0); (forvar250 < (2'h2)); forvar250 = (forvar250 + (1'h1)))
            begin
              reg251 = ({(^~reg242[(3'h7):(2'h2)])} ^~ (+reg229[(1'h0):(1'h0)]));
              reg252 <= $unsigned(({$unsigned($signed((8'hbe))),
                      reg164[(4'hf):(3'h5)]} ?
                  $signed(($unsigned(reg216) ?
                      (reg157 ?
                          reg245 : reg181) : $signed(reg223))) : (+$unsigned((!(8'ha9))))));
            end
        end
      else
        begin
          if ($unsigned(((reg241[(4'hc):(4'h9)] ?
                  ($unsigned(reg191) + (reg239 ?
                      reg252 : (8'had))) : $signed($signed(reg179))) ?
              {((reg235 ? reg157 : (8'hbc)) <= $signed(reg168)),
                  $signed(((8'ha6) | reg202))} : reg199)))
            begin
              reg234 = reg205[(3'h5):(3'h4)];
              reg238 <= ((|(&$unsigned($unsigned(reg251)))) ?
                  reg201[(3'h5):(3'h4)] : (-((reg193[(3'h6):(2'h3)] ?
                          (^~reg155) : $signed((8'ha2))) ?
                      ($unsigned(reg233) & $unsigned((8'hbc))) : $unsigned($signed(reg196)))));
            end
          else
            begin
              reg238 <= ($unsigned(((|$unsigned(reg160)) ?
                      $unsigned($unsigned(wire152)) : $signed((reg208 | reg186)))) ?
                  reg242 : (reg249 << $signed(($signed(reg234) >> $unsigned((8'hb0))))));
              reg239 <= reg206[(2'h2):(2'h2)];
              reg240 <= ((!{$unsigned(wire152[(2'h3):(2'h3)])}) ^ (-(|{reg186,
                  $unsigned(reg243)})));
              reg241 <= {$unsigned(reg233), $signed(reg240)};
            end
          for (forvar242 = (1'h0); (forvar242 < (2'h3)); forvar242 = (forvar242 + (1'h1)))
            begin
              reg244 <= $unsigned($signed(reg238[(1'h1):(1'h0)]));
              reg245 = ((&{$unsigned(reg228[(4'h9):(4'h8)]),
                  ($unsigned(reg176) || $unsigned(reg204))}) | ($unsigned((reg179 ?
                      $signed(reg186) : (wire153 ? reg216 : reg229))) ?
                  $signed($unsigned($signed(reg194))) : reg240[(2'h2):(1'h0)]));
              reg246 <= $signed(reg251[(1'h1):(1'h1)]);
              reg250 = forvar234;
            end
          if (reg249[(4'ha):(4'h9)])
            begin
              reg251 = {reg219, reg252};
              reg252 <= reg198[(2'h2):(1'h0)];
              reg253 <= (reg177[(2'h3):(2'h2)] ^ $unsigned((~&(+reg177[(3'h4):(2'h3)]))));
            end
          else
            begin
              reg251 = wire151[(3'h7):(3'h5)];
              reg252 <= (^(~|(&$unsigned($unsigned(reg166)))));
              reg253 <= (forvar250[(4'hc):(4'ha)] ~^ ({(((8'hbf) ?
                      reg198 : reg205) < reg199[(4'h8):(3'h5)])} >> reg209[(2'h2):(2'h2)]));
            end
          if ((reg248[(1'h0):(1'h0)] || ($signed(reg250) ?
              (reg246 >> {(reg213 != reg165)}) : $unsigned((reg203 ?
                  {reg250, reg192} : (!reg183))))))
            begin
              reg254 <= (reg193 ? reg252[(1'h1):(1'h1)] : reg211);
              reg255 <= $unsigned({$unsigned((reg228[(1'h1):(1'h1)] * $unsigned(wire149)))});
            end
          else
            begin
              reg254 <= reg177;
            end
          if ((reg239 ?
              $unsigned($signed((&$signed(reg253)))) : ($unsigned($unsigned($signed(reg221))) ~^ $unsigned(($signed(reg243) ?
                  (8'hb1) : forvar173[(3'h5):(1'h0)])))))
            begin
              reg256 <= (-{{$unsigned(((8'had) ? reg195 : reg170)),
                      ($signed((8'haa)) ?
                          $unsigned(reg164) : reg195[(4'h8):(3'h5)])}});
              reg257 = ($unsigned($unsigned((forvar240[(3'h5):(3'h4)] != (reg219 == reg254)))) > $signed($unsigned((~reg177))));
              reg258 <= reg222[(1'h1):(1'h0)];
              reg259 = $unsigned($unsigned(reg232));
            end
          else
            begin
              reg256 <= (((+(~^$unsigned(reg247))) || $signed((!(8'hae)))) ?
                  ($unsigned($signed((reg188 ? reg232 : reg255))) ?
                      $unsigned(reg242) : (~{(|(8'ha5)),
                          $unsigned(reg202)})) : (!$unsigned(((~&reg169) ?
                      $signed(reg243) : reg256[(4'h8):(4'h8)]))));
              reg257 = $signed($unsigned((8'haf)));
            end
        end
    end
endmodule
