(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param1136 = {{(&(^(7'h40)))}, {(((7'h44) ^~ (~&(7'h46))) && (|{(7'h49), (8'ha4)}))}}, 
parameter param1137 = ({{param1136}, (((param1136 ^~ param1136) * (&(7'h40))) ^~ param1136)} ? param1136 : (8'hb4)))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h7c1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h18):(1'h0)] wire3;
  input wire [(2'h2):(1'h0)] wire2;
  input wire signed [(5'h18):(1'h0)] wire1;
  input wire [(5'h11):(1'h0)] wire0;
  wire signed [(5'h17):(1'h0)] wire1092;
  wire signed [(5'h12):(1'h0)] wire1090;
  wire [(4'hf):(1'h0)] wire1089;
  wire [(4'hd):(1'h0)] wire1088;
  wire signed [(5'h18):(1'h0)] wire1064;
  wire [(4'hc):(1'h0)] wire1063;
  wire [(5'h13):(1'h0)] wire1028;
  wire signed [(5'h11):(1'h0)] wire1030;
  wire signed [(5'h14):(1'h0)] wire1031;
  wire [(2'h2):(1'h0)] wire1032;
  reg [(3'h7):(1'h0)] reg1135 = (1'h0);
  reg [(3'h7):(1'h0)] reg1127 = (1'h0);
  reg [(5'h10):(1'h0)] reg1129 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1128 = (1'h0);
  reg [(4'hd):(1'h0)] reg1123 = (1'h0);
  reg [(5'h18):(1'h0)] reg1122 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1121 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1120 = (1'h0);
  reg [(5'h10):(1'h0)] reg1118 = (1'h0);
  reg [(5'h10):(1'h0)] reg1112 = (1'h0);
  reg [(5'h17):(1'h0)] reg1109 = (1'h0);
  reg [(3'h5):(1'h0)] reg1107 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1106 = (1'h0);
  reg [(5'h14):(1'h0)] reg1103 = (1'h0);
  reg [(4'ha):(1'h0)] reg1102 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1100 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1099 = (1'h0);
  reg [(2'h3):(1'h0)] reg1097 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1095 = (1'h0);
  reg [(5'h13):(1'h0)] reg1091 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1086 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1085 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1083 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1082 = (1'h0);
  reg [(4'ha):(1'h0)] reg1081 = (1'h0);
  reg [(5'h16):(1'h0)] reg1080 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1076 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1072 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1071 = (1'h0);
  reg [(5'h18):(1'h0)] reg1070 = (1'h0);
  reg [(5'h12):(1'h0)] reg1069 = (1'h0);
  reg [(3'h4):(1'h0)] reg1067 = (1'h0);
  reg [(5'h13):(1'h0)] reg1066 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1061 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1060 = (1'h0);
  reg [(5'h17):(1'h0)] reg1059 = (1'h0);
  reg [(4'ha):(1'h0)] reg1057 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1055 = (1'h0);
  reg [(5'h11):(1'h0)] reg1054 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1050 = (1'h0);
  reg [(5'h10):(1'h0)] reg1045 = (1'h0);
  reg [(4'hc):(1'h0)] reg1047 = (1'h0);
  reg [(3'h5):(1'h0)] reg1046 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1042 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1038 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1037 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg34 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg33 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg32 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg28 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg27 = (1'h0);
  reg [(5'h12):(1'h0)] reg25 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg24 = (1'h0);
  reg [(4'hf):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg21 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg20 = (1'h0);
  reg [(4'ha):(1'h0)] reg19 = (1'h0);
  reg [(2'h3):(1'h0)] reg12 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg9 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1134 = (1'h0);
  reg [(4'h8):(1'h0)] reg1133 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1132 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1131 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1130 = (1'h0);
  reg [(5'h16):(1'h0)] reg1117 = (1'h0);
  reg [(4'he):(1'h0)] forvar1127 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1126 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1125 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1124 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1119 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1117 = (1'h0);
  reg [(4'ha):(1'h0)] reg1116 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1115 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1114 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1113 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1111 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1110 = (1'h0);
  reg [(3'h4):(1'h0)] reg1108 = (1'h0);
  reg [(4'he):(1'h0)] reg1105 = (1'h0);
  reg [(3'h7):(1'h0)] reg1104 = (1'h0);
  reg [(5'h11):(1'h0)] reg1101 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1098 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1094 = (1'h0);
  reg [(5'h16):(1'h0)] reg1093 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1087 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1084 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1079 = (1'h0);
  reg [(4'hb):(1'h0)] reg1078 = (1'h0);
  reg [(5'h12):(1'h0)] reg1077 = (1'h0);
  reg [(5'h10):(1'h0)] reg1075 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1074 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1073 = (1'h0);
  reg [(2'h3):(1'h0)] reg1068 = (1'h0);
  reg [(2'h2):(1'h0)] reg1065 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1062 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1058 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1056 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1053 = (1'h0);
  reg [(3'h7):(1'h0)] reg1052 = (1'h0);
  reg [(4'hc):(1'h0)] reg1051 = (1'h0);
  reg [(4'hd):(1'h0)] reg1049 = (1'h0);
  reg [(5'h16):(1'h0)] reg1048 = (1'h0);
  reg [(5'h16):(1'h0)] reg1043 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1045 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1044 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1043 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1041 = (1'h0);
  reg [(2'h2):(1'h0)] reg1040 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1039 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1036 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1035 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1034 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar31 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg29 = (1'h0);
  reg [(4'h9):(1'h0)] forvar26 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg22 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar21 = (1'h0);
  reg [(4'hd):(1'h0)] forvar10 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg18 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg17 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar14 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg13 = (1'h0);
  reg signed [(4'he):(1'h0)] reg11 = (1'h0);
  reg [(5'h15):(1'h0)] reg10 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4 = (1'h0);
  assign y = {wire1092,
                 wire1090,
                 wire1089,
                 wire1088,
                 wire1064,
                 wire1063,
                 wire1028,
                 wire1030,
                 wire1031,
                 wire1032,
                 reg1135,
                 reg1127,
                 reg1129,
                 reg1128,
                 reg1123,
                 reg1122,
                 reg1121,
                 reg1120,
                 reg1118,
                 reg1112,
                 reg1109,
                 reg1107,
                 reg1106,
                 reg1103,
                 reg1102,
                 reg1100,
                 reg1099,
                 reg1097,
                 reg1096,
                 reg1095,
                 reg1091,
                 reg1086,
                 reg1085,
                 reg1083,
                 reg1082,
                 reg1081,
                 reg1080,
                 reg1076,
                 reg1072,
                 reg1071,
                 reg1070,
                 reg1069,
                 reg1067,
                 reg1066,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1057,
                 reg1055,
                 reg1054,
                 reg1050,
                 reg1045,
                 reg1047,
                 reg1046,
                 reg1042,
                 reg1038,
                 reg1037,
                 reg34,
                 reg33,
                 reg32,
                 reg30,
                 reg28,
                 reg27,
                 reg25,
                 reg24,
                 reg14,
                 reg21,
                 reg20,
                 reg19,
                 reg12,
                 reg9,
                 reg8,
                 reg7,
                 reg5,
                 forvar1134,
                 reg1133,
                 forvar1132,
                 reg1131,
                 forvar1130,
                 reg1117,
                 forvar1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1119,
                 forvar1117,
                 reg1116,
                 reg1115,
                 reg1114,
                 reg1113,
                 forvar1111,
                 reg1110,
                 reg1108,
                 reg1105,
                 reg1104,
                 reg1101,
                 reg1098,
                 forvar1094,
                 reg1093,
                 reg1087,
                 reg1084,
                 forvar1079,
                 reg1078,
                 reg1077,
                 reg1075,
                 reg1074,
                 reg1073,
                 reg1068,
                 reg1065,
                 reg1062,
                 reg1058,
                 reg1056,
                 reg1053,
                 reg1052,
                 reg1051,
                 reg1049,
                 reg1048,
                 reg1043,
                 forvar1045,
                 reg1044,
                 forvar1043,
                 reg1041,
                 reg1040,
                 reg1039,
                 reg1036,
                 forvar1035,
                 reg1034,
                 forvar31,
                 reg29,
                 forvar26,
                 reg23,
                 reg22,
                 forvar21,
                 forvar10,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 forvar14,
                 reg13,
                 reg11,
                 reg10,
                 forvar6,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (2'h3)); forvar4 = (forvar4 + (1'h1)))
        begin
          reg5 <= wire3;
        end
      for (forvar6 = (1'h0); (forvar6 < (2'h3)); forvar6 = (forvar6 + (1'h1)))
        begin
          if ((8'hbc))
            begin
              reg7 <= (wire1 == forvar6);
              reg8 <= wire3;
            end
          else
            begin
              reg7 <= wire3[(5'h17):(3'h7)];
              reg8 <= (wire2[(1'h0):(1'h0)] ? wire3 : $unsigned((8'hbf)));
            end
          reg9 <= wire3;
        end
      if ($unsigned($unsigned(reg7)))
        begin
          reg10 = (reg7[(2'h2):(1'h1)] ?
              {$signed(($signed(reg7) * (~^(8'hbf)))),
                  (wire1 <<< reg7)} : forvar4);
          if (reg7[(4'ha):(4'h8)])
            begin
              reg11 = $unsigned(reg8);
              reg12 <= ($unsigned(wire2) ?
                  $signed($signed($unsigned({reg7}))) : (({$unsigned(reg7),
                          $signed(wire1)} ?
                      $unsigned((wire3 ?
                          reg5 : reg7)) : reg10[(5'h13):(5'h12)]) ^~ (~^(~|wire2))));
            end
          else
            begin
              reg12 <= ((-$signed($unsigned(reg10[(1'h0):(1'h0)]))) ?
                  ($unsigned({(+reg5), (reg9 << reg10)}) ?
                      (reg12 ^ (7'h43)) : ($signed(((7'h48) == reg12)) ?
                          $signed(forvar4) : $unsigned({forvar6,
                              wire0}))) : {($signed($signed(wire2)) ?
                          ((&wire2) && $signed(forvar6)) : forvar4[(1'h0):(1'h0)]),
                      $signed({$unsigned(forvar4), (forvar6 && reg7)})});
              reg13 = {$unsigned($unsigned((8'hb0))),
                  {{(forvar4 ? reg11[(4'h8):(2'h2)] : reg9)},
                      $signed($unsigned($signed(wire0)))}};
            end
          for (forvar14 = (1'h0); (forvar14 < (3'h4)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 = ($signed((reg11 ?
                      $unsigned($signed(reg5)) : $signed({reg5}))) ?
                  reg5[(3'h4):(1'h1)] : $unsigned(reg11));
              reg16 = reg12[(2'h2):(1'h0)];
              reg17 = forvar14;
              reg18 = (^~(~reg9[(3'h4):(2'h2)]));
              reg19 <= (!(($signed(reg18[(4'hd):(2'h3)]) ?
                      {reg8} : $signed(reg18[(3'h7):(2'h2)])) ?
                  {$unsigned((~^reg9))} : $unsigned((!(|reg13)))));
            end
          reg20 <= (reg10[(4'hd):(4'ha)] ^~ forvar14[(2'h3):(2'h3)]);
          reg21 <= wire3;
        end
      else
        begin
          for (forvar10 = (1'h0); (forvar10 < (3'h4)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg12 <= {wire1[(4'hd):(4'hc)]};
              reg14 <= $unsigned(({{$signed(wire3), {(7'h48)}}} ?
                  $unsigned((reg21 + $unsigned(reg20))) : $signed(($unsigned((7'h45)) ?
                      (reg20 + reg5) : reg15))));
              reg19 <= forvar6[(1'h1):(1'h1)];
              reg20 <= ($unsigned(reg8) ^ $unsigned(forvar14[(5'h12):(3'h4)]));
            end
          for (forvar21 = (1'h0); (forvar21 < (1'h0)); forvar21 = (forvar21 + (1'h1)))
            begin
              reg22 = $signed(($signed(forvar21) <= $signed(reg20)));
              reg23 = reg8[(3'h4):(1'h1)];
              reg24 <= {reg15};
            end
          reg25 <= forvar14;
          for (forvar26 = (1'h0); (forvar26 < (3'h4)); forvar26 = (forvar26 + (1'h1)))
            begin
              reg27 <= $unsigned((((reg17 ? $unsigned(wire2) : $signed(reg5)) ?
                  $signed((reg21 ?
                      reg24 : (8'hbb))) : reg7[(3'h4):(2'h2)]) >>> $signed((^(~^(8'hb1))))));
              reg28 <= reg17[(2'h2):(1'h0)];
              reg29 = $signed(($signed((reg9[(1'h1):(1'h1)] ?
                  $signed(reg9) : (8'hac))) >= reg15[(5'h13):(4'h9)]));
              reg30 <= ((((~(reg13 ? reg8 : reg8)) ?
                          ((reg8 - reg22) != reg25[(5'h11):(4'h8)]) : {$unsigned(forvar6),
                              (reg25 > reg9)}) ?
                      $unsigned(forvar14) : (($signed(reg24) & (reg11 ?
                          wire0 : reg24)) ~^ ($unsigned(reg24) - reg24[(3'h5):(3'h4)]))) ?
                  reg8 : {$unsigned(reg24[(2'h3):(1'h0)]), (^(8'h9e))});
            end
        end
      for (forvar31 = (1'h0); (forvar31 < (1'h0)); forvar31 = (forvar31 + (1'h1)))
        begin
          if (reg9[(3'h5):(1'h1)])
            begin
              reg32 <= reg15[(2'h2):(1'h1)];
              reg33 <= ({reg14[(3'h6):(1'h0)], $signed(reg20[(2'h3):(1'h0)])} ?
                  $unsigned($unsigned((reg32 ?
                      $signed(reg29) : {reg18, reg7}))) : (!reg16));
              reg34 <= wire2[(1'h1):(1'h1)];
            end
          else
            begin
              reg32 <= (reg22 ?
                  {(reg7[(4'hc):(4'hc)] ? reg13 : reg24[(3'h5):(1'h1)]),
                      forvar26[(3'h7):(3'h6)]} : (({$unsigned(forvar14),
                      $signed(reg18)} == ($signed(forvar6) ?
                      $unsigned(reg25) : (~reg8))) << forvar6[(2'h2):(1'h0)]));
            end
        end
    end
  module35 #() modinst1029 (wire1028, clk, reg14, wire0, reg28, reg30, reg5);
  assign wire1030 = $signed(reg19);
  assign wire1031 = {$signed((($unsigned(reg5) >>> (wire1030 ?
                            reg24 : reg14)) != (~&((8'hba) ? reg9 : reg7))))};
  module266 #() modinst1033 (.wire270(wire1028), .y(wire1032), .wire269(reg7), .clk(clk), .wire268(reg14), .wire267(reg9), .wire271(reg8));
  always
    @(posedge clk) begin
      reg1034 = ((reg24[(2'h2):(1'h0)] ?
          (~(~reg32)) : $unsigned($signed((reg20 || wire1031)))) + {($unsigned(wire1032) ?
              reg24 : ((reg24 ? (8'ha1) : reg28) >= wire1031[(3'h7):(3'h6)])),
          reg30});
      for (forvar1035 = (1'h0); (forvar1035 < (1'h0)); forvar1035 = (forvar1035 + (1'h1)))
        begin
          reg1036 = reg5;
          if ((7'h43))
            begin
              reg1037 <= ({{wire2[(1'h1):(1'h1)]},
                  $unsigned((^$unsigned(wire3)))} & (~&reg7[(4'hb):(3'h4)]));
            end
          else
            begin
              reg1037 <= reg8;
              reg1038 <= wire1032[(2'h2):(2'h2)];
              reg1039 = reg14;
            end
          reg1040 = $unsigned(wire1031[(1'h0):(1'h0)]);
          reg1041 = (~|(~^reg32));
        end
      reg1042 <= {($unsigned(reg1036[(4'hf):(1'h1)]) ?
              ((reg34[(4'h9):(4'h8)] != $unsigned(reg1041)) ?
                  $unsigned({wire2}) : ($signed((8'hbc)) == reg33)) : ($unsigned(reg8) ?
                  (!(7'h46)) : wire1028[(5'h11):(3'h6)]))};
      if (reg8)
        begin
          for (forvar1043 = (1'h0); (forvar1043 < (3'h4)); forvar1043 = (forvar1043 + (1'h1)))
            begin
              reg1044 = {((!reg24) ? reg1038 : $signed(wire1030)),
                  (wire1028[(5'h11):(1'h0)] ? {forvar1043} : reg7)};
            end
          for (forvar1045 = (1'h0); (forvar1045 < (2'h3)); forvar1045 = (forvar1045 + (1'h1)))
            begin
              reg1046 <= $unsigned(wire3[(5'h18):(5'h16)]);
            end
          reg1047 <= reg24;
        end
      else
        begin
          if ((reg9 >>> (~^wire3[(5'h11):(4'hb)])))
            begin
              reg1043 = $signed(($unsigned(((8'haa) ?
                      (wire1 ^ wire1030) : $signed(reg1034))) ?
                  reg1039[(4'ha):(3'h5)] : reg8[(5'h11):(5'h10)]));
              reg1045 <= $unsigned(($signed($unsigned($unsigned(wire3))) + (((wire1 ^~ reg19) * (^(8'hac))) || $unsigned($signed(wire3)))));
              reg1048 = reg30[(4'h9):(4'h9)];
            end
          else
            begin
              reg1043 = ($signed((((reg1044 ? (7'h41) : (8'ha7)) ?
                          reg9[(3'h7):(3'h4)] : wire1032[(1'h0):(1'h0)]) ?
                      reg28 : $signed(((7'h45) * (7'h4a))))) ?
                  wire0 : $unsigned($signed($signed((wire1 ? wire3 : reg28)))));
              reg1044 = reg5;
              reg1045 <= (^~$signed($unsigned($unsigned({reg1043}))));
              reg1048 = $signed(($signed($signed($unsigned(wire1))) <<< {($signed(reg1036) >>> (wire0 ?
                      reg1043 : reg21)),
                  reg14}));
              reg1049 = ((|({(reg1046 ? (8'ha0) : reg8),
                  (wire1 || reg1037)} < $unsigned(reg28[(4'hd):(4'h8)]))) ^~ forvar1035);
            end
          reg1050 <= {reg1040, reg1037};
          if ($unsigned((reg12[(2'h3):(2'h3)] ?
              reg21[(3'h6):(3'h4)] : reg32[(3'h6):(2'h2)])))
            begin
              reg1051 = (~^reg24[(2'h3):(2'h2)]);
              reg1052 = $unsigned((+($unsigned({reg1043}) <<< $unsigned(reg7))));
              reg1053 = (^reg1038);
            end
          else
            begin
              reg1054 <= (8'hbe);
              reg1055 <= ((^{{(!reg1051), $signed(wire3)},
                  (~^(+reg9))}) | reg1044);
            end
          if (wire3[(2'h3):(2'h2)])
            begin
              reg1056 = $unsigned((((!reg8) ?
                      $signed((^~reg7)) : $unsigned(wire3)) ?
                  (~^((~^(7'h46)) ?
                      forvar1045[(4'hd):(1'h0)] : (^reg25))) : ({reg1041} ?
                      $signed($signed(wire3)) : $signed(wire1028))));
            end
          else
            begin
              reg1056 = $signed($unsigned(reg30[(4'hc):(2'h2)]));
              reg1057 <= reg1034;
              reg1058 = ($signed($signed(wire0)) ? reg1046 : reg1036);
              reg1059 <= reg9;
              reg1060 <= reg30;
            end
        end
      if (($unsigned($unsigned((((8'hb7) ? reg1039 : reg1045) ^~ (reg1057 ?
          wire1031 : (8'hba))))) <= (~|((!(reg1055 <<< wire0)) * reg21))))
        begin
          reg1061 <= ((~|((~^(~|(8'ha2))) ?
                  {(reg28 ? reg1051 : reg1037)} : {(~&reg5)})) ?
              $unsigned($signed(((reg21 * forvar1035) ?
                  (|(8'haa)) : $signed(forvar1043)))) : $unsigned($signed($signed($signed(reg1058)))));
        end
      else
        begin
          reg1061 <= ($signed((!$signed((wire3 ^ reg1044)))) ?
              reg32 : $unsigned(reg1048));
          reg1062 = (^~reg1061[(4'he):(1'h0)]);
        end
    end
  assign wire1063 = reg1042;
  assign wire1064 = (~^(&reg1060[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      if ($unsigned((!{{(reg24 + reg1045), reg1042}})))
        begin
          if ((~&($unsigned($signed((-reg34))) ^ ({(wire1 ?
                  (8'hb1) : reg27)} + (reg8[(4'hd):(4'ha)] ?
              (reg1061 ^~ reg21) : (+reg1061))))))
            begin
              reg1065 = ((-reg1046[(2'h2):(1'h1)]) ^~ $signed($unsigned((reg5[(2'h2):(1'h1)] ?
                  reg1060[(3'h4):(2'h3)] : $signed(wire1063)))));
              reg1066 <= (|reg24);
              reg1067 <= ((^~{(|reg1037[(5'h11):(4'ha)])}) ~^ $unsigned((+(-reg19))));
            end
          else
            begin
              reg1065 = wire3;
              reg1068 = {{($unsigned({wire1032}) ?
                          ($unsigned(reg1066) ?
                              $unsigned(wire1030) : ((8'haa) ?
                                  reg25 : reg1045)) : reg1047[(3'h7):(3'h4)]),
                      $signed($signed(reg21))},
                  {$unsigned(($signed(wire0) >= (~|reg1061)))}};
              reg1069 <= {(^~(^(reg1045 ~^ {wire1, (8'hb2)})))};
              reg1070 <= ((~^((~|$signed(reg1065)) ?
                      ($signed(reg1066) ?
                          (reg1066 ~^ reg12) : (wire1064 >>> reg5)) : $signed(reg33))) ?
                  $signed($signed((reg20[(4'hb):(4'h8)] ?
                      reg32[(1'h1):(1'h0)] : reg28))) : reg32[(3'h7):(2'h2)]);
            end
          if (reg1068)
            begin
              reg1071 <= (8'had);
              reg1072 <= wire1028[(5'h13):(4'hf)];
            end
          else
            begin
              reg1073 = reg19;
              reg1074 = ($unsigned($signed(({reg20, reg24} >> (reg1047 ?
                  reg21 : reg5)))) > wire1031);
              reg1075 = (($signed(($signed(reg1073) <<< (~^(8'hb6)))) ?
                      reg1038 : $signed(reg28[(2'h3):(2'h2)])) ?
                  reg1068 : ((((reg1069 << reg1042) | {reg7,
                          wire1031}) && (~(reg1061 ^~ reg24))) ?
                      ((8'ha7) ? reg1047 : (~(reg27 << (8'h9e)))) : (((wire2 ?
                                  reg1072 : reg14) ?
                              reg1071[(4'h8):(3'h5)] : (^reg32)) ?
                          (((8'hb4) ^ reg1069) & {wire3}) : ({wire1064} ?
                              $unsigned((8'h9e)) : (reg7 <= reg24)))));
              reg1076 <= $signed((({reg9[(1'h1):(1'h1)]} >= (8'hbf)) ?
                  wire1 : (^(~^$unsigned(reg25)))));
            end
          reg1077 = $unsigned({reg34});
          reg1078 = ($unsigned((|(+(-reg28)))) ?
              (~|$unsigned(reg1068)) : reg1068);
          for (forvar1079 = (1'h0); (forvar1079 < (1'h1)); forvar1079 = (forvar1079 + (1'h1)))
            begin
              reg1080 <= (^~(((8'haa) < $signed(((8'h9f) ?
                  reg1078 : (8'hb8)))) << (reg1068[(2'h3):(2'h2)] >= ($signed(wire1) != (reg1060 ?
                  reg24 : (8'hbf))))));
              reg1081 <= reg1071[(3'h5):(1'h1)];
              reg1082 <= ((|((reg1081[(1'h0):(1'h0)] ~^ $unsigned((8'hb0))) ?
                      ($unsigned((8'hb9)) ?
                          reg19[(3'h4):(3'h4)] : $unsigned(reg28)) : (~^(7'h4a)))) ?
                  $unsigned(reg1070) : $unsigned({{(^(8'hbc)), wire1064}}));
              reg1083 <= reg14;
            end
        end
      else
        begin
          reg1065 = reg1073;
          reg1066 <= ((^~$signed(reg1076[(4'hf):(1'h1)])) ? (8'hb1) : (+reg14));
          reg1067 <= $signed(reg1080);
        end
    end
  always
    @(posedge clk) begin
      reg1084 = $signed((~$signed((^~(wire1064 & reg1038)))));
    end
  always
    @(posedge clk) begin
      reg1085 <= (reg1061[(4'he):(3'h5)] ?
          $signed(reg1054[(3'h5):(1'h0)]) : (!$signed(($signed((8'haa)) ?
              (reg33 ? reg1080 : wire1063) : (^reg9)))));
      reg1086 <= $unsigned(reg8[(4'hb):(4'ha)]);
      reg1087 = (({wire1030,
              {(reg24 ? (8'hb4) : (8'ha0))}} >> (~(~|$signed((8'ha4))))) ?
          wire1 : reg1057[(2'h2):(2'h2)]);
    end
  assign wire1088 = ((!$signed((~^(!reg27)))) <<< $unsigned($signed((^$unsigned(reg1083)))));
  assign wire1089 = ($unsigned({(&$signed(reg1072))}) | $unsigned(reg24[(3'h4):(1'h0)]));
  assign wire1090 = ($unsigned(reg1045) ?
                        (reg1054[(1'h0):(1'h0)] >> $unsigned((8'ha7))) : reg1045[(3'h5):(2'h2)]);
  always
    @(posedge clk) begin
      reg1091 <= reg1070;
    end
  assign wire1092 = (~^$signed($signed($unsigned(((8'hb1) ?
                        reg1076 : reg1083)))));
  always
    @(posedge clk) begin
      reg1093 = ($signed($signed((!(reg25 ?
          reg1061 : reg1055)))) <= reg1067[(1'h0):(1'h0)]);
      for (forvar1094 = (1'h0); (forvar1094 < (2'h2)); forvar1094 = (forvar1094 + (1'h1)))
        begin
          reg1095 <= (8'hbd);
        end
    end
  always
    @(posedge clk) begin
      if ($signed({$signed($unsigned({reg1070, (8'hbe)}))}))
        begin
          if ($signed(((~$unsigned((^reg28))) != wire2[(2'h2):(1'h1)])))
            begin
              reg1096 <= ((~$unsigned(reg30[(1'h1):(1'h1)])) ?
                  (reg9[(4'h9):(3'h5)] ?
                      $signed($unsigned($signed((8'h9c)))) : $signed($signed($signed(reg1071)))) : (reg34[(3'h6):(2'h3)] >>> reg1076));
              reg1097 <= $signed(reg1083);
            end
          else
            begin
              reg1096 <= reg1091;
              reg1098 = (&reg1066);
            end
          reg1099 <= (!((&reg1050) ?
              {((reg1083 <<< (8'ha9)) || reg1060[(4'hc):(4'ha)]),
                  reg1067} : reg1072[(3'h5):(1'h1)]));
          reg1100 <= reg1038;
          if (wire1088[(4'hd):(4'hc)])
            begin
              reg1101 = $unsigned(reg24[(2'h2):(2'h2)]);
            end
          else
            begin
              reg1102 <= ($unsigned(reg1061) <<< ({(8'haa),
                  ($unsigned((8'h9f)) | reg1055)} || (wire1064[(4'he):(4'he)] - {(8'ha5)})));
              reg1103 <= {$unsigned(((~(wire1031 != (8'hb1))) ?
                      $signed({(8'hbb), reg24}) : (reg27 ?
                          reg1098[(3'h5):(2'h3)] : (-wire1088))))};
              reg1104 = ({{(reg1067 >= $unsigned(reg33))}} & reg21[(1'h0):(1'h0)]);
              reg1105 = (reg28[(5'h13):(3'h7)] ^ $signed((({(8'hbf),
                      reg1104} + $unsigned(reg1097)) ?
                  $unsigned($signed(reg7)) : $unsigned((|reg1070)))));
            end
        end
      else
        begin
          reg1096 <= (reg32[(1'h1):(1'h0)] ?
              $unsigned((&{{reg1096},
                  (^reg1054)})) : $unsigned({$signed({reg12}),
                  $signed(((8'hab) >> reg1037))}));
        end
      if (((-(-reg1038[(5'h13):(5'h10)])) ?
          reg1055[(2'h3):(2'h3)] : ($signed(reg1102[(4'h8):(3'h6)]) ?
              $unsigned(reg14) : (8'hb6))))
        begin
          reg1106 <= $unsigned($unsigned($signed((-$unsigned(reg1101)))));
          reg1107 <= (|$unsigned(((~$signed(reg1076)) ?
              ((~&reg1106) != ((8'hbf) ?
                  reg1083 : wire1031)) : (reg1085[(2'h2):(1'h1)] * (8'ha8)))));
        end
      else
        begin
          reg1106 <= reg25[(4'hb):(1'h1)];
        end
      reg1108 = (~wire0[(4'hb):(3'h5)]);
      reg1109 <= $signed($unsigned(((reg1050 - {(8'hba), reg1061}) ?
          ((8'h9c) & reg1060[(1'h0):(1'h0)]) : ((^~reg1097) <<< $signed(reg1098)))));
    end
  always
    @(posedge clk) begin
      reg1110 = reg1057;
      for (forvar1111 = (1'h0); (forvar1111 < (3'h4)); forvar1111 = (forvar1111 + (1'h1)))
        begin
          reg1112 <= (+reg19);
          reg1113 = reg1067;
          reg1114 = (+((^~((reg8 ? wire1 : reg1038) ?
              reg1085 : (reg1106 ? (8'hba) : reg28))) * {$unsigned({(8'ha2),
                  wire1089}),
              (8'hac)}));
          reg1115 = (reg1082[(3'h6):(3'h6)] ?
              (reg1071[(4'hb):(4'ha)] ?
                  reg1046[(3'h5):(2'h3)] : reg1095) : reg1080);
          reg1116 = ((~|(+$signed(reg1114))) >> ((reg1061[(1'h0):(1'h0)] ?
              reg1066[(4'ha):(1'h0)] : reg21) ^~ wire3[(5'h16):(3'h4)]));
        end
      if (reg9[(4'h9):(3'h4)])
        begin
          for (forvar1117 = (1'h0); (forvar1117 < (1'h1)); forvar1117 = (forvar1117 + (1'h1)))
            begin
              reg1118 <= (($unsigned((!$unsigned(reg14))) + {$signed(reg1055)}) < forvar1117);
              reg1119 = $signed({reg1115});
              reg1120 <= ($signed(reg21) || wire3);
            end
          reg1121 <= ($signed(((~reg1120) + (reg1038 >>> (~|reg1099)))) ?
              {wire1[(1'h1):(1'h1)]} : ((8'hab) * wire1092));
          if ($unsigned(((+(reg1055 + (^~reg1046))) >> reg1114[(2'h3):(1'h0)])))
            begin
              reg1122 <= $signed((reg1061[(4'hf):(1'h0)] + ({reg1045,
                  reg1109} << $signed((reg1086 ? reg1076 : wire1088)))));
              reg1123 <= reg7;
              reg1124 = $signed(((~^((~|reg1123) ?
                      $unsigned(wire3) : (~|reg1086))) ?
                  (~&$unsigned(((8'hbe) ?
                      reg1114 : reg1085))) : $signed((^~(reg1085 ?
                      reg1070 : reg33)))));
              reg1125 = reg33[(4'h8):(3'h4)];
            end
          else
            begin
              reg1122 <= (wire2 ?
                  $signed(reg1124[(3'h6):(3'h4)]) : ((|wire3) && {$signed((!reg1085)),
                      {reg1046}}));
            end
          reg1126 = $unsigned(($signed({reg1118, (8'hb9)}) << wire1031));
          for (forvar1127 = (1'h0); (forvar1127 < (2'h2)); forvar1127 = (forvar1127 + (1'h1)))
            begin
              reg1128 <= (^(&($signed($signed(wire1064)) ?
                  (reg27 <= $unsigned(reg1095)) : $signed($unsigned(reg1070)))));
              reg1129 <= ((~^{(~^(8'ha3))}) ?
                  $signed((-reg1042)) : (reg1109 ?
                      (reg1060[(3'h6):(1'h0)] ?
                          (!reg1091) : reg30[(3'h6):(3'h6)]) : $unsigned((~^reg1114))));
            end
        end
      else
        begin
          if ($unsigned($unsigned((({wire1090, reg20} ~^ (reg1109 ?
              (8'hb6) : reg14)) & (~reg19[(4'h9):(3'h7)])))))
            begin
              reg1117 = reg1102;
              reg1119 = ((reg1123[(4'ha):(1'h0)] ?
                  $signed({(reg1096 ~^ (8'hbd))}) : wire1088) >= ((reg1055 ?
                  {reg9} : $signed(reg1102)) ~^ ((reg1103 ~^ reg1110[(2'h3):(1'h1)]) ?
                  $signed((reg1070 || reg9)) : (reg1045[(1'h1):(1'h1)] ?
                      (!reg32) : {wire2}))));
              reg1120 <= reg1066[(4'hb):(1'h1)];
              reg1124 = $signed(($signed(reg30[(3'h6):(1'h1)]) <= (reg1106 ?
                  ({(8'hb4)} ? $signed(reg1042) : {reg1122}) : (((7'h46) ?
                          reg1057 : reg1038) ?
                      (reg1045 <= wire1032) : (-reg1085)))));
              reg1127 <= reg21;
            end
          else
            begin
              reg1117 = (((+reg1124[(3'h6):(3'h4)]) | reg28[(4'hb):(3'h6)]) ?
                  wire1089 : $signed(reg1114));
              reg1118 <= forvar1127[(4'h9):(4'h9)];
              reg1120 <= reg1042;
              reg1124 = {((~((~^(8'ha8)) < (+(8'ha4)))) ?
                      (&reg1110[(2'h2):(1'h1)]) : {($unsigned(reg5) >= $unsigned(reg1072))})};
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1130 = (1'h0); (forvar1130 < (1'h1)); forvar1130 = (forvar1130 + (1'h1)))
        begin
          reg1131 = ($unsigned({(reg1047 & (|(7'h49)))}) ?
              (reg1091 & wire3[(5'h16):(5'h15)]) : (($unsigned((^~(8'hab))) <= reg14) <= reg1100[(2'h3):(2'h2)]));
          for (forvar1132 = (1'h0); (forvar1132 < (3'h4)); forvar1132 = (forvar1132 + (1'h1)))
            begin
              reg1133 = ($signed(reg34[(4'hc):(3'h6)]) ?
                  wire1028[(1'h1):(1'h0)] : ((($unsigned(reg34) ?
                              (reg1046 ? (8'ha5) : wire1031) : $signed(reg25)) ?
                          reg1055[(2'h3):(2'h2)] : ($signed(reg1057) ?
                              (8'hb4) : (reg1121 >>> reg1057))) ?
                      (8'hac) : ($signed({reg1071, reg1076}) ?
                          reg1085 : ({reg1099,
                              reg25} ~^ (reg1118 ^ wire1088)))));
            end
          for (forvar1134 = (1'h0); (forvar1134 < (2'h2)); forvar1134 = (forvar1134 + (1'h1)))
            begin
              reg1135 <= (((~&reg1037) ?
                  (~(~&reg1076)) : ((^~$unsigned(reg14)) ~^ ($unsigned(reg1120) * $signed(reg25)))) + $signed(reg1082));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module35
#(parameter param1026 = ((((&((8'hae) ? (8'h9f) : (7'h49))) > {{(8'hb4), (8'h9d)}}) < (7'h42)) == (|({((8'h9d) ? (8'hb0) : (8'hba))} + (|((8'ha8) ^ (8'ha0)))))), 
parameter param1027 = {({(&(^~param1026))} ? {(+(param1026 > param1026))} : (8'haf))})
(y, clk, wire40, wire39, wire38, wire37, wire36);
  output wire [(32'hdf2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire40;
  input wire [(3'h6):(1'h0)] wire39;
  input wire signed [(5'h18):(1'h0)] wire38;
  input wire [(4'h9):(1'h0)] wire37;
  input wire signed [(4'hc):(1'h0)] wire36;
  wire signed [(4'he):(1'h0)] wire1025;
  wire [(5'h13):(1'h0)] wire854;
  wire signed [(5'h17):(1'h0)] wire853;
  wire signed [(5'h14):(1'h0)] wire834;
  wire signed [(2'h2):(1'h0)] wire819;
  wire [(5'h12):(1'h0)] wire86;
  wire signed [(4'h8):(1'h0)] wire53;
  wire signed [(2'h3):(1'h0)] wire41;
  reg signed [(4'h8):(1'h0)] reg1023 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1019 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1018 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1008 = (1'h0);
  reg [(5'h14):(1'h0)] reg1006 = (1'h0);
  reg [(5'h15):(1'h0)] reg1003 = (1'h0);
  reg [(5'h12):(1'h0)] reg1002 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1001 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1000 = (1'h0);
  reg [(5'h12):(1'h0)] reg999 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg995 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg993 = (1'h0);
  reg [(2'h3):(1'h0)] reg988 = (1'h0);
  reg [(5'h16):(1'h0)] reg985 = (1'h0);
  reg [(5'h10):(1'h0)] reg984 = (1'h0);
  reg [(4'hf):(1'h0)] reg983 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg980 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg979 = (1'h0);
  reg [(4'hf):(1'h0)] reg977 = (1'h0);
  reg [(5'h17):(1'h0)] reg975 = (1'h0);
  reg signed [(4'he):(1'h0)] reg973 = (1'h0);
  reg [(5'h12):(1'h0)] reg971 = (1'h0);
  reg [(3'h7):(1'h0)] reg970 = (1'h0);
  reg signed [(4'he):(1'h0)] reg969 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg968 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg962 = (1'h0);
  reg [(2'h2):(1'h0)] reg960 = (1'h0);
  reg [(4'he):(1'h0)] reg958 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg957 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg956 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg952 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg946 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg945 = (1'h0);
  reg signed [(4'he):(1'h0)] reg943 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg938 = (1'h0);
  reg [(5'h16):(1'h0)] reg935 = (1'h0);
  reg [(4'hd):(1'h0)] reg933 = (1'h0);
  reg [(4'hf):(1'h0)] reg929 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg924 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg921 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg920 = (1'h0);
  reg [(5'h12):(1'h0)] reg917 = (1'h0);
  reg [(5'h17):(1'h0)] reg916 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg914 = (1'h0);
  reg [(4'he):(1'h0)] reg913 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg912 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg909 = (1'h0);
  reg [(5'h17):(1'h0)] reg908 = (1'h0);
  reg [(5'h15):(1'h0)] reg905 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg904 = (1'h0);
  reg [(5'h12):(1'h0)] reg901 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg897 = (1'h0);
  reg signed [(4'he):(1'h0)] reg896 = (1'h0);
  reg [(3'h6):(1'h0)] reg895 = (1'h0);
  reg [(5'h15):(1'h0)] reg892 = (1'h0);
  reg signed [(4'he):(1'h0)] reg890 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg887 = (1'h0);
  reg [(4'ha):(1'h0)] reg886 = (1'h0);
  reg [(5'h11):(1'h0)] reg885 = (1'h0);
  reg [(5'h18):(1'h0)] reg883 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg877 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg875 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg873 = (1'h0);
  reg [(4'he):(1'h0)] reg872 = (1'h0);
  reg [(4'h8):(1'h0)] reg871 = (1'h0);
  reg [(2'h2):(1'h0)] reg870 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg867 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg862 = (1'h0);
  reg [(3'h6):(1'h0)] reg858 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg857 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg856 = (1'h0);
  reg [(4'h8):(1'h0)] reg855 = (1'h0);
  reg signed [(4'he):(1'h0)] reg851 = (1'h0);
  reg [(4'h9):(1'h0)] reg850 = (1'h0);
  reg [(4'h9):(1'h0)] reg847 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg846 = (1'h0);
  reg [(4'ha):(1'h0)] reg841 = (1'h0);
  reg [(4'ha):(1'h0)] reg837 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg835 = (1'h0);
  reg [(4'hc):(1'h0)] reg833 = (1'h0);
  reg [(5'h11):(1'h0)] reg827 = (1'h0);
  reg [(4'hd):(1'h0)] reg823 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg830 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg828 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg824 = (1'h0);
  reg [(5'h16):(1'h0)] reg72 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg80 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg79 = (1'h0);
  reg [(5'h11):(1'h0)] reg77 = (1'h0);
  reg [(5'h15):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg70 = (1'h0);
  reg [(5'h10):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg63 = (1'h0);
  reg [(3'h5):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg60 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg [(5'h14):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg55 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg52 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg50 = (1'h0);
  reg [(4'hb):(1'h0)] reg45 = (1'h0);
  reg [(5'h17):(1'h0)] reg43 = (1'h0);
  reg [(4'hf):(1'h0)] reg1024 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1022 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1021 = (1'h0);
  reg [(3'h7):(1'h0)] reg1020 = (1'h0);
  reg [(5'h16):(1'h0)] reg1017 = (1'h0);
  reg [(4'hc):(1'h0)] reg1016 = (1'h0);
  reg [(3'h4):(1'h0)] reg1015 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1014 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1013 = (1'h0);
  reg [(4'he):(1'h0)] forvar1012 = (1'h0);
  reg [(5'h12):(1'h0)] reg1011 = (1'h0);
  reg [(5'h15):(1'h0)] reg1010 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1009 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1007 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1001 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1005 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1004 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg998 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg997 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg996 = (1'h0);
  reg [(5'h16):(1'h0)] reg994 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg992 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg991 = (1'h0);
  reg [(4'hd):(1'h0)] reg990 = (1'h0);
  reg [(5'h16):(1'h0)] reg989 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg987 = (1'h0);
  reg [(5'h18):(1'h0)] reg986 = (1'h0);
  reg [(5'h16):(1'h0)] reg982 = (1'h0);
  reg [(4'h8):(1'h0)] reg981 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar978 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg976 = (1'h0);
  reg signed [(4'he):(1'h0)] reg974 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar973 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg972 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg967 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg966 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg965 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar964 = (1'h0);
  reg [(2'h2):(1'h0)] reg963 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg961 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg959 = (1'h0);
  reg [(2'h3):(1'h0)] forvar955 = (1'h0);
  reg [(5'h17):(1'h0)] reg954 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg955 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar954 = (1'h0);
  reg [(3'h7):(1'h0)] reg953 = (1'h0);
  reg [(5'h16):(1'h0)] reg951 = (1'h0);
  reg [(4'hc):(1'h0)] reg950 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg949 = (1'h0);
  reg [(5'h12):(1'h0)] reg948 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar947 = (1'h0);
  reg [(3'h5):(1'h0)] reg944 = (1'h0);
  reg [(3'h4):(1'h0)] reg942 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg941 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg940 = (1'h0);
  reg [(5'h12):(1'h0)] forvar939 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar937 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar936 = (1'h0);
  reg [(4'hc):(1'h0)] reg934 = (1'h0);
  reg [(4'hf):(1'h0)] reg932 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar931 = (1'h0);
  reg [(2'h3):(1'h0)] reg930 = (1'h0);
  reg [(3'h4):(1'h0)] reg928 = (1'h0);
  reg [(5'h11):(1'h0)] reg927 = (1'h0);
  reg [(5'h10):(1'h0)] reg926 = (1'h0);
  reg [(5'h14):(1'h0)] reg925 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar923 = (1'h0);
  reg [(3'h4):(1'h0)] reg922 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg919 = (1'h0);
  reg [(5'h16):(1'h0)] forvar918 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar915 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg911 = (1'h0);
  reg [(4'hd):(1'h0)] reg910 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar907 = (1'h0);
  reg [(4'hd):(1'h0)] reg906 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg907 = (1'h0);
  reg [(5'h16):(1'h0)] forvar906 = (1'h0);
  reg [(3'h4):(1'h0)] reg903 = (1'h0);
  reg [(4'h9):(1'h0)] reg902 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar900 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg899 = (1'h0);
  reg [(5'h16):(1'h0)] reg898 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg894 = (1'h0);
  reg [(2'h3):(1'h0)] reg893 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg891 = (1'h0);
  reg [(5'h11):(1'h0)] reg889 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg888 = (1'h0);
  reg [(4'hb):(1'h0)] reg884 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg882 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg881 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar880 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg879 = (1'h0);
  reg [(5'h14):(1'h0)] forvar878 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar876 = (1'h0);
  reg [(4'hb):(1'h0)] forvar874 = (1'h0);
  reg [(2'h2):(1'h0)] reg869 = (1'h0);
  reg [(3'h7):(1'h0)] reg866 = (1'h0);
  reg [(4'h8):(1'h0)] reg865 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg863 = (1'h0);
  reg [(5'h13):(1'h0)] reg861 = (1'h0);
  reg signed [(4'he):(1'h0)] reg860 = (1'h0);
  reg [(4'h9):(1'h0)] reg859 = (1'h0);
  reg [(4'h9):(1'h0)] reg852 = (1'h0);
  reg [(4'hd):(1'h0)] reg849 = (1'h0);
  reg [(4'he):(1'h0)] reg848 = (1'h0);
  reg [(4'ha):(1'h0)] forvar845 = (1'h0);
  reg [(5'h14):(1'h0)] reg844 = (1'h0);
  reg [(3'h6):(1'h0)] reg843 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg842 = (1'h0);
  reg [(5'h17):(1'h0)] forvar837 = (1'h0);
  reg signed [(4'he):(1'h0)] reg836 = (1'h0);
  reg [(5'h10):(1'h0)] reg840 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg839 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg838 = (1'h0);
  reg [(4'h8):(1'h0)] forvar836 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg832 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg831 = (1'h0);
  reg [(4'h9):(1'h0)] reg829 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar827 = (1'h0);
  reg [(4'hf):(1'h0)] reg826 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg825 = (1'h0);
  reg [(5'h13):(1'h0)] forvar823 = (1'h0);
  reg [(5'h11):(1'h0)] reg822 = (1'h0);
  reg signed [(4'he):(1'h0)] reg821 = (1'h0);
  reg [(4'hd):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar83 = (1'h0);
  reg [(5'h12):(1'h0)] forvar71 = (1'h0);
  reg [(4'ha):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg82 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg81 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg78 = (1'h0);
  reg [(4'ha):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg75 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg73 = (1'h0);
  reg [(5'h13):(1'h0)] forvar72 = (1'h0);
  reg [(4'hf):(1'h0)] reg71 = (1'h0);
  reg [(5'h16):(1'h0)] reg69 = (1'h0);
  reg [(5'h17):(1'h0)] reg67 = (1'h0);
  reg [(5'h11):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg62 = (1'h0);
  reg [(4'hf):(1'h0)] forvar57 = (1'h0);
  reg [(4'h9):(1'h0)] forvar56 = (1'h0);
  reg [(5'h14):(1'h0)] reg54 = (1'h0);
  reg [(3'h4):(1'h0)] reg51 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg48 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg46 = (1'h0);
  reg [(4'ha):(1'h0)] forvar44 = (1'h0);
  reg [(5'h17):(1'h0)] reg42 = (1'h0);
  assign y = {wire1025,
                 wire854,
                 wire853,
                 wire834,
                 wire819,
                 wire86,
                 wire53,
                 wire41,
                 reg1023,
                 reg1019,
                 reg1018,
                 reg1012,
                 reg1008,
                 reg1006,
                 reg1003,
                 reg1002,
                 reg1001,
                 reg1000,
                 reg999,
                 reg995,
                 reg993,
                 reg988,
                 reg985,
                 reg984,
                 reg983,
                 reg980,
                 reg979,
                 reg977,
                 reg975,
                 reg973,
                 reg971,
                 reg970,
                 reg969,
                 reg968,
                 reg962,
                 reg960,
                 reg958,
                 reg957,
                 reg956,
                 reg952,
                 reg946,
                 reg945,
                 reg943,
                 reg938,
                 reg935,
                 reg933,
                 reg929,
                 reg924,
                 reg921,
                 reg920,
                 reg917,
                 reg916,
                 reg914,
                 reg913,
                 reg912,
                 reg900,
                 reg909,
                 reg908,
                 reg905,
                 reg904,
                 reg901,
                 reg897,
                 reg896,
                 reg895,
                 reg892,
                 reg890,
                 reg887,
                 reg886,
                 reg885,
                 reg883,
                 reg877,
                 reg875,
                 reg873,
                 reg872,
                 reg871,
                 reg870,
                 reg868,
                 reg867,
                 reg864,
                 reg862,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg851,
                 reg850,
                 reg847,
                 reg846,
                 reg841,
                 reg837,
                 reg835,
                 reg833,
                 reg827,
                 reg823,
                 reg830,
                 reg828,
                 reg824,
                 reg72,
                 reg80,
                 reg79,
                 reg77,
                 reg74,
                 reg70,
                 reg68,
                 reg65,
                 reg64,
                 reg63,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg55,
                 reg52,
                 reg50,
                 reg45,
                 reg43,
                 reg1024,
                 reg1022,
                 reg1021,
                 reg1020,
                 reg1017,
                 reg1016,
                 reg1015,
                 reg1014,
                 reg1013,
                 forvar1012,
                 reg1011,
                 reg1010,
                 reg1009,
                 reg1007,
                 forvar1001,
                 reg1005,
                 reg1004,
                 reg998,
                 reg997,
                 reg996,
                 reg994,
                 reg992,
                 reg991,
                 reg990,
                 reg989,
                 reg987,
                 reg986,
                 reg982,
                 reg981,
                 forvar978,
                 reg976,
                 reg974,
                 forvar973,
                 reg972,
                 reg967,
                 reg966,
                 reg965,
                 forvar964,
                 reg963,
                 reg961,
                 reg959,
                 forvar955,
                 reg954,
                 reg955,
                 forvar954,
                 reg953,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 forvar947,
                 reg944,
                 reg942,
                 reg941,
                 reg940,
                 forvar939,
                 forvar937,
                 forvar936,
                 reg934,
                 reg932,
                 forvar931,
                 reg930,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 forvar923,
                 reg922,
                 reg919,
                 forvar918,
                 forvar915,
                 reg911,
                 reg910,
                 forvar907,
                 reg906,
                 reg907,
                 forvar906,
                 reg903,
                 reg902,
                 forvar900,
                 reg899,
                 reg898,
                 reg894,
                 reg893,
                 reg891,
                 reg889,
                 reg888,
                 reg884,
                 reg882,
                 reg881,
                 forvar880,
                 reg879,
                 forvar878,
                 forvar876,
                 forvar874,
                 reg869,
                 reg866,
                 reg865,
                 reg863,
                 reg861,
                 reg860,
                 reg859,
                 reg852,
                 reg849,
                 reg848,
                 forvar845,
                 reg844,
                 reg843,
                 reg842,
                 forvar837,
                 reg836,
                 reg840,
                 reg839,
                 reg838,
                 forvar836,
                 reg832,
                 reg831,
                 reg829,
                 forvar827,
                 reg826,
                 reg825,
                 forvar823,
                 reg822,
                 reg821,
                 reg85,
                 reg84,
                 forvar83,
                 forvar71,
                 reg83,
                 reg82,
                 reg81,
                 reg78,
                 reg76,
                 reg75,
                 reg73,
                 forvar72,
                 reg71,
                 reg69,
                 reg67,
                 reg66,
                 reg62,
                 forvar57,
                 forvar56,
                 reg54,
                 reg51,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 forvar44,
                 reg42,
                 (1'h0)};
  assign wire41 = ($signed($unsigned($unsigned((wire36 ?
                      wire40 : wire40)))) - $unsigned((($signed(wire37) <<< $signed(wire37)) ?
                      (-wire37[(1'h1):(1'h0)]) : (~^$unsigned(wire36)))));
  always
    @(posedge clk) begin
      reg42 = $signed($signed((wire36 >> wire37[(1'h0):(1'h0)])));
      reg43 <= ($signed((^wire37[(3'h7):(1'h0)])) ?
          $unsigned($signed(wire38[(5'h12):(3'h5)])) : (wire40 <<< (+$signed($signed((8'hbb))))));
      for (forvar44 = (1'h0); (forvar44 < (2'h3)); forvar44 = (forvar44 + (1'h1)))
        begin
          reg45 <= $signed(wire37);
          if (((!$signed((~^(wire37 * reg45)))) >> wire37))
            begin
              reg46 = $signed(($signed({$unsigned((8'hb2))}) ?
                  $unsigned(({wire41} ?
                      ((8'hbb) < reg45) : $unsigned(reg43))) : {((forvar44 ?
                          reg43 : (8'hac)) >> {wire39})}));
            end
          else
            begin
              reg46 = reg45;
              reg47 = reg42[(5'h10):(4'hd)];
              reg48 = {wire38[(3'h6):(3'h4)], reg43};
              reg49 = $signed($unsigned((&(^~wire37[(3'h7):(3'h6)]))));
            end
          reg50 <= ((~wire40) ?
              reg45 : (|(&((reg43 >= reg43) - (wire40 ? wire38 : wire38)))));
          reg51 = reg49;
          reg52 <= reg42[(4'hf):(2'h2)];
        end
    end
  assign wire53 = (~($unsigned(wire41[(2'h2):(2'h2)]) ?
                      (((~^wire36) ~^ wire37) ?
                          $unsigned({wire39}) : (reg43[(2'h2):(1'h1)] ?
                              $unsigned(wire39) : reg50[(2'h2):(1'h1)])) : wire37));
  always
    @(posedge clk) begin
      reg54 = (~|($signed(wire41) ?
          (reg50[(3'h5):(3'h4)] ^~ $unsigned({(8'h9c)})) : (8'h9c)));
      reg55 <= ($signed(reg45[(4'hb):(2'h2)]) || (~|$unsigned(reg52[(1'h1):(1'h0)])));
      for (forvar56 = (1'h0); (forvar56 < (2'h3)); forvar56 = (forvar56 + (1'h1)))
        begin
          for (forvar57 = (1'h0); (forvar57 < (2'h3)); forvar57 = (forvar57 + (1'h1)))
            begin
              reg58 <= reg52;
              reg59 <= $signed($signed($signed($signed($unsigned(forvar56)))));
              reg60 <= $signed(wire40);
              reg61 <= reg45[(1'h1):(1'h1)];
              reg62 = (|reg61);
            end
          if (({reg61[(1'h1):(1'h1)]} != ($unsigned($signed(reg60)) <<< wire39[(3'h4):(1'h0)])))
            begin
              reg63 <= (~^(wire53 + $signed(wire39)));
              reg64 <= ($signed($signed((~|(reg50 <<< (8'hbf))))) ^ ($unsigned({$unsigned(wire37)}) ?
                  reg43 : reg61[(1'h1):(1'h1)]));
              reg65 <= ($unsigned($signed($unsigned(((7'h47) ?
                  wire36 : reg58)))) ~^ forvar56[(4'h8):(1'h1)]);
              reg66 = reg43[(4'hc):(1'h1)];
            end
          else
            begin
              reg63 <= reg58;
            end
          reg67 = (^~((((-wire40) ? $unsigned(wire39) : {forvar56, (7'h45)}) ?
                  forvar57 : reg52[(2'h3):(2'h2)]) ?
              wire38 : ((+(reg58 & reg65)) ?
                  $unsigned({wire41}) : $unsigned(reg65[(1'h0):(1'h0)]))));
          if ((~&reg55))
            begin
              reg68 <= wire37[(2'h2):(1'h1)];
              reg69 = wire38;
            end
          else
            begin
              reg68 <= $unsigned(forvar56);
              reg70 <= ({$signed(($unsigned(reg50) ?
                          wire38[(4'he):(4'he)] : (wire38 ? reg54 : reg45))),
                      (($signed(reg66) ?
                          ((8'hbc) | reg52) : (wire36 ?
                              reg60 : (7'h47))) >= (+$signed(forvar56)))} ?
                  $signed($signed(reg55)) : ((~^wire36[(1'h0):(1'h0)]) >= $unsigned(wire37)));
            end
        end
      if (({($unsigned(reg52[(3'h5):(1'h1)]) | ($unsigned((7'h43)) != reg52)),
              (reg67[(1'h1):(1'h0)] ? (7'h47) : reg45[(2'h2):(2'h2)])} ?
          ((~&$unsigned((^~reg63))) >= ((((8'hbf) ^~ reg59) ?
                  $unsigned((8'h9f)) : $unsigned(wire53)) ?
              (((8'hbd) ^ (8'hb6)) <<< (&(7'h45))) : $unsigned((reg61 ?
                  reg52 : reg68)))) : ($signed($signed(reg61)) == {$unsigned((forvar56 ?
                  reg70 : reg66))})))
        begin
          reg71 = (~reg70);
          for (forvar72 = (1'h0); (forvar72 < (1'h1)); forvar72 = (forvar72 + (1'h1)))
            begin
              reg73 = $unsigned((+$signed((-(^reg70)))));
              reg74 <= reg59;
              reg75 = (+reg70[(4'ha):(3'h7)]);
              reg76 = {$signed((reg71 * ({reg67} ~^ reg55[(3'h4):(1'h1)])))};
            end
          if ($signed(reg63))
            begin
              reg77 <= ((-(reg65 <<< reg74)) & (((((7'h49) << reg67) <<< forvar56) ?
                  reg55 : $unsigned(reg45)) >>> wire41[(1'h0):(1'h0)]));
              reg78 = (wire37 ?
                  $unsigned((^$signed((reg64 ^~ reg64)))) : wire38[(5'h12):(3'h7)]);
              reg79 <= $signed($signed(($unsigned(((7'h4a) ?
                      forvar57 : reg43)) ?
                  ($unsigned(reg73) ^~ (reg62 & reg58)) : forvar57[(2'h2):(1'h1)])));
              reg80 <= ((!reg67[(5'h11):(1'h0)]) ?
                  ((|((reg50 ? reg77 : wire38) > {wire40, reg55})) ?
                      (+($unsigned(reg75) < $signed(reg76))) : (((reg43 ~^ reg79) ?
                              reg65[(1'h1):(1'h0)] : (reg60 ? reg64 : reg74)) ?
                          reg61 : (^~reg74[(2'h3):(2'h3)]))) : reg62[(1'h0):(1'h0)]);
              reg81 = $unsigned(reg73);
            end
          else
            begin
              reg78 = $unsigned(forvar56[(4'h8):(3'h7)]);
              reg81 = {($unsigned($signed(forvar57)) ?
                      (($unsigned((8'hbd)) ^ $unsigned(reg66)) * reg60[(5'h11):(4'he)]) : (~&reg63))};
              reg82 = reg54;
              reg83 = ((!reg82) ?
                  (-reg67) : ((^((reg66 ? reg64 : reg74) ?
                          $signed(reg74) : reg74)) ?
                      wire40 : (-$signed((forvar72 ? reg70 : wire39)))));
            end
        end
      else
        begin
          for (forvar71 = (1'h0); (forvar71 < (2'h2)); forvar71 = (forvar71 + (1'h1)))
            begin
              reg72 <= $unsigned(reg80);
              reg73 = reg63;
              reg74 <= (!reg83);
              reg75 = reg61;
              reg77 <= $unsigned((reg63[(4'hc):(2'h2)] >= {(~|$signed(reg50))}));
            end
          reg79 <= reg82;
          reg81 = $unsigned((reg52[(3'h6):(3'h5)] >= {((reg71 ?
                      (8'hb7) : reg80) ?
                  reg65[(3'h4):(3'h4)] : (forvar71 <<< (8'ha1))),
              $signed(reg59)}));
          reg82 = reg63[(4'hd):(3'h5)];
          for (forvar83 = (1'h0); (forvar83 < (2'h2)); forvar83 = (forvar83 + (1'h1)))
            begin
              reg84 = ($signed($signed(wire37)) ~^ (reg62[(1'h1):(1'h0)] ?
                  forvar71 : $signed($signed($signed(reg72)))));
              reg85 = {(forvar71 << $unsigned(((~|(8'hba)) ?
                      {forvar56} : wire39[(3'h6):(1'h0)])))};
            end
        end
    end
  assign wire86 = wire53;
  module87 #() modinst820 (.y(wire819), .wire90(reg61), .wire91(reg68), .clk(clk), .wire89(wire40), .wire88(wire86));
  always
    @(posedge clk) begin
      reg821 = (~$signed(reg72[(2'h3):(2'h2)]));
      reg822 = $unsigned((reg61 > $unsigned({$signed(reg59)})));
      if (reg64[(4'hb):(3'h7)])
        begin
          for (forvar823 = (1'h0); (forvar823 < (2'h2)); forvar823 = (forvar823 + (1'h1)))
            begin
              reg824 <= (8'ha7);
              reg825 = $signed((~&reg43[(4'hc):(4'h8)]));
              reg826 = reg50;
            end
          for (forvar827 = (1'h0); (forvar827 < (1'h1)); forvar827 = (forvar827 + (1'h1)))
            begin
              reg828 <= reg58[(5'h14):(5'h14)];
              reg829 = (((reg68[(4'h9):(2'h3)] ?
                      ((!(8'haa)) * $unsigned(reg60)) : ((reg59 ?
                          forvar827 : wire36) + (&(7'h40)))) ?
                  $unsigned(reg77) : reg77[(4'hc):(1'h1)]) + $signed($unsigned(({(7'h49),
                      wire38} ?
                  (reg50 ? (8'ha2) : reg63) : $signed(wire53)))));
              reg830 <= ((wire86 != reg72[(4'h9):(3'h4)]) + ($unsigned(reg829) ?
                  (((8'hbf) ?
                      (&(8'ha6)) : $signed(forvar827)) >>> (reg45[(2'h3):(2'h3)] ?
                      (7'h41) : (wire36 + reg828))) : $signed((+(^wire39)))));
              reg831 = (reg58[(3'h6):(1'h1)] ?
                  $signed(((reg63[(1'h1):(1'h1)] ^ (wire819 != reg826)) && reg59)) : reg80[(4'h9):(2'h2)]);
            end
        end
      else
        begin
          reg823 <= ((8'had) ^ $signed(reg79[(3'h4):(1'h0)]));
          reg824 <= ((|(8'hab)) && {$unsigned((-(reg55 - reg52))),
              (+$unsigned((-reg830)))});
          if (($unsigned(((&$unsigned(reg50)) <= $unsigned((wire36 ?
                  reg63 : wire37)))) ?
              (&$signed(wire36[(4'hc):(3'h7)])) : ((((reg80 ?
                      reg72 : (8'had)) * $signed(reg58)) != (~^$unsigned(reg830))) ?
                  reg43 : ($unsigned($unsigned((8'hb0))) ?
                      reg822[(4'hc):(2'h2)] : (-reg65)))))
            begin
              reg827 <= $signed(reg58[(3'h6):(2'h2)]);
              reg829 = ($unsigned(reg77[(4'hf):(3'h7)]) >= $unsigned(wire86[(3'h4):(1'h1)]));
              reg830 <= reg63;
              reg831 = ((-$unsigned($signed(reg61[(3'h4):(2'h3)]))) ?
                  ({{(wire37 <= reg79), (reg43 - wire38)}} ?
                      ((|$unsigned(reg74)) > reg80[(4'ha):(3'h4)]) : (|$unsigned(wire37))) : $unsigned(({(^~reg72)} ?
                      ($signed(reg824) ?
                          reg821 : $signed(reg58)) : {wire53[(3'h4):(3'h4)],
                          (forvar823 ? (7'h46) : reg58)})));
              reg832 = $signed((forvar823[(1'h1):(1'h1)] != reg72));
            end
          else
            begin
              reg827 <= $unsigned($unsigned(((~|(reg45 << reg59)) ?
                  (~&$signed(wire38)) : {reg828[(4'h9):(1'h0)]})));
              reg828 <= {$signed((~$signed(reg58)))};
            end
        end
      reg833 <= ((reg52[(2'h2):(1'h1)] ?
              ((wire40[(4'h8):(1'h0)] | reg70) >= $signed({reg68})) : $unsigned(wire41[(2'h2):(1'h1)])) ?
          $unsigned({{reg68, $signed(reg55)},
              (~$signed(wire37))}) : {(((reg828 ? reg822 : reg58) ?
                      ((8'hac) ? wire37 : reg832) : (-reg830)) ?
                  reg825 : reg824[(1'h0):(1'h0)]),
              (((wire37 ?
                  wire39 : reg72) ~^ (~&reg68)) == wire41[(2'h3):(1'h1)])});
    end
  assign wire834 = ($signed((|reg43[(1'h1):(1'h1)])) ?
                       $signed(((reg45 ^~ reg59[(1'h1):(1'h1)]) ?
                           reg55 : $signed((reg61 && (8'ha4))))) : $signed(wire40[(3'h5):(2'h2)]));
  always
    @(posedge clk) begin
      if ((wire53 ?
          reg827 : ((reg833 ?
              {(reg55 < reg72),
                  $signed(wire36)} : reg80[(1'h0):(1'h0)]) && (+(wire40 ?
              (reg55 ? reg823 : reg823) : $signed(wire53))))))
        begin
          reg835 <= ((~($unsigned(reg64[(2'h2):(2'h2)]) | (wire38[(3'h4):(2'h2)] - (~^wire40)))) ?
              $unsigned(($signed({wire86, (7'h41)}) ?
                  wire39 : reg70[(4'hf):(4'h9)])) : $signed($signed((8'hab))));
          for (forvar836 = (1'h0); (forvar836 < (1'h1)); forvar836 = (forvar836 + (1'h1)))
            begin
              reg837 <= $unsigned({(!({(8'hbe)} ?
                      reg45 : (reg52 ? reg77 : (8'h9c)))),
                  reg828});
              reg838 = $signed((reg45[(3'h6):(2'h2)] - (7'h40)));
              reg839 = (!(|(|$unsigned((reg70 ? reg61 : wire819)))));
            end
          reg840 = (8'ha6);
        end
      else
        begin
          reg836 = $unsigned(wire40[(2'h3):(2'h2)]);
          for (forvar837 = (1'h0); (forvar837 < (1'h1)); forvar837 = (forvar837 + (1'h1)))
            begin
              reg838 = $unsigned($unsigned(wire819[(2'h2):(2'h2)]));
              reg841 <= reg839;
              reg842 = $unsigned(wire39[(3'h5):(3'h4)]);
              reg843 = reg840;
              reg844 = $signed((wire41[(1'h0):(1'h0)] ? (7'h42) : forvar837));
            end
          for (forvar845 = (1'h0); (forvar845 < (1'h0)); forvar845 = (forvar845 + (1'h1)))
            begin
              reg846 <= (~$unsigned($signed((8'hb4))));
              reg847 <= ((reg64 > reg59[(1'h0):(1'h0)]) < $unsigned(($unsigned(((8'hb8) || (8'hbb))) ?
                  $signed($unsigned(reg843)) : $signed(reg823[(3'h4):(3'h4)]))));
            end
          if ((reg837[(3'h6):(1'h0)] >>> (reg844 >= ((-reg840) ?
              reg60 : $signed((reg79 ? wire39 : wire86))))))
            begin
              reg848 = (($signed((~|$unsigned(reg43))) || reg58) ?
                  $signed((((reg837 <<< (8'hbe)) ?
                      reg833[(1'h1):(1'h1)] : (!reg830)) <<< ((reg847 >> reg839) ?
                      (|reg59) : wire36))) : $unsigned((($unsigned(reg840) <<< reg823) ?
                      (reg68[(2'h2):(2'h2)] ?
                          ((8'hb3) ? reg65 : reg68) : (forvar837 ?
                              reg61 : reg70)) : $unsigned($unsigned(wire834)))));
              reg849 = $unsigned(reg830[(4'hb):(3'h7)]);
              reg850 <= ({$unsigned($unsigned(reg65))} | $unsigned((^~$signed(wire86[(1'h1):(1'h0)]))));
              reg851 <= ((reg52[(1'h1):(1'h1)] ?
                  $unsigned($unsigned(reg59[(2'h2):(2'h2)])) : (((reg50 != reg824) ?
                      (reg80 < reg74) : {wire39,
                          (8'hb9)}) >>> (~^$signed(wire819)))) - $signed($unsigned(((-reg60) ?
                  (reg844 != reg840) : forvar836))));
            end
          else
            begin
              reg848 = forvar845;
            end
        end
      reg852 = $unsigned((&{($signed(reg61) ?
              ((7'h45) ? (8'hbb) : reg851) : $unsigned(reg63)),
          wire41}));
    end
  assign wire853 = (wire41 ? $signed(wire819[(1'h1):(1'h0)]) : reg59);
  assign wire854 = (($unsigned((!{reg60,
                       reg847})) <<< $unsigned(reg828[(4'he):(2'h3)])) & (&($signed($unsigned(wire819)) >>> $signed(reg851))));
  always
    @(posedge clk) begin
      if ($signed(reg823))
        begin
          if (($unsigned((7'h47)) <= reg63))
            begin
              reg855 <= $signed(reg827);
              reg856 <= ({(({reg55} && (wire39 ? reg52 : reg855)) ?
                          $unsigned(reg60) : $unsigned(reg72)),
                      (($unsigned(reg827) * reg50[(3'h4):(1'h1)]) ?
                          reg855[(1'h0):(1'h0)] : $signed((reg58 ?
                              reg851 : reg74)))} ?
                  ($unsigned((~^(reg43 ?
                      reg828 : reg59))) >= {reg58[(4'hd):(4'h9)]}) : (((|(reg837 >> wire853)) & (reg833 ?
                          (reg847 ? reg60 : wire41) : reg74[(3'h7):(2'h2)])) ?
                      reg63 : ($unsigned(wire41) & (reg79 ?
                          $signed(reg60) : (reg828 ? wire40 : reg61)))));
              reg857 <= (^{$unsigned((~|$unsigned(reg72))),
                  ((^~(wire36 ? reg72 : (8'hb6))) ?
                      $signed({reg65, reg55}) : (((8'h9e) >>> reg45) ?
                          reg827 : $unsigned(reg50)))});
              reg858 <= reg835;
            end
          else
            begin
              reg855 <= ({$signed(wire86[(4'hb):(4'hb)])} ?
                  wire37[(4'h8):(1'h1)] : $signed({reg64[(4'h9):(3'h6)]}));
              reg856 <= (|(|{$signed(reg830), (^~(!wire853))}));
            end
        end
      else
        begin
          if ($unsigned(((((8'h9f) >= $signed(reg65)) | (reg857 | (wire39 ~^ reg856))) ?
              reg68 : reg59)))
            begin
              reg859 = $signed((reg858 >> wire37[(1'h1):(1'h0)]));
            end
          else
            begin
              reg859 = wire39[(3'h4):(1'h1)];
              reg860 = {(($unsigned(reg45[(1'h1):(1'h1)]) ?
                      ((|reg65) ^~ $signed((7'h49))) : ($unsigned(reg45) ?
                          $signed((8'hb3)) : (reg837 << reg72))) != (((reg59 <= (8'hbf)) ?
                          reg59[(1'h1):(1'h1)] : reg58) ?
                      (reg824 ?
                          $signed(reg64) : reg856[(4'hf):(4'he)]) : ($unsigned(reg55) >>> (reg58 || (8'hb4)))))};
              reg861 = (&wire853);
              reg862 <= (((~&{reg52[(3'h4):(2'h2)]}) ?
                  reg74 : wire834[(3'h6):(1'h1)]) ^ ({$signed((reg837 << reg64))} ?
                  $unsigned((8'hb9)) : reg52[(1'h1):(1'h1)]));
              reg863 = $signed((~|reg857[(2'h3):(1'h0)]));
            end
          reg864 <= wire853;
        end
      if (reg846[(3'h5):(3'h4)])
        begin
          if ((+reg862[(4'h8):(3'h4)]))
            begin
              reg865 = ($signed((^~$unsigned((&reg52)))) ?
                  reg857 : $signed({wire834}));
              reg866 = wire39[(1'h0):(1'h0)];
              reg867 <= (reg857 || reg60[(5'h11):(4'he)]);
              reg868 <= reg837;
            end
          else
            begin
              reg867 <= $signed($signed((reg59 >> (reg850[(4'h9):(3'h4)] ?
                  $signed(reg860) : reg862[(2'h3):(1'h1)]))));
              reg869 = $unsigned((reg80[(3'h7):(3'h5)] ?
                  reg833[(3'h4):(3'h4)] : $signed(((reg828 == reg855) ?
                      $unsigned(reg827) : reg79))));
              reg870 <= {reg50};
              reg871 <= reg65[(2'h2):(1'h1)];
            end
          reg872 <= wire854;
          reg873 <= ((reg865[(1'h0):(1'h0)] ?
                  reg64[(4'h8):(3'h4)] : reg861[(3'h4):(2'h3)]) ?
              (reg860 ?
                  $signed($unsigned((~&reg72))) : ($unsigned((reg59 && reg824)) < $unsigned(reg861[(3'h5):(1'h0)]))) : reg872[(4'h9):(3'h6)]);
        end
      else
        begin
          reg867 <= reg828;
        end
    end
  always
    @(posedge clk) begin
      for (forvar874 = (1'h0); (forvar874 < (2'h2)); forvar874 = (forvar874 + (1'h1)))
        begin
          reg875 <= $signed(wire36[(4'h9):(2'h2)]);
          for (forvar876 = (1'h0); (forvar876 < (2'h2)); forvar876 = (forvar876 + (1'h1)))
            begin
              reg877 <= (7'h42);
            end
          for (forvar878 = (1'h0); (forvar878 < (2'h2)); forvar878 = (forvar878 + (1'h1)))
            begin
              reg879 = (wire41[(1'h0):(1'h0)] ?
                  (((-(~&reg60)) ?
                      reg828[(2'h2):(2'h2)] : {reg45[(3'h4):(1'h0)],
                          $unsigned(reg875)}) & (~|(reg851 ?
                      ((8'hb5) ~^ reg52) : reg870))) : (($unsigned($unsigned((7'h48))) >>> (8'ha3)) < wire834[(4'he):(3'h6)]));
            end
          for (forvar880 = (1'h0); (forvar880 < (3'h4)); forvar880 = (forvar880 + (1'h1)))
            begin
              reg881 = ($signed(($signed((reg851 > reg858)) | {$signed(reg873),
                      reg74[(2'h2):(1'h1)]})) ?
                  (~|wire86[(4'h9):(4'h9)]) : {(((reg72 >= reg858) ?
                              {forvar876, reg862} : $signed(reg79)) ?
                          wire38 : ((-reg858) >= $unsigned(wire86))),
                      ((&(reg60 ? reg875 : reg828)) & wire53)});
              reg882 = (!(-(((8'hb3) ?
                  reg60[(1'h0):(1'h0)] : $signed(reg851)) + ((wire53 ?
                  wire37 : reg827) == (reg875 > wire36)))));
              reg883 <= ((|(~{wire853[(1'h0):(1'h0)], reg63})) && reg65);
              reg884 = reg58[(5'h14):(4'h8)];
              reg885 <= $signed($signed(reg872));
            end
          if (reg877)
            begin
              reg886 <= (reg862[(4'h9):(4'h9)] ~^ reg828[(4'h8):(4'h8)]);
              reg887 <= (7'h40);
              reg888 = (~^$unsigned(((~|wire38[(3'h5):(1'h1)]) ?
                  (^~(~(8'hb2))) : ({reg58} ? {reg827, wire834} : {reg65}))));
              reg889 = $signed(reg847[(1'h1):(1'h1)]);
            end
          else
            begin
              reg888 = $signed((&reg74));
              reg890 <= $signed((|reg823[(4'hb):(3'h5)]));
              reg891 = $unsigned(((wire40 ?
                  $unsigned(reg886) : reg60) ~^ ((reg835[(5'h14):(1'h1)] ?
                      $unsigned(reg855) : reg867[(1'h0):(1'h0)]) ?
                  (reg45[(3'h4):(1'h1)] > (^~reg862)) : {{reg72, reg43},
                      (-reg79)})));
              reg892 <= reg871[(3'h6):(2'h3)];
              reg893 = $unsigned($signed((wire39 ?
                  reg855[(4'h8):(1'h1)] : (-(reg871 > reg68)))));
            end
        end
      if ($unsigned(reg890))
        begin
          if ((($unsigned({reg68, reg45}) ?
                  reg881[(3'h7):(1'h0)] : ($unsigned((reg862 ?
                      reg61 : (7'h47))) || (reg80[(4'h8):(1'h1)] * {reg824,
                      reg55}))) ?
              reg881 : (8'hbc)))
            begin
              reg894 = ((~&$signed(reg886[(3'h6):(3'h5)])) >>> $unsigned(($unsigned((reg827 ?
                  reg864 : reg59)) > wire853)));
            end
          else
            begin
              reg895 <= ((&$signed(($unsigned(wire39) & (^reg887)))) ~^ ({((reg864 <= reg79) ?
                      reg68[(1'h1):(1'h0)] : reg886[(3'h5):(1'h1)]),
                  (&reg888)} <= $unsigned((-$unsigned((8'hae))))));
              reg896 <= {forvar878[(2'h2):(2'h2)], (8'hb7)};
              reg897 <= ({($unsigned($signed(reg873)) ?
                          $unsigned((reg61 ?
                              reg857 : forvar880)) : $unsigned($signed(reg45)))} ?
                  $unsigned({reg864}) : wire40);
              reg898 = (($unsigned(reg892) ?
                      ({$signed((8'hb9)), reg879} < ((~reg55) ?
                          {reg889} : (reg68 ?
                              reg43 : reg895))) : $unsigned($signed((reg827 ?
                          (7'h49) : reg830)))) ?
                  (~|$unsigned($unsigned(reg887[(2'h3):(1'h0)]))) : $unsigned(($signed($unsigned(wire854)) + $unsigned($unsigned(wire819)))));
              reg899 = ((&(forvar878[(3'h7):(2'h3)] * (|(wire41 < wire41)))) ?
                  $unsigned((|wire53)) : $unsigned(reg864[(4'h9):(2'h3)]));
            end
          for (forvar900 = (1'h0); (forvar900 < (2'h2)); forvar900 = (forvar900 + (1'h1)))
            begin
              reg901 <= {wire819, reg846};
              reg902 = $signed(reg828[(4'hc):(3'h6)]);
              reg903 = $signed($signed((((|(7'h42)) ^ $signed(reg58)) ?
                  $signed(reg74) : (-$signed(wire38)))));
              reg904 <= $signed(reg890[(4'hc):(2'h2)]);
              reg905 <= reg879[(1'h1):(1'h1)];
            end
          for (forvar906 = (1'h0); (forvar906 < (3'h4)); forvar906 = (forvar906 + (1'h1)))
            begin
              reg907 = reg60;
            end
          reg908 <= reg877[(4'ha):(1'h0)];
          reg909 <= reg898[(1'h0):(1'h0)];
        end
      else
        begin
          if (($signed((8'hb1)) ?
              $unsigned($unsigned(reg79[(3'h4):(2'h3)])) : reg827[(4'he):(3'h4)]))
            begin
              reg895 <= ((8'h9c) ?
                  $unsigned($unsigned((|(reg871 ?
                      forvar878 : reg902)))) : $signed((!(wire53[(3'h5):(1'h0)] ?
                      (-wire53) : (reg873 ? reg875 : reg847)))));
              reg896 <= reg855[(1'h0):(1'h0)];
              reg897 <= $signed($unsigned({({reg80} ?
                      $signed((8'ha5)) : $signed(forvar880)),
                  $signed(((8'ha3) ? forvar880 : reg61))}));
              reg900 <= forvar900[(1'h1):(1'h0)];
            end
          else
            begin
              reg894 = {$unsigned((~wire86[(4'hb):(4'ha)]))};
              reg895 <= $unsigned((reg58 > $unsigned(reg846[(3'h4):(2'h3)])));
            end
          if (({($signed(reg72) << $unsigned(reg899[(3'h6):(2'h3)]))} ?
              forvar876[(2'h2):(1'h0)] : (7'h4a)))
            begin
              reg902 = (8'hb6);
              reg904 <= ((((8'ha2) ? reg904 : (+(reg59 || (7'h46)))) ?
                  reg72[(3'h7):(3'h6)] : {$unsigned(reg862)}) || (|{($signed((8'hb4)) < reg875[(3'h6):(1'h1)])}));
              reg906 = wire53;
            end
          else
            begin
              reg901 <= wire853;
              reg902 = {($signed($unsigned($unsigned(forvar878))) >> (((reg45 < reg884) * $unsigned(forvar906)) <= $unsigned($signed((7'h4a))))),
                  $unsigned((wire36[(3'h6):(1'h1)] && ($signed(reg43) ?
                      {reg888} : {reg900, reg886})))};
              reg904 <= (((wire86 ?
                  $unsigned(wire40) : {(reg835 >>> (8'hb8))}) * (~|$signed(reg872))) <<< ((({reg887,
                      reg898} ?
                  reg850[(1'h1):(1'h1)] : $signed((8'hb4))) ^~ $signed((reg60 << reg847))) << (reg885[(3'h5):(2'h3)] <= $unsigned($signed(forvar880)))));
              reg905 <= reg50[(1'h1):(1'h0)];
            end
          for (forvar907 = (1'h0); (forvar907 < (1'h0)); forvar907 = (forvar907 + (1'h1)))
            begin
              reg910 = ({reg79, reg59} < ({({(8'ha8)} ?
                      (wire36 - wire37) : $signed(reg837)),
                  ($unsigned((8'ha8)) || (wire854 >>> wire41))} * (&(8'hb2))));
              reg911 = reg899[(4'he):(4'he)];
              reg912 <= (reg896[(4'hc):(3'h5)] | reg896[(4'hc):(2'h2)]);
            end
          reg913 <= {$unsigned(reg855),
              $unsigned($signed(reg886[(3'h5):(3'h4)]))};
          reg914 <= reg912;
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned({($unsigned($unsigned(reg877)) ?
              $signed($unsigned(reg872)) : $unsigned(reg886)),
          $signed((+(reg60 != reg70)))}))
        begin
          for (forvar915 = (1'h0); (forvar915 < (2'h2)); forvar915 = (forvar915 + (1'h1)))
            begin
              reg916 <= $signed((~|(reg43 ?
                  $unsigned((8'ha5)) : {reg868, ((8'had) * reg45)})));
            end
          reg917 <= forvar915[(1'h0):(1'h0)];
          for (forvar918 = (1'h0); (forvar918 < (1'h0)); forvar918 = (forvar918 + (1'h1)))
            begin
              reg919 = ($unsigned($signed($signed($signed(reg886)))) ^~ $unsigned((~&{(^~wire853)})));
              reg920 <= (!reg43);
              reg921 <= (reg841 < ((7'h42) ?
                  $unsigned($unsigned((reg61 >>> reg827))) : {$unsigned($unsigned(reg892)),
                      reg886[(3'h5):(2'h3)]}));
              reg922 = reg79[(3'h4):(1'h0)];
            end
          for (forvar923 = (1'h0); (forvar923 < (1'h1)); forvar923 = (forvar923 + (1'h1)))
            begin
              reg924 <= ($unsigned(reg885[(5'h11):(1'h0)]) ?
                  ((((reg850 <<< reg905) ?
                              $signed(reg896) : ((8'hab) >= reg827)) ?
                          (~^$signed(reg68)) : $signed(wire38)) ?
                      $unsigned(reg864) : ($signed(reg895) ?
                          ((reg64 ? reg45 : reg904) ?
                              (reg870 ?
                                  reg841 : wire854) : $unsigned(reg68)) : (|reg68[(4'hc):(1'h0)]))) : $unsigned(($signed(reg858[(1'h1):(1'h0)]) * ($unsigned(reg856) ^~ $signed(reg867)))));
              reg925 = $signed(reg856);
              reg926 = {reg867, wire834};
              reg927 = reg873;
            end
          reg928 = $signed($signed(reg830[(1'h0):(1'h0)]));
        end
      else
        begin
          for (forvar915 = (1'h0); (forvar915 < (2'h3)); forvar915 = (forvar915 + (1'h1)))
            begin
              reg916 <= {reg65,
                  (!{((reg919 ? reg913 : reg63) * (reg50 ? reg862 : reg45)),
                      $signed($signed(reg850))})};
            end
        end
    end
  always
    @(posedge clk) begin
      reg929 <= $signed($unsigned((^~(reg830 ? reg872 : $signed(reg875)))));
      reg930 = ($unsigned((wire41 ?
          (~|reg868[(1'h0):(1'h0)]) : (wire853[(4'h9):(2'h2)] >> (8'h9e)))) < (reg847 == (reg875[(1'h1):(1'h0)] ?
          {reg887, $signed((8'ha2))} : (+(wire86 << (8'ha0))))));
      for (forvar931 = (1'h0); (forvar931 < (1'h0)); forvar931 = (forvar931 + (1'h1)))
        begin
          reg932 = {reg887[(1'h1):(1'h1)]};
          reg933 <= (8'ha5);
          reg934 = reg932[(3'h5):(2'h2)];
          reg935 <= $unsigned(({(wire86[(3'h4):(1'h0)] << $unsigned(reg905)),
              reg60[(5'h15):(3'h5)]} - reg851[(3'h4):(1'h0)]));
        end
    end
  always
    @(posedge clk) begin
      for (forvar936 = (1'h0); (forvar936 < (2'h2)); forvar936 = (forvar936 + (1'h1)))
        begin
          for (forvar937 = (1'h0); (forvar937 < (3'h4)); forvar937 = (forvar937 + (1'h1)))
            begin
              reg938 <= (^reg55);
            end
          for (forvar939 = (1'h0); (forvar939 < (1'h0)); forvar939 = (forvar939 + (1'h1)))
            begin
              reg940 = $unsigned(reg64);
              reg941 = $unsigned((($unsigned((reg58 << reg872)) - reg855[(1'h0):(1'h0)]) + {(^$signed(wire86)),
                  (((8'h9d) || reg904) >> reg905)}));
              reg942 = $unsigned(wire53[(1'h0):(1'h0)]);
              reg943 <= $signed(reg846[(2'h2):(1'h0)]);
              reg944 = $signed(($signed(reg921) ^~ reg823));
            end
          reg945 <= $signed($unsigned(((~reg920) ?
              $unsigned(reg895[(1'h1):(1'h0)]) : ((-wire854) ?
                  reg921 : $signed(reg909)))));
          reg946 <= reg65;
          for (forvar947 = (1'h0); (forvar947 < (1'h1)); forvar947 = (forvar947 + (1'h1)))
            begin
              reg948 = (($signed((~|reg924)) >> $unsigned($signed((wire41 ?
                      reg824 : reg828)))) ?
                  $unsigned($signed($unsigned($unsigned((8'hbd))))) : $unsigned((($signed(reg924) <<< (wire38 ?
                          reg55 : reg875)) ?
                      reg52 : reg867)));
              reg949 = reg909[(5'h13):(4'h8)];
              reg950 = reg896;
              reg951 = $unsigned(($unsigned(wire53[(2'h2):(1'h0)]) ?
                  $unsigned(($unsigned((7'h47)) >= reg935)) : reg77[(2'h2):(2'h2)]));
            end
        end
      reg952 <= (reg830[(1'h0):(1'h0)] >= $unsigned({(reg80 ?
              (reg938 + reg945) : {reg950})}));
      reg953 = $unsigned($unsigned($signed((8'ha4))));
      if (($signed(forvar936) ?
          ({reg896, $signed($signed(wire53))} ?
              $signed(({reg942} ?
                  reg58[(5'h14):(1'h0)] : forvar936)) : $signed(reg873)) : $signed(((!reg900) >> reg65))))
        begin
          for (forvar954 = (1'h0); (forvar954 < (2'h2)); forvar954 = (forvar954 + (1'h1)))
            begin
              reg955 = {$signed(($unsigned($signed(reg952)) ?
                      (7'h49) : $signed({reg833, wire39})))};
              reg956 <= reg824;
            end
          if (($unsigned(reg948) == (~&reg933)))
            begin
              reg957 <= {(-reg905[(4'hb):(1'h0)])};
              reg958 <= ((|reg952[(4'hd):(3'h6)]) ?
                  (reg875 ?
                      reg846 : ((-(reg943 || reg875)) ?
                          (+(8'ha5)) : (!$signed(reg904)))) : {$unsigned((reg846[(3'h5):(2'h3)] ?
                          {reg45, wire41} : $unsigned(reg914)))});
            end
          else
            begin
              reg957 <= ($unsigned(wire53) ?
                  $unsigned($signed(reg935[(3'h6):(3'h5)])) : $unsigned(({$unsigned(reg941)} ?
                      (&reg944[(2'h2):(1'h0)]) : $unsigned(reg944[(1'h1):(1'h1)]))));
              reg958 <= $unsigned(reg846[(2'h3):(2'h2)]);
            end
        end
      else
        begin
          reg954 = reg949[(5'h12):(3'h6)];
          for (forvar955 = (1'h0); (forvar955 < (2'h3)); forvar955 = (forvar955 + (1'h1)))
            begin
              reg956 <= $unsigned(((wire53 ?
                      wire38[(5'h17):(4'h9)] : $signed({reg951})) ?
                  (^~forvar947[(4'h9):(2'h2)]) : $unsigned(((reg873 | reg873) ?
                      (|reg68) : ((7'h40) + reg904)))));
              reg959 = reg61;
              reg960 <= reg52;
              reg961 = (reg945[(4'ha):(3'h5)] ?
                  $signed($unsigned(reg943[(3'h5):(1'h0)])) : (((~^$unsigned((8'hbb))) <<< $signed($unsigned(reg957))) && ({(reg952 ?
                              (8'h9d) : reg883),
                          (8'ha7)} ?
                      $signed((^~(8'hb6))) : (&$signed(forvar947)))));
            end
          reg962 <= {$unsigned($unsigned(wire854)),
              $unsigned($signed(((reg74 != reg846) ?
                  reg957[(3'h4):(2'h3)] : $unsigned(reg80))))};
        end
      reg963 = (((wire53[(3'h4):(2'h2)] | $signed((~^reg72))) & reg949) * $signed((-reg61[(1'h0):(1'h0)])));
    end
  always
    @(posedge clk) begin
      if ((|$signed((+(&(~reg890))))))
        begin
          for (forvar964 = (1'h0); (forvar964 < (1'h1)); forvar964 = (forvar964 + (1'h1)))
            begin
              reg965 = wire36;
              reg966 = reg43;
              reg967 = (^((({reg824, (7'h45)} ?
                          reg883[(4'he):(2'h2)] : reg846) ?
                      reg77[(5'h10):(4'h8)] : $signed((reg72 ?
                          reg837 : reg823))) ?
                  (reg877 ? $unsigned((~^reg841)) : $signed(reg55)) : reg61));
            end
          reg968 <= (~|wire38[(5'h14):(4'h8)]);
          if (wire41[(1'h1):(1'h0)])
            begin
              reg969 <= ((&reg61) >= {reg830});
              reg970 <= $signed({(reg933 ?
                      (reg875 - (reg862 ? reg70 : reg871)) : $unsigned((reg74 ?
                          wire38 : wire38)))});
              reg971 <= reg877;
            end
          else
            begin
              reg972 = reg872;
              reg973 <= ((reg952 ?
                      (((reg943 ~^ reg952) == reg858[(1'h1):(1'h1)]) ?
                          (^$unsigned(reg886)) : $unsigned(((8'hbc) ^ wire40))) : reg830) ?
                  $unsigned($signed(($signed(reg877) ?
                      {reg68} : {reg830, reg862}))) : reg77[(5'h11):(3'h7)]);
            end
        end
      else
        begin
          for (forvar964 = (1'h0); (forvar964 < (2'h3)); forvar964 = (forvar964 + (1'h1)))
            begin
              reg965 = {$signed((reg887[(3'h7):(3'h7)] ?
                      reg945 : $signed((reg969 >= reg873))))};
              reg966 = ($unsigned((({reg63,
                  (8'ha6)} >= $unsigned(wire86)) << $signed((reg921 > reg946)))) <= $unsigned(($signed(((8'ha3) <= reg68)) ?
                  {(-reg967)} : $signed({reg64}))));
              reg968 <= (reg962[(4'h9):(1'h0)] ?
                  (~|($unsigned((reg74 ^~ reg968)) <= $signed((^~(8'hbe))))) : $unsigned((~(reg890[(4'hc):(4'ha)] ?
                      (~^reg80) : reg828[(1'h1):(1'h1)]))));
              reg969 <= (~(($unsigned((~reg916)) ^~ $unsigned((reg887 | (8'ha5)))) ?
                  reg68[(4'hc):(4'h9)] : ($signed({reg966}) ?
                      (|(!reg970)) : reg938[(2'h3):(2'h3)])));
            end
          reg972 = (8'hb5);
          for (forvar973 = (1'h0); (forvar973 < (3'h4)); forvar973 = (forvar973 + (1'h1)))
            begin
              reg974 = $unsigned(($unsigned(reg59[(2'h2):(2'h2)]) > (((reg873 ?
                      reg920 : reg55) ?
                  reg45 : $unsigned(reg905)) - reg921)));
              reg975 <= (+(reg966 ^ {reg883[(4'h9):(3'h5)],
                  $signed((|(8'haa)))}));
              reg976 = (reg851 ?
                  (^((reg841 && $unsigned((7'h47))) ?
                      (^~{reg974,
                          reg858}) : $unsigned($unsigned((8'hbd))))) : ((reg952 ?
                          (-{reg43, reg868}) : ((~^reg862) >>> (reg887 ?
                              reg827 : forvar973))) ?
                      $signed((8'haf)) : ($signed(reg969) ?
                          reg850[(4'h8):(3'h6)] : $unsigned(reg64[(4'ha):(1'h1)]))));
              reg977 <= (reg61 ? wire53 : $unsigned(reg887));
            end
          for (forvar978 = (1'h0); (forvar978 < (1'h1)); forvar978 = (forvar978 + (1'h1)))
            begin
              reg979 <= {(($unsigned($signed((8'hb3))) << (~(~reg50))) < (($signed(reg929) <= (^(8'hb9))) ~^ reg935))};
              reg980 <= (&(8'hbb));
            end
          reg981 = wire819[(1'h0):(1'h0)];
        end
      if ($signed(($signed($unsigned(reg870)) ?
          (-$unsigned((^~reg833))) : reg895[(3'h4):(2'h3)])))
        begin
          if ({$signed(reg952[(4'h9):(1'h1)])})
            begin
              reg982 = ($signed($unsigned((reg921[(1'h0):(1'h0)] - reg72))) ?
                  $signed($unsigned(reg921)) : $signed(reg877[(1'h1):(1'h0)]));
            end
          else
            begin
              reg983 <= (~^$signed($signed($unsigned((&(8'hab))))));
            end
          if ($unsigned(({($signed(reg970) ?
                      (reg969 <= reg956) : ((7'h41) + (7'h42))),
                  $signed({(8'hb8)})} ?
              {(~|$unsigned(reg856)),
                  ($unsigned(reg945) ~^ $unsigned((8'hbc)))} : reg921)))
            begin
              reg984 <= reg883[(2'h2):(1'h1)];
              reg985 <= $signed((~|$unsigned($unsigned($signed(reg895)))));
              reg986 = (wire854 ?
                  reg985 : $unsigned((^~(reg61 ?
                      (reg945 <<< (8'hbf)) : $unsigned(wire53)))));
              reg987 = reg77;
            end
          else
            begin
              reg984 <= $unsigned(reg901[(5'h11):(1'h1)]);
              reg986 = ((reg833[(1'h1):(1'h1)] == (((reg979 - reg969) ?
                      (+reg901) : {wire53}) >= $unsigned(reg980[(3'h4):(2'h3)]))) ?
                  (reg929 ?
                      $unsigned(reg968) : ((reg985[(4'hf):(4'h9)] ?
                          {reg967} : reg969[(2'h2):(1'h1)]) ~^ {reg833[(3'h7):(2'h3)],
                          {reg973, reg867}})) : reg938);
              reg988 <= $unsigned(reg985[(2'h3):(2'h3)]);
              reg989 = reg897;
            end
        end
      else
        begin
          if (reg980[(4'hd):(3'h4)])
            begin
              reg982 = (reg887[(3'h7):(3'h7)] & reg920);
              reg983 <= reg886;
              reg984 <= reg908;
              reg986 = (^(reg921 ?
                  $unsigned($signed((reg870 && reg80))) : ($unsigned($signed(reg920)) != $signed(reg80[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg983 <= (reg914 == reg984);
            end
          if ($signed((8'ha7)))
            begin
              reg987 = reg980;
              reg989 = reg870;
              reg990 = reg979[(3'h6):(2'h3)];
              reg991 = ({(!reg924),
                  ({reg952, reg935[(5'h13):(3'h6)]} ?
                      (^(wire38 << reg59)) : wire41[(1'h1):(1'h0)])} ~^ {(+(|(~&(7'h45)))),
                  reg870[(1'h0):(1'h0)]});
              reg992 = $signed(($unsigned((8'ha0)) >> ({(reg883 >>> (8'ha9)),
                      $signed(reg886)} ?
                  {$unsigned(reg912),
                      wire86[(3'h5):(3'h4)]} : ($unsigned((8'hab)) & $unsigned(reg972)))));
            end
          else
            begin
              reg987 = ($signed((({reg43} ^~ (reg823 ? wire819 : (8'haa))) ?
                      reg912 : wire39)) ?
                  reg835[(4'hc):(3'h6)] : ($signed(((!reg908) ?
                          (reg913 ? reg858 : wire38) : reg913)) ?
                      $signed((~&(forvar978 ^~ reg883))) : reg992));
              reg989 = $signed(({(-(reg55 == reg63)),
                  ($unsigned((8'ha4)) == reg958[(4'hb):(3'h4)])} * reg55));
              reg990 = ((&$signed(((reg984 ? reg929 : reg987) - (&wire819)))) ?
                  reg914[(4'he):(3'h5)] : reg975);
              reg993 <= (reg988 ?
                  reg962 : $unsigned($unsigned($signed((reg68 || reg856)))));
              reg994 = {$unsigned($unsigned($unsigned($signed((7'h49)))))};
            end
        end
      reg995 <= (reg895 ?
          ($signed(({reg935, wire38} == reg981[(1'h0):(1'h0)])) ?
              ((&(~reg901)) < $unsigned((8'hbb))) : $signed(reg857)) : reg864[(4'ha):(4'ha)]);
      reg996 = (!$unsigned(((8'ha2) ?
          $unsigned($signed(reg827)) : reg924[(2'h2):(1'h0)])));
    end
  always
    @(posedge clk) begin
      if (((reg909[(3'h6):(3'h5)] ? (~&wire854[(5'h13):(3'h4)]) : wire36) ?
          reg900[(4'hd):(3'h5)] : reg823))
        begin
          if (($signed($signed($signed(((8'ha4) ?
              (8'hbf) : reg908)))) >= wire39))
            begin
              reg997 = $signed($unsigned((reg960 ^~ $signed(reg871))));
              reg998 = ($signed(reg877) ?
                  $unsigned(wire38[(5'h16):(3'h7)]) : ($signed((~^(reg79 ?
                          reg924 : reg912))) ?
                      (-reg858) : reg846[(2'h2):(2'h2)]));
            end
          else
            begin
              reg999 <= (reg823[(4'h8):(3'h5)] ? reg984[(3'h4):(1'h0)] : reg79);
              reg1000 <= $signed((^~($signed(reg55[(2'h2):(1'h0)]) && reg79[(2'h3):(1'h0)])));
            end
          reg1001 <= ((~|reg909[(4'h8):(3'h5)]) | $signed($signed((reg960 <<< {wire40}))));
          reg1002 <= {reg938, reg855[(1'h1):(1'h0)]};
          if ($signed({((reg914[(4'he):(4'h9)] - (reg823 & reg909)) & $unsigned((reg921 >= reg850)))}))
            begin
              reg1003 <= reg824[(1'h1):(1'h1)];
              reg1004 = $unsigned(reg877);
              reg1005 = reg61;
              reg1006 <= {(reg50[(3'h4):(2'h3)] > (8'hbe)), reg835};
            end
          else
            begin
              reg1004 = $unsigned($unsigned($signed(reg998)));
            end
        end
      else
        begin
          if (wire36)
            begin
              reg997 = (reg50[(3'h5):(2'h3)] ?
                  reg938[(1'h0):(1'h0)] : reg871[(3'h5):(1'h1)]);
            end
          else
            begin
              reg997 = (~|wire53);
              reg999 <= reg979;
              reg1000 <= (reg921[(3'h7):(3'h7)] << $signed($unsigned($unsigned(((8'ha2) ?
                  reg864 : reg896)))));
            end
          for (forvar1001 = (1'h0); (forvar1001 < (1'h0)); forvar1001 = (forvar1001 + (1'h1)))
            begin
              reg1002 <= (^(({$unsigned(reg998)} ^~ $unsigned(reg908)) ?
                  reg968[(2'h2):(1'h1)] : (8'hb0)));
              reg1003 <= (((((&reg52) >> reg58[(1'h1):(1'h0)]) >> (reg79 ?
                  reg887[(3'h6):(1'h0)] : (reg846 ?
                      reg61 : (8'ha9)))) ^~ {$unsigned((reg912 ?
                      reg64 : reg917))}) && $unsigned(($signed(reg938[(1'h1):(1'h1)]) ?
                  $unsigned((wire37 >>> reg64)) : $unsigned(reg971[(2'h3):(2'h2)]))));
              reg1006 <= (8'hb8);
              reg1007 = {reg890};
            end
          reg1008 <= ((reg980 < reg856[(4'hc):(3'h5)]) ?
              reg841 : $unsigned($signed(((-reg960) ?
                  $unsigned(reg871) : $signed(reg79)))));
        end
      reg1009 = reg55[(2'h3):(1'h0)];
    end
  always
    @(posedge clk) begin
      if (({($unsigned((reg900 ?
              (8'h9c) : (8'hb8))) < $unsigned(reg985))} << ($unsigned($signed((^reg50))) >>> ((-reg43) ?
          reg824[(2'h2):(1'h0)] : $signed((reg847 < reg835))))))
        begin
          reg1010 = {$signed($signed((~(reg60 != reg864)))), reg999};
          reg1011 = $unsigned({reg968});
          for (forvar1012 = (1'h0); (forvar1012 < (1'h1)); forvar1012 = (forvar1012 + (1'h1)))
            begin
              reg1013 = (8'hb9);
              reg1014 = reg909;
            end
          if ($unsigned(((7'h46) ? $unsigned((-(!reg1010))) : reg871)))
            begin
              reg1015 = (($unsigned((+$signed((8'hac)))) ?
                  (8'hbb) : $signed($unsigned((reg890 > reg912)))) || ({(+$unsigned(reg1010)),
                      (reg855[(3'h5):(3'h4)] ~^ reg80)} ?
                  (reg63[(5'h12):(3'h4)] ~^ {$unsigned(wire854)}) : reg837[(2'h3):(1'h0)]));
            end
          else
            begin
              reg1015 = ($signed($signed($signed($signed(reg61)))) + (^((8'ha1) == $unsigned(reg979))));
              reg1016 = $unsigned((~^wire834[(4'he):(4'h8)]));
            end
          reg1017 = ((reg856 ?
              (($unsigned(reg896) ? reg868[(3'h4):(1'h1)] : $unsigned(reg837)) ?
                  (8'hb8) : (~&{reg50})) : reg975) | ((|reg985) ?
              (reg52[(3'h5):(2'h2)] ^~ (8'had)) : $unsigned(reg867[(5'h10):(4'h9)])));
        end
      else
        begin
          reg1010 = $signed({reg968[(1'h1):(1'h0)]});
          if ((~|{wire37[(3'h7):(3'h4)]}))
            begin
              reg1012 <= ((-$unsigned(((reg1002 ?
                  reg857 : (7'h45)) >>> reg883))) * $signed((reg913 ?
                  reg938[(1'h0):(1'h0)] : ((&reg985) ?
                      (^~reg877) : reg871[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg1012 <= ($unsigned(reg905[(3'h5):(1'h0)]) | wire53[(3'h6):(1'h1)]);
              reg1013 = ($unsigned((&reg851[(3'h7):(2'h2)])) ?
                  ($signed(($signed(reg957) ?
                      {reg912} : reg64)) << (|reg1003)) : (7'h46));
              reg1014 = reg1006[(5'h14):(4'hb)];
              reg1015 = ((8'hbd) ?
                  (reg885 ?
                      $signed(reg52) : (~&($signed((8'h9f)) && (-reg850)))) : ($unsigned(reg835[(1'h1):(1'h0)]) || $signed({(reg64 ?
                          reg958 : (7'h40)),
                      reg913})));
              reg1018 <= $signed(reg904);
            end
          if (reg1000[(1'h1):(1'h0)])
            begin
              reg1019 <= (~|reg909);
              reg1020 = ({$unsigned((reg909[(5'h14):(5'h10)] ?
                          reg846[(2'h3):(2'h3)] : $signed(reg835))),
                      (~&(((7'h40) ? reg837 : wire39) < (reg80 ?
                          reg827 : reg833)))} ?
                  $signed((~((reg917 ? reg983 : wire853) ?
                      (reg827 - reg904) : (&reg883)))) : (^~($signed({reg1013,
                      reg887}) < (~(reg58 ? reg872 : reg70)))));
              reg1021 = $signed({(((~&(8'hb5)) ?
                      $signed(reg58) : wire41) >> reg908[(4'he):(2'h2)])});
            end
          else
            begin
              reg1019 <= (&{$signed({$unsigned(reg1016), (~|reg970)}),
                  $signed((~|(reg1017 * reg1020)))});
            end
        end
      reg1022 = $signed((~&reg1021[(2'h2):(1'h1)]));
      reg1023 <= (~((reg970 >> (~^reg958)) ?
          (~^(reg45[(3'h7):(3'h4)] * (&reg872))) : (wire41 ?
              (^~(reg79 && reg900)) : $signed((reg841 - (8'hb8))))));
    end
  always
    @(posedge clk) begin
      reg1024 = (reg868 != (reg74 | reg938));
    end
  assign wire1025 = wire41;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module87  (y, clk, wire88, wire89, wire90, wire91);
  output wire [(32'he52):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire88;
  input wire signed [(2'h2):(1'h0)] wire89;
  input wire [(3'h4):(1'h0)] wire90;
  input wire [(4'hc):(1'h0)] wire91;
  wire signed [(4'ha):(1'h0)] wire818;
  wire [(4'hf):(1'h0)] wire745;
  wire signed [(3'h7):(1'h0)] wire703;
  wire [(4'hb):(1'h0)] wire702;
  wire signed [(5'h17):(1'h0)] wire662;
  wire [(4'he):(1'h0)] wire651;
  wire signed [(4'hc):(1'h0)] wire649;
  wire [(4'hc):(1'h0)] wire434;
  wire signed [(2'h3):(1'h0)] wire433;
  wire signed [(5'h16):(1'h0)] wire112;
  wire signed [(2'h2):(1'h0)] wire124;
  wire [(4'h9):(1'h0)] wire216;
  wire [(5'h18):(1'h0)] wire431;
  reg [(4'ha):(1'h0)] reg807 = (1'h0);
  reg [(3'h7):(1'h0)] reg817 = (1'h0);
  reg [(5'h10):(1'h0)] reg816 = (1'h0);
  reg [(3'h4):(1'h0)] reg812 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg809 = (1'h0);
  reg [(2'h3):(1'h0)] reg806 = (1'h0);
  reg [(2'h2):(1'h0)] reg803 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg800 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg799 = (1'h0);
  reg [(5'h15):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg795 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg791 = (1'h0);
  reg [(2'h3):(1'h0)] reg788 = (1'h0);
  reg [(5'h15):(1'h0)] reg786 = (1'h0);
  reg [(5'h12):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg780 = (1'h0);
  reg [(5'h17):(1'h0)] reg779 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg776 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg773 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg772 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg770 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg767 = (1'h0);
  reg [(5'h11):(1'h0)] reg766 = (1'h0);
  reg [(4'hf):(1'h0)] reg761 = (1'h0);
  reg [(5'h18):(1'h0)] reg759 = (1'h0);
  reg [(4'hc):(1'h0)] reg758 = (1'h0);
  reg [(4'he):(1'h0)] reg750 = (1'h0);
  reg [(4'ha):(1'h0)] reg749 = (1'h0);
  reg [(3'h5):(1'h0)] reg744 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg742 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg740 = (1'h0);
  reg [(5'h12):(1'h0)] reg739 = (1'h0);
  reg [(3'h4):(1'h0)] reg734 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg733 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg732 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg730 = (1'h0);
  reg [(3'h5):(1'h0)] reg729 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg722 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg721 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg720 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg704 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg716 = (1'h0);
  reg [(3'h4):(1'h0)] reg713 = (1'h0);
  reg [(4'hf):(1'h0)] reg712 = (1'h0);
  reg [(2'h2):(1'h0)] reg711 = (1'h0);
  reg [(2'h2):(1'h0)] reg710 = (1'h0);
  reg [(4'he):(1'h0)] reg709 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg708 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg707 = (1'h0);
  reg [(4'hd):(1'h0)] reg705 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg700 = (1'h0);
  reg [(4'hf):(1'h0)] reg699 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg696 = (1'h0);
  reg [(5'h12):(1'h0)] reg695 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg694 = (1'h0);
  reg [(5'h14):(1'h0)] reg689 = (1'h0);
  reg signed [(4'he):(1'h0)] reg687 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg686 = (1'h0);
  reg [(4'h9):(1'h0)] reg684 = (1'h0);
  reg [(5'h13):(1'h0)] reg683 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg680 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg679 = (1'h0);
  reg [(3'h7):(1'h0)] reg678 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg677 = (1'h0);
  reg [(3'h6):(1'h0)] reg675 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg674 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg671 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg669 = (1'h0);
  reg [(4'he):(1'h0)] reg667 = (1'h0);
  reg [(5'h11):(1'h0)] reg664 = (1'h0);
  reg [(5'h10):(1'h0)] reg661 = (1'h0);
  reg [(4'hf):(1'h0)] reg659 = (1'h0);
  reg signed [(4'he):(1'h0)] reg657 = (1'h0);
  reg [(4'he):(1'h0)] reg653 = (1'h0);
  reg [(3'h7):(1'h0)] reg652 = (1'h0);
  reg [(5'h14):(1'h0)] reg126 = (1'h0);
  reg [(5'h16):(1'h0)] reg123 = (1'h0);
  reg [(5'h11):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg116 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg110 = (1'h0);
  reg [(5'h12):(1'h0)] reg109 = (1'h0);
  reg [(4'hb):(1'h0)] reg103 = (1'h0);
  reg [(5'h11):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg98 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg95 = (1'h0);
  reg [(3'h7):(1'h0)] reg218 = (1'h0);
  reg [(4'h9):(1'h0)] reg221 = (1'h0);
  reg [(5'h11):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg232 = (1'h0);
  reg [(5'h16):(1'h0)] reg234 = (1'h0);
  reg [(5'h14):(1'h0)] reg236 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg240 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg245 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg248 = (1'h0);
  reg [(3'h5):(1'h0)] reg253 = (1'h0);
  reg [(4'h9):(1'h0)] reg258 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg261 = (1'h0);
  reg [(5'h17):(1'h0)] reg262 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg815 = (1'h0);
  reg [(5'h18):(1'h0)] reg814 = (1'h0);
  reg [(4'hd):(1'h0)] forvar813 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg811 = (1'h0);
  reg [(5'h18):(1'h0)] reg810 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg808 = (1'h0);
  reg [(3'h4):(1'h0)] forvar807 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar805 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg804 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg802 = (1'h0);
  reg [(4'hb):(1'h0)] reg801 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg797 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar796 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg794 = (1'h0);
  reg [(4'hd):(1'h0)] reg793 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg792 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar790 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar789 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg787 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg785 = (1'h0);
  reg [(5'h10):(1'h0)] forvar784 = (1'h0);
  reg [(5'h15):(1'h0)] forvar783 = (1'h0);
  reg [(3'h6):(1'h0)] reg782 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg778 = (1'h0);
  reg [(4'hd):(1'h0)] reg777 = (1'h0);
  reg [(5'h15):(1'h0)] forvar775 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg774 = (1'h0);
  reg signed [(4'he):(1'h0)] reg771 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg769 = (1'h0);
  reg [(4'hd):(1'h0)] reg768 = (1'h0);
  reg [(4'h9):(1'h0)] reg765 = (1'h0);
  reg [(5'h12):(1'h0)] reg764 = (1'h0);
  reg [(5'h14):(1'h0)] reg763 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg762 = (1'h0);
  reg [(5'h18):(1'h0)] forvar760 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg757 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar756 = (1'h0);
  reg [(5'h15):(1'h0)] reg755 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar754 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg753 = (1'h0);
  reg [(2'h3):(1'h0)] reg752 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg751 = (1'h0);
  reg [(4'hd):(1'h0)] reg748 = (1'h0);
  reg [(5'h14):(1'h0)] forvar747 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar746 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg743 = (1'h0);
  reg [(3'h6):(1'h0)] forvar741 = (1'h0);
  reg [(4'he):(1'h0)] reg738 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg737 = (1'h0);
  reg [(4'hc):(1'h0)] reg736 = (1'h0);
  reg [(5'h10):(1'h0)] reg735 = (1'h0);
  reg [(3'h7):(1'h0)] reg731 = (1'h0);
  reg [(5'h17):(1'h0)] forvar729 = (1'h0);
  reg [(5'h17):(1'h0)] reg728 = (1'h0);
  reg [(5'h10):(1'h0)] reg727 = (1'h0);
  reg [(4'ha):(1'h0)] reg726 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg725 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg723 = (1'h0);
  reg [(4'hd):(1'h0)] reg719 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg718 = (1'h0);
  reg [(4'h9):(1'h0)] reg717 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg715 = (1'h0);
  reg [(5'h16):(1'h0)] reg714 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg706 = (1'h0);
  reg [(4'hc):(1'h0)] forvar704 = (1'h0);
  reg [(4'ha):(1'h0)] forvar686 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg701 = (1'h0);
  reg [(3'h5):(1'h0)] reg697 = (1'h0);
  reg [(4'ha):(1'h0)] reg693 = (1'h0);
  reg [(4'hd):(1'h0)] reg692 = (1'h0);
  reg [(4'hf):(1'h0)] reg691 = (1'h0);
  reg [(4'hb):(1'h0)] reg690 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg688 = (1'h0);
  reg [(3'h5):(1'h0)] reg685 = (1'h0);
  reg [(5'h18):(1'h0)] reg682 = (1'h0);
  reg [(3'h5):(1'h0)] forvar681 = (1'h0);
  reg [(5'h15):(1'h0)] reg676 = (1'h0);
  reg [(5'h13):(1'h0)] reg673 = (1'h0);
  reg [(4'hf):(1'h0)] reg672 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar670 = (1'h0);
  reg [(5'h11):(1'h0)] forvar668 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg666 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar665 = (1'h0);
  reg [(4'he):(1'h0)] reg663 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg660 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg658 = (1'h0);
  reg [(4'hc):(1'h0)] forvar656 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar655 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg654 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg265 = (1'h0);
  reg [(5'h12):(1'h0)] forvar263 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg260 = (1'h0);
  reg [(3'h4):(1'h0)] reg259 = (1'h0);
  reg [(3'h5):(1'h0)] reg257 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar256 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar255 = (1'h0);
  reg [(5'h17):(1'h0)] reg254 = (1'h0);
  reg [(4'h9):(1'h0)] reg252 = (1'h0);
  reg [(4'ha):(1'h0)] reg251 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg250 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar249 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg247 = (1'h0);
  reg [(4'h9):(1'h0)] reg246 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg244 = (1'h0);
  reg [(3'h5):(1'h0)] reg243 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg239 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg238 = (1'h0);
  reg [(5'h16):(1'h0)] forvar237 = (1'h0);
  reg [(4'hf):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg233 = (1'h0);
  reg [(5'h14):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg230 = (1'h0);
  reg [(2'h2):(1'h0)] reg228 = (1'h0);
  reg [(5'h14):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg225 = (1'h0);
  reg [(2'h2):(1'h0)] forvar224 = (1'h0);
  reg [(5'h18):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg219 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg125 = (1'h0);
  reg [(5'h17):(1'h0)] forvar121 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg120 = (1'h0);
  reg [(5'h14):(1'h0)] reg119 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar118 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg115 = (1'h0);
  reg [(5'h15):(1'h0)] reg114 = (1'h0);
  reg [(4'hf):(1'h0)] reg111 = (1'h0);
  reg [(4'he):(1'h0)] reg108 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg105 = (1'h0);
  reg [(4'h9):(1'h0)] reg104 = (1'h0);
  reg [(5'h14):(1'h0)] reg100 = (1'h0);
  reg [(4'hf):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar100 = (1'h0);
  reg [(5'h11):(1'h0)] reg99 = (1'h0);
  reg [(2'h2):(1'h0)] reg97 = (1'h0);
  reg [(5'h17):(1'h0)] reg94 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg93 = (1'h0);
  reg [(5'h10):(1'h0)] reg92 = (1'h0);
  assign y = {wire818,
                 wire745,
                 wire703,
                 wire702,
                 wire662,
                 wire651,
                 wire649,
                 wire434,
                 wire433,
                 wire112,
                 wire124,
                 wire216,
                 wire431,
                 reg807,
                 reg817,
                 reg816,
                 reg812,
                 reg809,
                 reg806,
                 reg803,
                 reg800,
                 reg799,
                 reg798,
                 reg795,
                 reg791,
                 reg788,
                 reg786,
                 reg781,
                 reg780,
                 reg779,
                 reg776,
                 reg773,
                 reg772,
                 reg770,
                 reg767,
                 reg766,
                 reg761,
                 reg759,
                 reg758,
                 reg750,
                 reg749,
                 reg744,
                 reg742,
                 reg740,
                 reg739,
                 reg734,
                 reg733,
                 reg732,
                 reg730,
                 reg729,
                 reg724,
                 reg722,
                 reg721,
                 reg720,
                 reg704,
                 reg716,
                 reg713,
                 reg712,
                 reg711,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 reg705,
                 reg700,
                 reg699,
                 reg698,
                 reg696,
                 reg695,
                 reg694,
                 reg689,
                 reg687,
                 reg686,
                 reg684,
                 reg683,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg675,
                 reg674,
                 reg671,
                 reg669,
                 reg667,
                 reg664,
                 reg661,
                 reg659,
                 reg657,
                 reg653,
                 reg652,
                 reg126,
                 reg123,
                 reg122,
                 reg117,
                 reg116,
                 reg113,
                 reg110,
                 reg109,
                 reg103,
                 reg101,
                 reg98,
                 reg96,
                 reg95,
                 reg218,
                 reg221,
                 reg226,
                 reg229,
                 reg224,
                 reg232,
                 reg234,
                 reg236,
                 reg240,
                 reg241,
                 reg245,
                 reg248,
                 reg253,
                 reg258,
                 reg261,
                 reg262,
                 reg264,
                 reg815,
                 reg814,
                 forvar813,
                 reg811,
                 reg810,
                 reg808,
                 forvar807,
                 forvar805,
                 reg804,
                 reg802,
                 reg801,
                 reg797,
                 forvar796,
                 reg794,
                 reg793,
                 reg792,
                 forvar790,
                 forvar789,
                 reg787,
                 reg785,
                 forvar784,
                 forvar783,
                 reg782,
                 reg778,
                 reg777,
                 forvar775,
                 reg774,
                 reg771,
                 reg769,
                 reg768,
                 reg765,
                 reg764,
                 reg763,
                 reg762,
                 forvar760,
                 reg757,
                 forvar756,
                 reg755,
                 forvar754,
                 reg753,
                 reg752,
                 reg751,
                 reg748,
                 forvar747,
                 forvar746,
                 reg743,
                 forvar741,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 reg731,
                 forvar729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg723,
                 reg719,
                 reg718,
                 reg717,
                 reg715,
                 reg714,
                 reg706,
                 forvar704,
                 forvar686,
                 reg701,
                 reg697,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg688,
                 reg685,
                 reg682,
                 forvar681,
                 reg676,
                 reg673,
                 reg672,
                 forvar670,
                 forvar668,
                 reg666,
                 forvar665,
                 reg663,
                 reg660,
                 reg658,
                 forvar656,
                 forvar655,
                 reg654,
                 reg265,
                 forvar263,
                 reg260,
                 reg259,
                 reg257,
                 forvar256,
                 forvar255,
                 reg254,
                 reg252,
                 reg251,
                 reg250,
                 forvar249,
                 reg247,
                 reg246,
                 reg237,
                 reg244,
                 reg243,
                 reg242,
                 reg239,
                 reg238,
                 forvar237,
                 reg235,
                 reg233,
                 reg231,
                 reg230,
                 reg228,
                 reg227,
                 reg225,
                 forvar224,
                 reg223,
                 reg222,
                 reg220,
                 reg219,
                 reg125,
                 forvar121,
                 reg120,
                 reg119,
                 forvar118,
                 reg115,
                 reg114,
                 reg111,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg100,
                 reg102,
                 forvar100,
                 reg99,
                 reg97,
                 reg94,
                 reg93,
                 reg92,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire89)
        begin
          reg92 = $signed(wire90[(1'h0):(1'h0)]);
        end
      else
        begin
          if (({wire88[(2'h2):(2'h2)]} ?
              ((wire91 != wire91[(3'h6):(1'h0)]) * {$unsigned((wire89 > (8'hb7)))}) : $unsigned(wire89)))
            begin
              reg92 = (8'hac);
              reg93 = $unsigned(wire88[(2'h3):(1'h0)]);
              reg94 = wire90;
              reg95 <= $signed((!(({reg94, (8'h9c)} ?
                      wire91[(1'h1):(1'h1)] : $signed(wire91)) ?
                  wire88 : reg92[(4'hc):(3'h4)])));
              reg96 <= (wire90 >>> (($unsigned(wire90) <<< wire91) ?
                  ((wire91[(3'h4):(2'h2)] - ((8'h9d) >> reg92)) ?
                      $unsigned(reg95[(5'h14):(2'h3)]) : (wire88 != (8'hbf))) : reg92));
            end
          else
            begin
              reg92 = reg95[(1'h0):(1'h0)];
              reg95 <= $signed((^~($signed($signed(reg96)) + wire88[(3'h7):(1'h1)])));
              reg96 <= (-{((reg95 ?
                      $unsigned(wire90) : $unsigned(reg92)) == (^$unsigned(reg93))),
                  $unsigned($unsigned((reg96 | wire91)))});
              reg97 = $signed($unsigned({((^reg92) >> $unsigned(wire90))}));
              reg98 <= {$unsigned(((7'h48) ? reg94 : ({wire90} ^ wire90))),
                  ($unsigned($signed($unsigned(wire91))) * wire89)};
            end
        end
      reg99 = (^(wire88[(2'h2):(1'h1)] <<< {(7'h47)}));
      if (({$unsigned(reg97[(1'h0):(1'h0)])} ? wire88[(2'h2):(2'h2)] : (7'h48)))
        begin
          for (forvar100 = (1'h0); (forvar100 < (1'h0)); forvar100 = (forvar100 + (1'h1)))
            begin
              reg101 <= {($signed((~(!wire90))) <<< ($unsigned($unsigned(wire91)) == $unsigned((reg94 ?
                      wire88 : reg97)))),
                  reg94};
              reg102 = $unsigned($signed((wire91[(4'h8):(3'h5)] ^~ wire91)));
            end
          reg103 <= (((({reg94,
              (7'h46)} << ((8'hb8) == reg94)) <<< wire88[(3'h5):(2'h2)]) ^ wire91) ^~ {$unsigned($unsigned(reg101[(4'he):(4'he)]))});
        end
      else
        begin
          reg100 = {wire89};
          reg102 = $signed($unsigned((((reg93 ? forvar100 : reg98) ?
              {forvar100} : $unsigned(reg94)) && {{wire91}})));
          reg104 = (~^wire88);
          reg105 = reg98;
          if ({$signed(wire89[(1'h0):(1'h0)])})
            begin
              reg106 = ($unsigned({(7'h4a), (~^$unsigned(wire89))}) ?
                  (wire91 << ($unsigned($unsigned(reg97)) >> (^(~^reg99)))) : {{(^$unsigned(reg102)),
                          reg95},
                      ((reg103 ? (~|reg92) : (reg99 || reg104)) ?
                          ($signed((8'ha7)) ?
                              (reg95 ?
                                  (7'h46) : reg105) : reg95) : ($unsigned(reg100) ?
                              reg92 : $unsigned(reg103)))});
              reg107 = ($unsigned((-{{reg97},
                  $signed(forvar100)})) * $signed($unsigned(reg100)));
              reg108 = $unsigned(((($unsigned(reg99) ?
                          (&forvar100) : $signed(reg97)) ?
                      reg106[(5'h13):(3'h6)] : $unsigned((wire89 ?
                          wire89 : reg92))) ?
                  {$signed(((8'hbe) ? reg105 : reg101)),
                      reg98} : reg99[(5'h11):(3'h7)]));
              reg109 <= ($signed($unsigned($unsigned((reg96 ?
                  forvar100 : (8'ha9))))) << {reg97[(1'h0):(1'h0)],
                  reg104[(3'h5):(2'h3)]});
              reg110 <= $signed(wire89);
            end
          else
            begin
              reg106 = (^$signed(($unsigned(wire89) > reg95[(5'h17):(3'h7)])));
              reg109 <= wire91[(4'hc):(4'hc)];
              reg111 = $signed(($unsigned($signed(((7'h4a) ?
                      forvar100 : (8'hbf)))) ?
                  $unsigned({reg105[(4'h9):(3'h4)]}) : $unsigned(($signed(reg102) | {reg107}))));
            end
        end
    end
  assign wire112 = {{({(8'h9d)} ? reg103[(3'h7):(2'h3)] : $signed(reg109)),
                           (((&wire91) == $unsigned((7'h44))) ?
                               ((~|(7'h40)) ?
                                   {wire89} : reg109[(5'h12):(4'hc)]) : $signed((reg110 < reg95)))}};
  always
    @(posedge clk) begin
      reg113 <= wire90;
      reg114 = (~&(reg96[(1'h1):(1'h0)] < (!(7'h47))));
      reg115 = reg101;
      reg116 <= wire88[(3'h7):(3'h6)];
      reg117 <= (reg113 ?
          (!(&($signed(reg110) > ((8'hb3) >> reg115)))) : {(wire90 ~^ reg103[(3'h7):(3'h4)]),
              wire89[(2'h2):(1'h1)]});
    end
  always
    @(posedge clk) begin
      for (forvar118 = (1'h0); (forvar118 < (2'h3)); forvar118 = (forvar118 + (1'h1)))
        begin
          reg119 = (7'h48);
          reg120 = ((^(|{{wire88, reg109}, (!(7'h4a))})) >> $unsigned(reg101));
        end
      for (forvar121 = (1'h0); (forvar121 < (3'h4)); forvar121 = (forvar121 + (1'h1)))
        begin
          reg122 <= {forvar121[(4'hd):(4'hd)]};
        end
      reg123 <= forvar121;
    end
  assign wire124 = reg116[(3'h6):(2'h2)];
  always
    @(posedge clk) begin
      reg125 = $unsigned(({reg116[(1'h1):(1'h0)], $unsigned($signed(wire88))} ?
          reg113[(5'h14):(4'ha)] : (($unsigned(reg113) ?
                  {wire112, (8'ha9)} : wire88[(1'h1):(1'h1)]) ?
              {(reg101 ? reg103 : (8'h9e))} : reg103[(4'h9):(3'h5)])));
      reg126 <= (~reg117);
    end
  module127 #() modinst217 (.wire130(reg123), .wire131(wire112), .wire129(reg122), .wire132(wire88), .wire128(reg113), .y(wire216), .clk(clk));
  always
    @(posedge clk) begin
      reg218 <= (~reg110);
      if ($signed($unsigned($unsigned(wire90))))
        begin
          if ((~&{((~reg123) + $unsigned((wire124 ? (8'ha9) : wire112))),
              $unsigned($unsigned(reg113[(2'h2):(1'h1)]))}))
            begin
              reg219 = (!(~reg95));
              reg220 = (|reg103);
            end
          else
            begin
              reg221 <= ($unsigned((reg95 + $signed((wire91 ?
                      wire216 : (7'h47))))) ?
                  reg110[(5'h17):(5'h13)] : wire90);
              reg222 = $unsigned($unsigned(((~reg98[(1'h1):(1'h0)]) & {$signed(reg123)})));
            end
          reg223 = $unsigned(((7'h45) ?
              $unsigned($unsigned(reg117[(3'h4):(2'h3)])) : $signed({$unsigned(wire88)})));
          for (forvar224 = (1'h0); (forvar224 < (3'h4)); forvar224 = (forvar224 + (1'h1)))
            begin
              reg225 = reg222;
              reg226 <= ((7'h44) ^~ (reg103 ?
                  ($unsigned((reg126 ?
                      reg126 : reg117)) + wire91[(4'hc):(4'h9)]) : reg101));
              reg227 = ($unsigned($signed($unsigned($signed(reg116)))) + (((^$signed(reg223)) ?
                  reg221 : ($unsigned(reg109) ?
                      (^~wire89) : (wire112 ?
                          wire90 : reg126))) == $unsigned(wire89[(2'h2):(1'h0)])));
              reg228 = reg227;
              reg229 <= reg225[(3'h7):(3'h7)];
            end
        end
      else
        begin
          if (reg229[(5'h10):(4'h8)])
            begin
              reg221 <= $unsigned((+(((reg103 != reg117) ?
                  (+reg222) : $signed(wire112)) ~^ $signed((8'hbd)))));
            end
          else
            begin
              reg221 <= reg221;
              reg224 <= ((({forvar224} >> (reg225[(4'hc):(4'h9)] << (^~reg116))) ?
                      $unsigned($unsigned($unsigned(reg223))) : reg113[(5'h12):(4'ha)]) ?
                  (&$signed($signed($signed(reg229)))) : {reg109[(4'he):(4'h9)]});
              reg226 <= forvar224[(2'h2):(2'h2)];
            end
          if ((~^$signed($signed(((^~reg227) ?
              {reg225, wire89} : $unsigned(reg116))))))
            begin
              reg227 = $unsigned({(~(+(wire216 >= (7'h49)))),
                  (reg221[(1'h0):(1'h0)] >>> ($unsigned(wire112) ~^ {reg103}))});
              reg229 <= ($unsigned((|reg226)) ? (8'hb4) : (8'hb3));
              reg230 = (($unsigned((~((8'hae) >= reg228))) ^ $signed((~&(reg116 ?
                      reg109 : reg98)))) ?
                  wire88[(2'h3):(1'h0)] : (($unsigned((reg227 || wire91)) ?
                      reg113[(4'h8):(1'h0)] : ((~&wire88) > (reg101 <= reg95))) == {((reg109 >> reg220) ?
                          forvar224 : wire90),
                      {reg218[(2'h2):(2'h2)], reg96}}));
            end
          else
            begin
              reg227 = $unsigned((wire124[(2'h2):(1'h1)] ?
                  {{$signed(reg218),
                          reg117[(5'h10):(2'h2)]}} : (~|$signed($signed(reg228)))));
            end
          reg231 = ((reg113[(4'he):(4'he)] || $unsigned(reg95)) ^~ {{(~|reg226),
                  wire124[(1'h1):(1'h1)]},
              reg221});
          if ({(reg117[(4'hb):(4'hb)] ^~ (|$unsigned($signed(reg117)))),
              reg221})
            begin
              reg232 <= $signed(($signed(($signed(wire89) >>> {reg101})) ?
                  (+reg230[(4'hd):(4'hb)]) : (wire88[(3'h6):(3'h4)] ?
                      wire88[(1'h0):(1'h0)] : ({reg230, reg95} ?
                          ((7'h44) ^~ (8'hba)) : reg229[(4'h8):(1'h1)]))));
              reg233 = ($unsigned($unsigned($unsigned(reg116[(3'h5):(1'h1)]))) || (((reg96 ?
                      (reg123 >= wire88) : {reg113}) + reg225) ?
                  $unsigned($unsigned((reg110 ?
                      reg123 : reg116))) : {($unsigned((7'h41)) ?
                          $unsigned(reg95) : $signed(reg122))}));
              reg234 <= {{$unsigned($signed(reg226))},
                  $signed((~|wire124[(2'h2):(1'h0)]))};
              reg235 = $unsigned((reg227 ?
                  $signed(((~&reg223) ?
                      reg226 : $unsigned(reg221))) : (|reg231)));
            end
          else
            begin
              reg233 = (|reg232);
              reg235 = {$signed((reg222[(2'h2):(1'h0)] >>> reg226))};
              reg236 <= ($signed($unsigned(reg109)) ?
                  (^wire216) : reg219[(4'hd):(1'h0)]);
            end
        end
      if ({(reg223[(4'hb):(4'h9)] ?
              (($signed(reg223) && ((8'hb3) ? reg117 : (7'h4a))) * {((8'hab) ?
                      reg227 : reg219),
                  {(8'hb5), (8'haa)}}) : ((|(8'hb5)) & wire216)),
          reg227})
        begin
          for (forvar237 = (1'h0); (forvar237 < (3'h4)); forvar237 = (forvar237 + (1'h1)))
            begin
              reg238 = ($unsigned(wire90) - reg117[(4'hc):(4'hc)]);
              reg239 = $unsigned((^($signed($unsigned((8'had))) & ($unsigned(reg123) ?
                  (~^reg234) : reg116[(1'h0):(1'h0)]))));
              reg240 <= wire91;
              reg241 <= $unsigned({(!$signed($unsigned(wire91))),
                  (~|$signed($signed(forvar237)))});
            end
          reg242 = (((-$signed((~|reg96))) > wire88) ?
              ((reg225 ? (+{reg98}) : ((&wire89) & $signed(reg241))) ?
                  reg103 : (reg116[(4'h8):(3'h4)] ?
                      (!((8'hb6) - (7'h41))) : ((reg236 ?
                          reg233 : reg241) ~^ $signed((8'ha1))))) : $unsigned(reg240));
          reg243 = reg109[(1'h1):(1'h0)];
          reg244 = wire89[(1'h1):(1'h1)];
        end
      else
        begin
          if ($signed(({(+$signed(reg103))} >= reg126)))
            begin
              reg237 = $signed((wire91[(2'h2):(1'h0)] << (((reg113 ?
                  reg244 : (8'hbe)) + reg101[(4'hb):(2'h3)]) >= reg231)));
              reg240 <= $unsigned($unsigned((~&$unsigned($signed(wire124)))));
              reg242 = (($signed(reg244) <= (~|$unsigned($unsigned((7'h40))))) ?
                  (+$unsigned((wire124 ?
                      (reg231 | (7'h49)) : $signed(reg231)))) : ($unsigned(((-reg227) ?
                          reg219 : $signed(reg110))) ?
                      reg122[(3'h7):(1'h1)] : reg98));
              reg245 <= (^(wire216[(3'h5):(1'h0)] ?
                  reg226[(4'h8):(3'h4)] : reg242));
            end
          else
            begin
              reg240 <= $unsigned($unsigned(($unsigned((~^reg110)) ?
                  reg122[(3'h4):(3'h4)] : ((reg223 ?
                      wire91 : reg95) - reg231))));
            end
          reg246 = {reg229};
        end
      if (reg220)
        begin
          reg247 = $unsigned(reg101[(4'he):(1'h0)]);
        end
      else
        begin
          reg248 <= forvar224[(1'h0):(1'h0)];
          for (forvar249 = (1'h0); (forvar249 < (3'h4)); forvar249 = (forvar249 + (1'h1)))
            begin
              reg250 = reg240;
            end
          if ((|(reg126 ? reg248 : (+$unsigned($unsigned((8'haf)))))))
            begin
              reg251 = $unsigned(((8'h9c) <= $unsigned(($unsigned(reg235) ?
                  $unsigned(wire89) : $unsigned(reg117)))));
              reg252 = {(reg220 ?
                      reg113[(5'h13):(5'h13)] : reg239[(4'ha):(1'h1)])};
            end
          else
            begin
              reg253 <= reg226;
            end
        end
    end
  always
    @(posedge clk) begin
      reg254 = $signed(((((reg234 == reg248) << {(8'h9f)}) <<< wire216[(4'h9):(3'h6)]) || $signed({reg232,
          $signed(reg98)})));
      for (forvar255 = (1'h0); (forvar255 < (2'h3)); forvar255 = (forvar255 + (1'h1)))
        begin
          for (forvar256 = (1'h0); (forvar256 < (3'h4)); forvar256 = (forvar256 + (1'h1)))
            begin
              reg257 = (|((8'hac) || reg95[(4'hb):(3'h5)]));
            end
          reg258 <= (^$unsigned($signed($signed((~^(8'hbd))))));
          if (reg254[(3'h4):(1'h0)])
            begin
              reg259 = (($signed(reg101[(3'h5):(3'h4)]) * ((~|(8'hbc)) ?
                      $signed((^reg101)) : forvar256)) ?
                  (~|$signed(reg245)) : {$unsigned($signed(((8'hb6) ?
                          reg122 : reg103))),
                      $signed((&(^reg113)))});
            end
          else
            begin
              reg259 = ($unsigned((((reg110 && reg221) * (reg126 ?
                      reg117 : wire90)) ?
                  reg101[(3'h4):(2'h2)] : wire124)) * (wire91 ?
                  ((forvar255 ?
                      (+reg259) : $signed(reg254)) || $unsigned((reg117 ?
                      forvar256 : reg253))) : reg240));
              reg260 = $unsigned(reg218);
              reg261 <= (+$signed(({(reg221 ? reg96 : reg259),
                      $unsigned(reg123)} ?
                  ((+(8'hb4)) ?
                      (+wire90) : (-wire88)) : ({(8'hb1)} * (wire216 << wire89)))));
            end
          reg262 <= {reg261[(1'h0):(1'h0)]};
          for (forvar263 = (1'h0); (forvar263 < (1'h1)); forvar263 = (forvar263 + (1'h1)))
            begin
              reg264 <= reg257[(2'h2):(1'h0)];
            end
        end
      reg265 = reg103;
    end
  module266 #() modinst432 (.wire267(wire112), .wire269(reg113), .wire271(reg234), .wire270(reg116), .clk(clk), .y(wire431), .wire268(reg101));
  assign wire433 = reg98[(3'h5):(3'h5)];
  assign wire434 = (|$unsigned($signed($unsigned((reg240 ?
                       reg221 : wire431)))));
  module435 #() modinst650 (.wire438(reg262), .wire436(reg110), .clk(clk), .wire439(reg241), .wire437(reg229), .y(wire649), .wire440(reg113));
  assign wire651 = $signed($signed($signed(reg122)));
  always
    @(posedge clk) begin
      reg652 <= wire88;
      reg653 <= reg248;
      reg654 = $unsigned(($signed((+reg652[(2'h2):(1'h1)])) > ($signed(reg240) ?
          $signed(reg110) : ($signed(reg116) ?
              (reg126 ? (8'ha9) : reg241) : (wire649 ? reg652 : wire112)))));
    end
  always
    @(posedge clk) begin
      for (forvar655 = (1'h0); (forvar655 < (3'h4)); forvar655 = (forvar655 + (1'h1)))
        begin
          for (forvar656 = (1'h0); (forvar656 < (1'h1)); forvar656 = (forvar656 + (1'h1)))
            begin
              reg657 <= wire90;
              reg658 = ($signed((((^reg232) || reg258[(3'h7):(3'h4)]) & (7'h49))) ?
                  wire216[(3'h7):(1'h0)] : (8'hb6));
              reg659 <= $unsigned((reg248 >= reg122));
              reg660 = (reg96[(1'h1):(1'h1)] ~^ $unsigned(reg113[(1'h1):(1'h1)]));
              reg661 <= reg226[(2'h3):(1'h0)];
            end
        end
    end
  assign wire662 = {$unsigned(reg224),
                       {((!wire434[(4'ha):(3'h7)]) ?
                               (~&$unsigned(wire88)) : $signed({reg221,
                                   reg657}))}};
  always
    @(posedge clk) begin
      if (reg229)
        begin
          reg663 = $unsigned(({reg258[(4'h9):(3'h5)], reg253[(2'h2):(1'h1)]} ?
              $unsigned((~^$signed(reg258))) : (!$unsigned(reg262[(5'h16):(3'h6)]))));
          reg664 <= ({wire89[(2'h2):(1'h0)], $unsigned(wire216)} ?
              reg661[(3'h6):(2'h2)] : reg248);
        end
      else
        begin
          reg664 <= reg264[(2'h2):(2'h2)];
          for (forvar665 = (1'h0); (forvar665 < (3'h4)); forvar665 = (forvar665 + (1'h1)))
            begin
              reg666 = $signed({reg122, reg110});
              reg667 <= (~&wire431);
            end
        end
      for (forvar668 = (1'h0); (forvar668 < (1'h1)); forvar668 = (forvar668 + (1'h1)))
        begin
          reg669 <= (8'hb3);
          for (forvar670 = (1'h0); (forvar670 < (1'h0)); forvar670 = (forvar670 + (1'h1)))
            begin
              reg671 <= {(~|$signed($signed((+reg98))))};
              reg672 = $signed(((($signed(reg666) == $unsigned(reg98)) >= $signed($unsigned((8'hbd)))) && wire649[(3'h7):(2'h2)]));
              reg673 = $unsigned((^~$signed($unsigned((reg262 ?
                  reg240 : reg96)))));
            end
          reg674 <= wire124;
          reg675 <= ((reg663[(4'hb):(1'h1)] || (8'hbb)) ?
              (|$unsigned(($signed(reg258) ~^ {reg98}))) : reg109[(3'h4):(2'h3)]);
          if ($unsigned((reg240[(1'h1):(1'h0)] ~^ (~(~^(reg226 ?
              reg673 : reg653))))))
            begin
              reg676 = reg666;
              reg677 <= (&($signed(({reg95} ~^ reg116[(4'hf):(3'h7)])) ?
                  $unsigned($unsigned({reg98, wire112})) : reg663));
              reg678 <= ($signed((^~$unsigned(reg253))) ?
                  $signed({$signed($signed((7'h45)))}) : (&$unsigned((8'ha1))));
              reg679 <= (wire434 >>> $signed(($unsigned((reg664 ?
                      wire651 : reg657)) ?
                  $unsigned($signed(reg241)) : $signed($unsigned(wire88)))));
              reg680 <= reg672;
            end
          else
            begin
              reg677 <= reg113;
              reg678 <= ($signed((&(~^reg113[(4'hb):(3'h5)]))) >= $unsigned($signed(reg110[(3'h6):(1'h0)])));
            end
        end
      for (forvar681 = (1'h0); (forvar681 < (2'h2)); forvar681 = (forvar681 + (1'h1)))
        begin
          reg682 = ($unsigned((($signed(reg226) ?
                  $unsigned(reg664) : wire649) >>> ($unsigned(reg659) ?
                  ((8'hac) ? reg659 : wire90) : reg669[(4'h8):(2'h2)]))) ?
              ((+{(&(8'ha4)), reg98[(4'hb):(3'h4)]}) ?
                  ({(reg675 ? reg261 : reg663), reg103[(4'h9):(2'h2)]} ?
                      (((8'ha4) >> reg123) ?
                          $signed(wire434) : ((8'hbd) ~^ reg258)) : reg113) : reg661[(4'hc):(2'h2)]) : (&$signed($unsigned({(8'hab)}))));
          reg683 <= (~&((8'hbb) ?
              $unsigned(reg221) : $signed(($unsigned(reg226) | reg675[(3'h6):(3'h4)]))));
        end
      if (wire89[(1'h0):(1'h0)])
        begin
          if (($unsigned(reg663) ? reg98 : reg659[(4'hd):(1'h0)]))
            begin
              reg684 <= $unsigned((reg236[(3'h6):(3'h5)] > (~$unsigned($signed(reg675)))));
              reg685 = ($unsigned(reg652[(3'h5):(3'h5)]) ?
                  (8'ha7) : {$signed(((reg661 ? wire651 : reg123) - reg679)),
                      (!((8'hba) >> reg218))});
            end
          else
            begin
              reg685 = (~^($unsigned(wire91) ?
                  $unsigned((reg95[(5'h15):(4'ha)] ^~ (8'ha4))) : reg669[(5'h15):(1'h1)]));
              reg686 <= wire91;
              reg687 <= $unsigned({reg113,
                  ({$unsigned(reg229), reg232[(5'h14):(4'hf)]} ?
                      reg678[(3'h7):(3'h6)] : ($unsigned(reg678) || reg669[(2'h2):(2'h2)]))});
              reg688 = wire216;
            end
          if (reg262[(5'h10):(5'h10)])
            begin
              reg689 <= reg653[(2'h3):(2'h3)];
              reg690 = reg671;
            end
          else
            begin
              reg690 = (|reg683[(1'h1):(1'h1)]);
              reg691 = {($signed((~&reg676)) | ((~^(~^reg117)) && (reg678 ?
                      (8'hbe) : $signed(reg678))))};
              reg692 = (($signed(({reg123} ?
                  (^~reg253) : (forvar665 - reg101))) - (8'haf)) & (^~$signed((wire90[(3'h4):(3'h4)] ?
                  $unsigned(forvar665) : reg682[(5'h14):(4'ha)]))));
              reg693 = (($unsigned((|(-reg678))) == reg95) ?
                  reg676[(4'hb):(1'h0)] : $signed(({$unsigned(forvar681),
                          {reg240, reg669}} ?
                      (^~(reg659 >= reg659)) : (reg113 ?
                          $unsigned(forvar670) : {(7'h44), wire90}))));
              reg694 <= $signed($signed(reg671));
            end
          reg695 <= (reg688 ?
              $unsigned(reg95) : $unsigned($signed({$signed(reg248),
                  {reg677}})));
          if ((~^((reg675[(1'h1):(1'h0)] ?
              ((~^reg675) ~^ {reg667}) : ((|reg667) ?
                  ((8'hab) - (8'hb2)) : (~&reg123))) ^~ (reg262[(1'h1):(1'h0)] + reg691[(3'h6):(2'h2)]))))
            begin
              reg696 <= (~|(~{reg673, $unsigned(reg679)}));
              reg697 = ($unsigned(((reg113[(4'hb):(4'ha)] < (reg241 ?
                      reg686 : reg240)) ?
                  $signed(reg122[(2'h2):(1'h0)]) : wire433[(2'h2):(1'h1)])) > ((~&($unsigned(reg262) ?
                      reg669 : reg113[(5'h17):(3'h5)])) ?
                  (reg677[(4'hb):(4'hb)] ?
                      reg253[(2'h3):(2'h2)] : (reg657 - (reg666 ?
                          reg262 : wire433))) : (~|$signed($signed(reg694)))));
              reg698 <= reg116;
              reg699 <= (~|(^~reg221));
              reg700 <= {reg110[(2'h3):(1'h1)], reg677[(2'h3):(2'h3)]};
            end
          else
            begin
              reg696 <= $unsigned($signed($signed($unsigned($unsigned(reg659)))));
            end
          reg701 = (((8'h9f) ?
                  ($unsigned((reg672 != reg699)) * $unsigned($unsigned(wire124))) : ($signed((~reg116)) <= reg117)) ?
              (~$signed({(!reg673), $unsigned((8'ha4))})) : (!reg699));
        end
      else
        begin
          if (reg693[(4'h9):(4'h9)])
            begin
              reg684 <= {wire431, (~&reg680[(4'h9):(3'h5)])};
            end
          else
            begin
              reg684 <= {{($unsigned(reg234[(1'h0):(1'h0)]) ?
                          $signed((wire662 || reg673)) : $signed((^reg693))),
                      $unsigned($unsigned(reg678))},
                  reg676[(3'h7):(3'h6)]};
              reg685 = ({$signed($unsigned(reg224)),
                  (&$unsigned((^~wire89)))} != $signed((&{reg261,
                  reg241[(1'h1):(1'h1)]})));
            end
          for (forvar686 = (1'h0); (forvar686 < (1'h0)); forvar686 = (forvar686 + (1'h1)))
            begin
              reg688 = $unsigned($unsigned((reg694 & {(reg693 < reg98)})));
              reg689 <= reg96;
            end
          reg694 <= $signed(reg678);
        end
    end
  assign wire702 = reg218[(3'h4):(3'h4)];
  assign wire703 = (8'hbc);
  always
    @(posedge clk) begin
      if ($unsigned((((+reg101) ? reg95 : $unsigned($unsigned((8'h9d)))) ?
          (^~wire703) : $signed((~|reg699)))))
        begin
          for (forvar704 = (1'h0); (forvar704 < (2'h3)); forvar704 = (forvar704 + (1'h1)))
            begin
              reg705 <= reg262;
              reg706 = wire433[(2'h2):(2'h2)];
              reg707 <= wire703[(2'h2):(2'h2)];
              reg708 <= ((reg674[(5'h13):(3'h4)] || $signed(reg677)) ?
                  $signed($signed($signed(wire112[(1'h1):(1'h1)]))) : (reg674[(4'he):(4'ha)] ?
                      ($signed((^wire433)) & wire702[(4'hb):(4'ha)]) : reg674));
              reg709 <= (((+wire91[(4'hc):(3'h4)]) ?
                  reg240[(4'ha):(4'ha)] : (8'ha4)) != {{(~$signed(reg262)),
                      (^~((8'hb1) ? wire703 : reg689))}});
            end
          if ((-(7'h40)))
            begin
              reg710 <= reg264[(3'h5):(3'h4)];
              reg711 <= (&$unsigned({reg126[(3'h4):(2'h3)], reg680}));
              reg712 <= reg661[(4'h9):(2'h3)];
              reg713 <= $unsigned((^~$unsigned(reg229)));
              reg714 = {$unsigned($signed(reg262[(3'h4):(2'h3)]))};
            end
          else
            begin
              reg714 = {((reg686[(4'ha):(2'h3)] == ((!wire702) ?
                      $signed((8'haf)) : (reg709 & reg126))) << $signed($unsigned({reg657})))};
              reg715 = $unsigned($signed((7'h45)));
              reg716 <= (|$unsigned((~((reg264 << reg674) == (reg116 ?
                  reg101 : reg689)))));
              reg717 = reg218[(2'h2):(2'h2)];
              reg718 = (((+reg712[(2'h3):(1'h1)]) | $signed((reg715[(2'h2):(1'h0)] << reg686))) ?
                  $unsigned(reg652) : (($signed((+reg126)) <<< $unsigned(reg245[(5'h12):(3'h7)])) <<< $signed(((&reg674) ?
                      $unsigned(reg659) : $unsigned(reg700)))));
            end
          reg719 = reg657;
        end
      else
        begin
          if (reg705)
            begin
              reg704 <= (~&({reg98[(2'h3):(1'h0)]} ?
                  (((~|reg218) ?
                          $signed(wire431) : (reg116 ? (8'ha5) : reg109)) ?
                      reg674 : {reg229}) : $unsigned($signed(wire88[(1'h0):(1'h0)]))));
              reg706 = $unsigned(reg704);
              reg707 <= (8'hb7);
              reg714 = {{$signed((7'h44)), reg126},
                  $signed(((-$signed(wire112)) ?
                      ({reg96,
                          reg680} >= (7'h41)) : (&reg229[(3'h4):(1'h1)])))};
            end
          else
            begin
              reg706 = $unsigned((+reg248));
              reg714 = (|(7'h49));
              reg716 <= reg229;
              reg720 <= wire703[(3'h5):(3'h4)];
              reg721 <= ($signed(wire91) >> reg261);
            end
          reg722 <= (~^((($signed((8'hb7)) - reg671[(4'h9):(3'h4)]) ?
                  ((reg713 ?
                      reg704 : reg696) >> reg122[(2'h3):(2'h2)]) : ($signed((7'h43)) ?
                      reg101[(3'h4):(2'h3)] : {wire88, reg687})) ?
              ({(reg711 != forvar704), {(7'h40)}} ?
                  (^~$signed(reg126)) : $unsigned($signed(wire433))) : reg661[(4'h8):(1'h0)]));
          if (reg700[(2'h2):(1'h0)])
            begin
              reg723 = (8'hb7);
              reg724 <= reg674;
              reg725 = wire112;
              reg726 = $signed((&reg714));
            end
          else
            begin
              reg723 = ({reg721} > (+$signed({$unsigned(reg261), (&wire651)})));
              reg724 <= ({reg720, ({reg261} << {reg234})} ?
                  (reg113[(4'ha):(2'h3)] && ((!(reg116 ? wire216 : reg96)) ?
                      {(wire703 - (8'ha2)), reg677} : {{reg258}})) : (reg710 ?
                      reg241[(4'hd):(3'h7)] : (^(^reg653))));
              reg725 = {$unsigned($unsigned(({reg123,
                      reg705} | reg680[(1'h0):(1'h0)])))};
              reg726 = ($unsigned((($signed(reg687) - (+reg714)) ^ (|$unsigned(wire651)))) ~^ $signed((-(reg262[(5'h15):(4'he)] <<< wire90[(2'h2):(1'h0)]))));
              reg727 = ((-({(reg717 ~^ reg723),
                      (&reg98)} >>> $unsigned($unsigned(reg226)))) ?
                  wire90 : reg708);
            end
          reg728 = reg218[(1'h1):(1'h1)];
        end
      if ($unsigned((reg117[(5'h12):(4'hc)] - ($signed({(8'ha5),
          reg707}) || wire649))))
        begin
          reg729 <= (^(($signed($unsigned(reg718)) ^~ $unsigned((reg113 ?
              reg218 : reg708))) >> reg103[(4'hb):(3'h7)]));
        end
      else
        begin
          for (forvar729 = (1'h0); (forvar729 < (3'h4)); forvar729 = (forvar729 + (1'h1)))
            begin
              reg730 <= {reg221[(1'h0):(1'h0)]};
              reg731 = ((^~reg729) < wire89);
              reg732 <= (!$signed({(reg710 ? (~|reg667) : $signed(reg727)),
                  (&reg234)}));
              reg733 <= reg705[(4'hc):(1'h0)];
              reg734 <= (^~$unsigned((reg725[(2'h2):(2'h2)] ?
                  reg728 : (|reg709))));
            end
          if ($signed($signed(($unsigned($unsigned(reg123)) ^~ reg229[(1'h1):(1'h0)]))))
            begin
              reg735 = ($unsigned((({reg726} <= reg695[(3'h4):(2'h2)]) < (~(reg679 ?
                      reg680 : reg110)))) ?
                  (-(((^reg726) ~^ (reg234 ? reg734 : wire216)) + ({reg218} ?
                      (~^wire662) : (reg725 >>> reg699)))) : wire649);
              reg736 = (({wire702[(3'h5):(2'h3)],
                      (reg729 ? (reg686 == reg675) : reg704)} ~^ (((reg721 ?
                              reg696 : reg245) ?
                          (reg261 - reg236) : $unsigned(wire90)) ?
                      (reg262 ?
                          $signed(reg730) : reg707[(4'hd):(3'h7)]) : {(reg728 << reg229),
                          (reg735 ? reg726 : reg728)})) ?
                  $unsigned(reg234[(5'h12):(4'h8)]) : ((|$signed($unsigned(reg709))) ?
                      $signed((~|(|reg109))) : $signed($unsigned($signed(reg719)))));
              reg737 = (reg109[(4'hc):(4'ha)] ?
                  (^$signed($signed((wire431 >= (8'hb3))))) : $signed(reg669[(3'h5):(3'h4)]));
              reg738 = ($unsigned(((~&$unsigned((7'h42))) >>> $unsigned((^reg657)))) + ($unsigned($unsigned(reg677)) ?
                  reg721 : reg245));
              reg739 <= (|(!($signed(reg659) <= {{(8'h9e)},
                  (reg677 > (8'hb4))})));
            end
          else
            begin
              reg735 = reg736[(1'h1):(1'h0)];
              reg739 <= ($unsigned(wire433[(2'h2):(2'h2)]) ?
                  $signed($unsigned(wire89[(1'h1):(1'h1)])) : $signed((|((wire90 & reg721) >= (8'hb6)))));
              reg740 <= ($signed((+reg116)) ? reg671 : reg736[(2'h3):(2'h3)]);
            end
          for (forvar741 = (1'h0); (forvar741 < (3'h4)); forvar741 = (forvar741 + (1'h1)))
            begin
              reg742 <= reg95;
              reg743 = reg695;
            end
          reg744 <= (~|(~^$unsigned(reg117)));
        end
    end
  assign wire745 = reg258[(3'h7):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar746 = (1'h0); (forvar746 < (2'h3)); forvar746 = (forvar746 + (1'h1)))
        begin
          for (forvar747 = (1'h0); (forvar747 < (1'h1)); forvar747 = (forvar747 + (1'h1)))
            begin
              reg748 = reg117[(5'h11):(3'h5)];
              reg749 <= $unsigned($unsigned((($signed(wire702) ?
                  reg109 : (reg653 <= reg695)) || (~&(reg732 ?
                  reg667 : reg667)))));
              reg750 <= (~^reg699);
              reg751 = {reg262};
            end
          reg752 = reg675;
        end
      reg753 = ($signed(reg664[(2'h3):(2'h3)]) ?
          (($unsigned((reg258 > wire112)) <<< reg241) ?
              (-$signed((reg709 <<< reg117))) : $unsigned(((reg721 && reg229) | $unsigned((8'hbf))))) : (reg712[(3'h6):(3'h6)] ?
              ((&{reg671}) || ({reg248} ?
                  (reg710 < wire703) : ((8'h9c) - forvar746))) : (wire651[(4'ha):(4'h8)] | ((8'hb0) + (reg724 ?
                  reg733 : wire431)))));
      for (forvar754 = (1'h0); (forvar754 < (3'h4)); forvar754 = (forvar754 + (1'h1)))
        begin
          reg755 = ((($unsigned((~^reg700)) & $unsigned(reg711[(1'h1):(1'h0)])) <= ($unsigned((wire124 >> (8'h9e))) ?
              $unsigned({reg709}) : (|(reg749 || (7'h47))))) || ($unsigned((~&reg707[(4'h9):(2'h2)])) ?
              $unsigned((|$signed((8'ha4)))) : reg698));
          for (forvar756 = (1'h0); (forvar756 < (2'h3)); forvar756 = (forvar756 + (1'h1)))
            begin
              reg757 = reg751;
              reg758 <= reg675[(2'h3):(2'h2)];
            end
        end
      reg759 <= {wire431[(2'h2):(2'h2)],
          (reg742 ?
              (8'hb8) : ($unsigned($signed(reg694)) + $signed(reg264[(3'h4):(3'h4)])))};
      if ((reg122 ^~ (reg126 ? (-(8'hbb)) : $signed({(7'h47)}))))
        begin
          for (forvar760 = (1'h0); (forvar760 < (1'h1)); forvar760 = (forvar760 + (1'h1)))
            begin
              reg761 <= {($signed(((reg704 & reg229) + (reg721 ?
                      (8'hb2) : reg755))) == reg700[(2'h3):(2'h3)])};
              reg762 = $signed((+reg241));
              reg763 = {wire216[(1'h1):(1'h0)],
                  ($signed(reg696) ?
                      (^$signed(reg98[(3'h4):(2'h2)])) : reg749[(3'h5):(1'h0)])};
            end
          reg764 = ($signed((|((reg262 | reg744) < (reg677 ~^ reg716)))) ?
              reg704 : {(reg707[(3'h7):(3'h6)] - ((reg677 ?
                      (8'h9c) : reg680) <<< $unsigned(reg667)))});
          if (({($unsigned($unsigned(wire745)) ?
                  {(+reg748)} : (reg109 ^ $unsigned(reg716))),
              {$signed({reg680, reg763}),
                  ($signed(reg248) <<< {reg734,
                      reg221})}} == $signed($unsigned((|reg749[(1'h1):(1'h1)])))))
            begin
              reg765 = $signed($signed((reg755[(3'h5):(3'h4)] ?
                  (8'ha8) : wire90[(2'h2):(1'h1)])));
              reg766 <= reg669[(3'h6):(1'h1)];
            end
          else
            begin
              reg765 = forvar756;
              reg766 <= $signed((((reg687 ?
                      reg261[(1'h1):(1'h1)] : (!reg95)) == reg226[(4'ha):(4'h9)]) ?
                  reg687 : reg729[(3'h5):(2'h2)]));
              reg767 <= (($signed($signed(wire89)) | (~^reg232)) ?
                  (8'hbb) : reg765);
              reg768 = $unsigned({(($signed(forvar747) ?
                      $signed(reg759) : $unsigned(wire651)) <= reg710[(2'h2):(1'h1)]),
                  ((reg763[(3'h4):(1'h1)] << (^~reg744)) >> reg126[(4'h8):(4'h8)])});
            end
          reg769 = reg696;
          if (forvar756)
            begin
              reg770 <= $signed((($unsigned(reg659) || wire702[(1'h0):(1'h0)]) ?
                  $unsigned($signed((~reg755))) : ((reg700[(4'hc):(3'h5)] - reg757) ?
                      reg245[(3'h7):(1'h0)] : $unsigned((~^reg699)))));
              reg771 = ($signed(((reg712[(3'h5):(2'h2)] >>> reg675) ?
                      wire651 : reg704)) ?
                  reg720[(3'h4):(2'h2)] : $signed($signed($unsigned($unsigned(reg765)))));
              reg772 <= {reg732[(3'h7):(3'h7)]};
            end
          else
            begin
              reg770 <= (^~((~reg740) || (reg661[(4'he):(4'hc)] ~^ (+(forvar760 >> reg98)))));
            end
        end
      else
        begin
          for (forvar760 = (1'h0); (forvar760 < (3'h4)); forvar760 = (forvar760 + (1'h1)))
            begin
              reg762 = $signed($signed(reg264[(3'h4):(2'h2)]));
              reg763 = reg695[(5'h11):(2'h3)];
            end
          reg764 = $unsigned(({reg245[(2'h2):(1'h0)]} || (reg716 ?
              ((reg755 <<< (8'hb7)) ?
                  {reg751, reg234} : {reg716,
                      reg716}) : (reg698[(4'hd):(4'ha)] != (!wire434)))));
          if (reg762)
            begin
              reg765 = $signed((reg757[(2'h3):(2'h3)] ?
                  (|reg763) : ($signed((reg675 || wire702)) ?
                      reg755 : (reg716 <<< reg755))));
              reg768 = (($unsigned($unsigned($unsigned(reg224))) << ($unsigned({reg667,
                      (8'ha8)}) + (!reg680[(3'h4):(3'h4)]))) ?
                  reg96 : ((7'h45) + $signed((8'hac))));
              reg770 <= {{$signed(reg699[(4'ha):(2'h3)]), $unsigned(reg755)}};
              reg772 <= {(((reg753 >> $signed(reg221)) < reg122[(4'h9):(3'h4)]) ?
                      wire89 : (|$signed({wire124})))};
              reg773 <= reg245[(3'h6):(3'h5)];
            end
          else
            begin
              reg766 <= ($unsigned(reg766) + (~(7'h44)));
              reg768 = ($signed((((^(8'ha7)) * reg749) ?
                  $unsigned({reg261,
                      reg122}) : (7'h48))) == ((~^$unsigned((~&reg724))) & ($unsigned(reg710) ?
                  $signed((forvar756 << reg96)) : (~^$unsigned(reg755)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg774 = (!((^(~$unsigned(reg773))) ? reg698 : {$signed({reg98})}));
      for (forvar775 = (1'h0); (forvar775 < (3'h4)); forvar775 = (forvar775 + (1'h1)))
        begin
          if ({reg733[(1'h0):(1'h0)]})
            begin
              reg776 <= reg767[(1'h1):(1'h0)];
              reg777 = (({$signed(reg686), (8'ha1)} ?
                      $signed({wire702,
                          $unsigned(reg96)}) : (reg234[(4'he):(4'hc)] ?
                          {reg759[(4'hc):(1'h0)]} : (reg689[(3'h5):(3'h4)] && (|reg679)))) ?
                  ((|(reg759 != (forvar775 ? reg258 : reg772))) ?
                      $unsigned(reg744) : reg705) : $unsigned((reg229[(4'h9):(1'h1)] ?
                      $unsigned(reg226) : $signed((~|(7'h46))))));
              reg778 = $signed($unsigned((reg126 ?
                  (reg667 ?
                      {reg696, reg110} : (reg758 ? reg694 : reg709)) : (reg721 ?
                      (8'ha5) : {reg123}))));
              reg779 <= (~&(($unsigned((~&reg699)) & reg708[(3'h5):(2'h3)]) ?
                  ((reg700 ? $unsigned((8'hb9)) : $unsigned(reg241)) ?
                      $unsigned(reg661[(4'h9):(3'h7)]) : reg712) : $signed(wire702)));
            end
          else
            begin
              reg776 <= (($unsigned(reg126) ?
                      $signed(reg689[(5'h10):(1'h1)]) : (reg122[(4'h8):(3'h4)] >> wire91[(3'h6):(3'h6)])) ?
                  ((($unsigned(reg109) ?
                      (wire745 * (8'ha9)) : reg699[(3'h4):(2'h3)]) * $unsigned(reg224[(5'h13):(4'he)])) ^ ({(8'hb4)} ^ $signed((^~reg777)))) : reg245[(2'h2):(2'h2)]);
              reg779 <= (!$signed((|reg218[(2'h2):(1'h1)])));
              reg780 <= wire89[(1'h0):(1'h0)];
              reg781 <= (reg732[(1'h1):(1'h1)] ?
                  ({wire745} <= (reg234[(1'h1):(1'h0)] ?
                      $unsigned((reg724 >= wire433)) : reg712[(4'hb):(1'h1)])) : (&reg671));
            end
          reg782 = $unsigned($unsigned((7'h44)));
        end
    end
  always
    @(posedge clk) begin
      for (forvar783 = (1'h0); (forvar783 < (1'h0)); forvar783 = (forvar783 + (1'h1)))
        begin
          for (forvar784 = (1'h0); (forvar784 < (2'h2)); forvar784 = (forvar784 + (1'h1)))
            begin
              reg785 = $signed($unsigned((^~$signed((reg245 ?
                  reg780 : (7'h44))))));
              reg786 <= reg720[(4'h9):(1'h1)];
            end
          reg787 = (wire433[(1'h1):(1'h0)] ^ $signed(reg226));
        end
      reg788 <= $unsigned($signed((+$unsigned(reg732))));
      for (forvar789 = (1'h0); (forvar789 < (1'h1)); forvar789 = (forvar789 + (1'h1)))
        begin
          for (forvar790 = (1'h0); (forvar790 < (2'h2)); forvar790 = (forvar790 + (1'h1)))
            begin
              reg791 <= (~^$unsigned(reg749));
              reg792 = wire662;
              reg793 = $signed($unsigned({(((8'ha2) <= reg721) ?
                      $unsigned((7'h41)) : forvar783[(5'h10):(2'h3)])}));
              reg794 = $unsigned((reg767 != (wire651[(2'h3):(2'h2)] ?
                  ((reg786 ?
                      reg773 : reg710) ^ (~&reg779)) : ($signed(reg695) * $signed(reg680)))));
              reg795 <= (~^(reg713 ^~ {reg698,
                  (^~(reg234 ? reg218 : reg680))}));
            end
          for (forvar796 = (1'h0); (forvar796 < (1'h0)); forvar796 = (forvar796 + (1'h1)))
            begin
              reg797 = (~&($signed($signed(wire702[(3'h6):(3'h4)])) < reg684[(4'h9):(1'h0)]));
              reg798 <= $signed(($unsigned({(reg708 ? (8'ha8) : reg792),
                  wire702}) || $unsigned(reg684)));
            end
          reg799 <= reg767;
          if ((!(~reg659[(4'hb):(1'h1)])))
            begin
              reg800 <= (reg245 ?
                  reg705 : (!$unsigned(((^reg677) ?
                      (reg721 * reg707) : {(8'ha4), wire91}))));
              reg801 = reg221[(4'h8):(2'h2)];
              reg802 = {{($unsigned((reg657 ? reg679 : reg699)) ?
                          reg264 : ((|(8'ha2)) >= $unsigned(reg779))),
                      reg123}};
              reg803 <= $signed(reg264);
            end
          else
            begin
              reg801 = {(+$unsigned(({reg694,
                      (8'h9c)} >> wire649[(1'h1):(1'h1)]))),
                  (($unsigned({reg800, reg744}) & reg742) >= reg700)};
              reg802 = {reg226};
              reg804 = $unsigned(reg780[(5'h11):(3'h5)]);
            end
          for (forvar805 = (1'h0); (forvar805 < (1'h1)); forvar805 = (forvar805 + (1'h1)))
            begin
              reg806 <= reg750[(4'h9):(4'h8)];
            end
        end
      if (wire662)
        begin
          for (forvar807 = (1'h0); (forvar807 < (3'h4)); forvar807 = (forvar807 + (1'h1)))
            begin
              reg808 = reg766[(3'h6):(2'h2)];
              reg809 <= $signed($signed($signed((reg101[(4'he):(4'ha)] ?
                  (8'hb2) : wire216[(2'h2):(1'h1)]))));
            end
          reg810 = (!((^reg652) != (reg258[(1'h0):(1'h0)] ^~ reg659)));
          reg811 = ($unsigned({$unsigned($signed(reg739)),
                  (wire434[(3'h5):(2'h2)] * $unsigned(reg793))}) ?
              wire745[(2'h2):(1'h0)] : {(8'ha8), reg734[(1'h0):(1'h0)]});
          reg812 <= (8'hb1);
          for (forvar813 = (1'h0); (forvar813 < (2'h2)); forvar813 = (forvar813 + (1'h1)))
            begin
              reg814 = (&reg253);
              reg815 = reg794;
              reg816 <= ((((~&$unsigned(reg652)) | $signed(reg716)) ?
                      (($unsigned((8'hb4)) ? {(8'h9d)} : $unsigned(forvar805)) ?
                          ((^~wire662) ?
                              (reg264 >> reg101) : $signed(reg739)) : reg705) : (~&reg709)) ?
                  (8'h9e) : $signed(reg794[(4'ha):(4'h8)]));
              reg817 <= ((~&(!$signed($unsigned(forvar805)))) != $unsigned(($unsigned((reg758 ?
                      reg109 : reg811)) ?
                  {(reg122 >>> reg793)} : $signed($signed(reg664)))));
            end
        end
      else
        begin
          if ($unsigned((!(reg766[(3'h6):(3'h6)] ?
              reg680 : {((8'hac) | (8'ha1)), (reg116 ? reg248 : (7'h41))}))))
            begin
              reg807 <= reg713[(3'h4):(3'h4)];
              reg808 = reg803;
              reg809 <= (~{(&reg695[(2'h3):(2'h2)]),
                  $signed((((7'h42) ? reg678 : (8'ha1)) << {reg761}))});
            end
          else
            begin
              reg807 <= $signed(($signed($signed((reg117 <<< wire745))) == $unsigned($unsigned(reg720[(4'hb):(4'h8)]))));
              reg809 <= $signed($signed($unsigned((+(reg803 << reg226)))));
              reg810 = (~|({{(reg667 ^ reg236)}} || ({(reg674 - reg716)} >> (|(reg781 ?
                  (8'h9d) : (7'h44))))));
            end
        end
    end
  assign wire818 = (reg712 <<< $unsigned($unsigned(reg264[(3'h4):(3'h4)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module435  (y, clk, wire440, wire439, wire438, wire437, wire436);
  output wire [(32'hb21):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire440;
  input wire [(5'h15):(1'h0)] wire439;
  input wire signed [(5'h14):(1'h0)] wire438;
  input wire [(2'h3):(1'h0)] wire437;
  input wire [(5'h13):(1'h0)] wire436;
  wire signed [(5'h13):(1'h0)] wire627;
  wire signed [(5'h16):(1'h0)] wire540;
  wire signed [(2'h2):(1'h0)] wire539;
  wire signed [(4'h9):(1'h0)] wire523;
  wire signed [(4'h8):(1'h0)] wire522;
  wire signed [(5'h14):(1'h0)] wire521;
  wire signed [(4'h8):(1'h0)] wire498;
  wire [(2'h3):(1'h0)] wire497;
  wire [(3'h7):(1'h0)] wire445;
  wire signed [(2'h3):(1'h0)] wire441;
  reg signed [(4'h9):(1'h0)] reg640 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg646 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg643 = (1'h0);
  reg [(5'h10):(1'h0)] reg636 = (1'h0);
  reg [(5'h15):(1'h0)] reg634 = (1'h0);
  reg [(2'h3):(1'h0)] reg631 = (1'h0);
  reg [(4'hf):(1'h0)] reg628 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg621 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg617 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg613 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg620 = (1'h0);
  reg [(5'h14):(1'h0)] reg618 = (1'h0);
  reg [(4'he):(1'h0)] reg614 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg610 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg609 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg604 = (1'h0);
  reg [(3'h5):(1'h0)] reg601 = (1'h0);
  reg signed [(4'he):(1'h0)] reg599 = (1'h0);
  reg [(2'h2):(1'h0)] reg597 = (1'h0);
  reg [(3'h4):(1'h0)] reg596 = (1'h0);
  reg [(2'h2):(1'h0)] reg592 = (1'h0);
  reg signed [(4'he):(1'h0)] reg591 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg590 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg588 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg587 = (1'h0);
  reg [(3'h6):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg580 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg577 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg576 = (1'h0);
  reg [(5'h16):(1'h0)] reg574 = (1'h0);
  reg [(3'h7):(1'h0)] reg573 = (1'h0);
  reg [(5'h11):(1'h0)] reg570 = (1'h0);
  reg [(5'h16):(1'h0)] reg569 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg565 = (1'h0);
  reg [(4'he):(1'h0)] reg562 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg561 = (1'h0);
  reg [(4'hb):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg554 = (1'h0);
  reg [(4'hb):(1'h0)] reg549 = (1'h0);
  reg [(4'hf):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg550 = (1'h0);
  reg [(5'h10):(1'h0)] reg547 = (1'h0);
  reg [(5'h12):(1'h0)] reg546 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg541 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg535 = (1'h0);
  reg [(4'he):(1'h0)] reg533 = (1'h0);
  reg [(4'hb):(1'h0)] reg532 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg530 = (1'h0);
  reg [(5'h15):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg524 = (1'h0);
  reg [(5'h14):(1'h0)] reg520 = (1'h0);
  reg [(5'h13):(1'h0)] reg516 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg515 = (1'h0);
  reg [(3'h4):(1'h0)] reg513 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg511 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg508 = (1'h0);
  reg [(2'h3):(1'h0)] reg507 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg506 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg505 = (1'h0);
  reg [(5'h11):(1'h0)] reg502 = (1'h0);
  reg [(3'h7):(1'h0)] reg501 = (1'h0);
  reg [(4'h9):(1'h0)] reg496 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg493 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg489 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg488 = (1'h0);
  reg [(3'h5):(1'h0)] reg486 = (1'h0);
  reg [(5'h16):(1'h0)] reg484 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg478 = (1'h0);
  reg [(5'h10):(1'h0)] reg477 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg476 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg474 = (1'h0);
  reg [(3'h5):(1'h0)] reg470 = (1'h0);
  reg [(5'h17):(1'h0)] reg468 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg467 = (1'h0);
  reg [(3'h4):(1'h0)] reg466 = (1'h0);
  reg [(4'hf):(1'h0)] reg463 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg462 = (1'h0);
  reg [(5'h15):(1'h0)] reg461 = (1'h0);
  reg [(5'h13):(1'h0)] reg460 = (1'h0);
  reg [(2'h3):(1'h0)] reg459 = (1'h0);
  reg [(5'h15):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg455 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg453 = (1'h0);
  reg [(5'h16):(1'h0)] reg451 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg450 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg449 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg448 = (1'h0);
  reg [(4'hb):(1'h0)] reg443 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg442 = (1'h0);
  reg [(4'he):(1'h0)] reg648 = (1'h0);
  reg [(3'h4):(1'h0)] forvar647 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg645 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar644 = (1'h0);
  reg [(4'hc):(1'h0)] reg642 = (1'h0);
  reg [(5'h15):(1'h0)] reg641 = (1'h0);
  reg [(5'h15):(1'h0)] forvar640 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg639 = (1'h0);
  reg [(5'h13):(1'h0)] reg638 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg637 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg635 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg633 = (1'h0);
  reg [(4'ha):(1'h0)] reg632 = (1'h0);
  reg [(5'h12):(1'h0)] reg630 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar629 = (1'h0);
  reg [(4'he):(1'h0)] reg626 = (1'h0);
  reg [(4'hf):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg624 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg623 = (1'h0);
  reg [(5'h11):(1'h0)] forvar622 = (1'h0);
  reg [(3'h5):(1'h0)] reg619 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar617 = (1'h0);
  reg [(2'h2):(1'h0)] reg616 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg615 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar613 = (1'h0);
  reg [(3'h5):(1'h0)] reg612 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar611 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar608 = (1'h0);
  reg [(3'h7):(1'h0)] reg607 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg606 = (1'h0);
  reg [(4'h9):(1'h0)] reg605 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar603 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg602 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar600 = (1'h0);
  reg [(4'hd):(1'h0)] reg598 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg594 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar593 = (1'h0);
  reg [(4'h8):(1'h0)] reg584 = (1'h0);
  reg [(4'hc):(1'h0)] reg589 = (1'h0);
  reg [(3'h4):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg585 = (1'h0);
  reg [(5'h11):(1'h0)] forvar584 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg583 = (1'h0);
  reg [(4'he):(1'h0)] reg581 = (1'h0);
  reg [(4'hc):(1'h0)] reg579 = (1'h0);
  reg [(5'h14):(1'h0)] reg578 = (1'h0);
  reg [(5'h14):(1'h0)] forvar574 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg567 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg564 = (1'h0);
  reg [(3'h4):(1'h0)] forvar563 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg575 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg572 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg571 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg568 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar567 = (1'h0);
  reg [(5'h17):(1'h0)] reg566 = (1'h0);
  reg [(4'hf):(1'h0)] forvar564 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg563 = (1'h0);
  reg [(5'h10):(1'h0)] forvar560 = (1'h0);
  reg [(4'hd):(1'h0)] forvar557 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg556 = (1'h0);
  reg [(4'hd):(1'h0)] reg555 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg553 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar549 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg548 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg545 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg544 = (1'h0);
  reg [(4'h8):(1'h0)] reg543 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg542 = (1'h0);
  reg [(5'h17):(1'h0)] reg538 = (1'h0);
  reg [(5'h15):(1'h0)] forvar537 = (1'h0);
  reg [(5'h11):(1'h0)] reg536 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg534 = (1'h0);
  reg [(3'h4):(1'h0)] reg531 = (1'h0);
  reg [(4'ha):(1'h0)] forvar529 = (1'h0);
  reg [(4'hb):(1'h0)] forvar528 = (1'h0);
  reg [(4'hb):(1'h0)] reg527 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar525 = (1'h0);
  reg [(5'h15):(1'h0)] reg519 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg518 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar517 = (1'h0);
  reg [(5'h11):(1'h0)] reg514 = (1'h0);
  reg [(4'hf):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar510 = (1'h0);
  reg [(3'h6):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar504 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg503 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar500 = (1'h0);
  reg [(5'h13):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg473 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg495 = (1'h0);
  reg [(5'h16):(1'h0)] reg494 = (1'h0);
  reg [(2'h3):(1'h0)] reg492 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg491 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg490 = (1'h0);
  reg [(5'h11):(1'h0)] reg487 = (1'h0);
  reg signed [(4'he):(1'h0)] reg485 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg483 = (1'h0);
  reg [(3'h7):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg481 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg479 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg475 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar473 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg471 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar462 = (1'h0);
  reg [(4'hf):(1'h0)] reg469 = (1'h0);
  reg [(5'h15):(1'h0)] reg465 = (1'h0);
  reg [(5'h13):(1'h0)] reg464 = (1'h0);
  reg [(4'hf):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg457 = (1'h0);
  reg [(3'h5):(1'h0)] reg454 = (1'h0);
  reg [(2'h2):(1'h0)] reg452 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar447 = (1'h0);
  reg [(4'h8):(1'h0)] reg446 = (1'h0);
  reg [(5'h16):(1'h0)] reg444 = (1'h0);
  reg [(4'hb):(1'h0)] forvar442 = (1'h0);
  assign y = {wire627,
                 wire540,
                 wire539,
                 wire523,
                 wire522,
                 wire521,
                 wire498,
                 wire497,
                 wire445,
                 wire441,
                 reg640,
                 reg646,
                 reg643,
                 reg636,
                 reg634,
                 reg631,
                 reg628,
                 reg621,
                 reg617,
                 reg613,
                 reg620,
                 reg618,
                 reg614,
                 reg610,
                 reg609,
                 reg604,
                 reg601,
                 reg599,
                 reg597,
                 reg596,
                 reg592,
                 reg591,
                 reg590,
                 reg588,
                 reg587,
                 reg582,
                 reg580,
                 reg577,
                 reg576,
                 reg574,
                 reg573,
                 reg570,
                 reg569,
                 reg565,
                 reg562,
                 reg561,
                 reg559,
                 reg558,
                 reg554,
                 reg549,
                 reg552,
                 reg551,
                 reg550,
                 reg547,
                 reg546,
                 reg541,
                 reg535,
                 reg533,
                 reg532,
                 reg530,
                 reg526,
                 reg524,
                 reg520,
                 reg516,
                 reg515,
                 reg513,
                 reg511,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg502,
                 reg501,
                 reg496,
                 reg493,
                 reg489,
                 reg488,
                 reg486,
                 reg484,
                 reg478,
                 reg477,
                 reg476,
                 reg474,
                 reg470,
                 reg468,
                 reg467,
                 reg466,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg456,
                 reg455,
                 reg453,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg443,
                 reg442,
                 reg648,
                 forvar647,
                 reg645,
                 forvar644,
                 reg642,
                 reg641,
                 forvar640,
                 reg639,
                 reg638,
                 reg637,
                 reg635,
                 reg633,
                 reg632,
                 reg630,
                 forvar629,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 forvar622,
                 reg619,
                 forvar617,
                 reg616,
                 reg615,
                 forvar613,
                 reg612,
                 forvar611,
                 forvar608,
                 reg607,
                 reg606,
                 reg605,
                 forvar603,
                 reg602,
                 forvar600,
                 reg598,
                 reg595,
                 reg594,
                 forvar593,
                 reg584,
                 reg589,
                 reg586,
                 reg585,
                 forvar584,
                 reg583,
                 reg581,
                 reg579,
                 reg578,
                 forvar574,
                 reg567,
                 reg564,
                 forvar563,
                 reg575,
                 reg572,
                 reg571,
                 reg568,
                 forvar567,
                 reg566,
                 forvar564,
                 reg563,
                 forvar560,
                 forvar557,
                 reg556,
                 reg555,
                 reg553,
                 forvar549,
                 reg548,
                 reg545,
                 reg544,
                 reg543,
                 reg542,
                 reg538,
                 forvar537,
                 reg536,
                 reg534,
                 reg531,
                 forvar529,
                 forvar528,
                 reg527,
                 forvar525,
                 reg519,
                 reg518,
                 forvar517,
                 reg514,
                 reg512,
                 forvar510,
                 reg509,
                 forvar504,
                 reg503,
                 forvar500,
                 reg499,
                 reg473,
                 reg495,
                 reg494,
                 reg492,
                 reg491,
                 reg490,
                 reg487,
                 reg485,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 reg475,
                 forvar473,
                 reg472,
                 reg471,
                 forvar462,
                 reg469,
                 reg465,
                 reg464,
                 reg458,
                 reg457,
                 reg454,
                 reg452,
                 forvar447,
                 reg446,
                 reg444,
                 forvar442,
                 (1'h0)};
  assign wire441 = $signed({(^~$signed((~wire437))), {(8'hb2)}});
  always
    @(posedge clk) begin
      if ((wire439[(5'h12):(4'ha)] - wire436))
        begin
          reg442 <= ($signed((wire439[(3'h5):(1'h1)] > wire437[(1'h0):(1'h0)])) >>> (8'hb2));
        end
      else
        begin
          for (forvar442 = (1'h0); (forvar442 < (1'h0)); forvar442 = (forvar442 + (1'h1)))
            begin
              reg443 <= $signed(wire436[(3'h7):(1'h1)]);
            end
        end
      reg444 = (wire436 - (((forvar442[(4'h9):(3'h6)] ^ (8'hbb)) ?
              {(|wire437), $unsigned(reg443)} : (-wire436)) ?
          wire440 : reg442[(1'h0):(1'h0)]));
    end
  assign wire445 = $signed((^~reg443));
  always
    @(posedge clk) begin
      reg446 = wire437[(2'h3):(1'h1)];
    end
  always
    @(posedge clk) begin
      for (forvar447 = (1'h0); (forvar447 < (2'h3)); forvar447 = (forvar447 + (1'h1)))
        begin
          if (forvar447[(4'h9):(4'h9)])
            begin
              reg448 <= (~(+(((!reg443) ?
                      (wire438 < forvar447) : reg442[(4'ha):(1'h1)]) ?
                  ($signed(wire441) && wire439) : ((&wire439) >>> $unsigned((7'h49))))));
              reg449 <= $signed((reg442 ?
                  ((reg442 + $unsigned(forvar447)) ?
                      ((~^forvar447) ^ $unsigned((8'hb9))) : wire436[(1'h0):(1'h0)]) : $unsigned(wire439)));
              reg450 <= ({$unsigned((!reg448)), wire438} ?
                  wire445[(2'h2):(2'h2)] : ({wire441} & wire437[(2'h2):(1'h0)]));
            end
          else
            begin
              reg448 <= reg448[(4'h8):(1'h1)];
            end
          if ((~^wire440))
            begin
              reg451 <= $signed((~^($signed((~&wire445)) ?
                  ((forvar447 ? reg449 : wire445) ?
                      (reg443 ?
                          (8'hae) : reg442) : reg449[(4'h9):(4'h9)]) : {(wire445 ?
                          reg443 : reg450),
                      reg449})));
              reg452 = reg442;
              reg453 <= ((^~$signed(($unsigned(wire441) ?
                  (wire441 ^~ wire440) : $signed(wire436)))) - forvar447[(2'h2):(1'h1)]);
              reg454 = ({(^~($signed(reg442) <= $unsigned(reg448)))} ?
                  {$unsigned(($unsigned(wire440) ?
                          $unsigned(reg449) : (~|wire436)))} : {$unsigned($signed($signed(reg443))),
                      (reg448[(3'h5):(3'h5)] <<< wire441)});
            end
          else
            begin
              reg451 <= $signed((forvar447 ? $signed(wire438) : (^reg453)));
              reg452 = $signed({(((forvar447 <= wire438) ?
                      $unsigned(reg453) : (~&reg453)) - {(reg453 < wire440)})});
              reg454 = wire439[(2'h2):(1'h1)];
            end
          if ((({($signed(forvar447) * (wire439 | reg443)), {reg442, wire439}} ?
                  $signed((((8'hba) ? reg449 : reg452) | (wire441 ?
                      reg452 : wire439))) : ($signed((forvar447 ?
                      reg449 : reg454)) >= (((8'hb7) ? (8'ha6) : forvar447) ?
                      reg452[(1'h1):(1'h1)] : wire441[(2'h3):(1'h1)]))) ?
              {$signed((|(^(7'h44))))} : (~|(+(-((7'h41) ?
                  forvar447 : (8'hb3)))))))
            begin
              reg455 <= $unsigned(wire438);
              reg456 <= reg450[(2'h2):(2'h2)];
            end
          else
            begin
              reg457 = wire436;
              reg458 = (wire436 * (reg443 ?
                  $unsigned($signed($unsigned(reg443))) : (&((&reg443) >>> (8'hac)))));
              reg459 <= reg456;
            end
          reg460 <= (~(($signed((reg451 & wire437)) ?
                  ($unsigned(reg451) ?
                      ((7'h44) & wire438) : (reg456 <= (8'hb7))) : ($signed((8'hbc)) ?
                      $signed((8'hb0)) : wire445)) ?
              {(~^$unsigned(wire440))} : ((reg442 ?
                  {reg449,
                      wire436} : $unsigned(reg449)) <= (&$unsigned(reg456)))));
        end
      reg461 <= $unsigned(($signed((wire436[(4'hf):(4'h9)] > $unsigned(wire440))) != (&wire438[(4'hd):(4'hb)])));
      if (({(reg448[(1'h0):(1'h0)] ?
              $signed((reg461 ? reg443 : reg452)) : (~(7'h46))),
          $signed(((!reg456) ?
              $signed(reg456) : (reg442 ?
                  (8'haf) : reg442)))} >= reg448[(1'h0):(1'h0)]))
        begin
          if (reg456[(1'h1):(1'h1)])
            begin
              reg462 <= (&reg450[(1'h0):(1'h0)]);
              reg463 <= reg450;
            end
          else
            begin
              reg462 <= $unsigned((((reg443[(4'ha):(4'ha)] ?
                      (~&reg455) : (~|wire437)) >>> ($unsigned(reg449) > reg463[(2'h2):(1'h1)])) ?
                  $signed(((reg448 << reg459) ?
                      (wire445 * (8'hb7)) : $signed(reg451))) : $unsigned((8'hb4))));
              reg463 <= $signed($unsigned($signed(($unsigned(reg462) > $unsigned(wire436)))));
              reg464 = reg460;
              reg465 = reg452[(1'h0):(1'h0)];
              reg466 <= ((8'h9f) & $unsigned((^wire440)));
            end
          reg467 <= (reg462 ? forvar447 : $signed(reg458[(4'hc):(4'hc)]));
          reg468 <= {((-($unsigned(reg448) - {reg457})) ?
                  ($signed(reg463[(4'he):(4'hd)]) & $unsigned($signed(reg454))) : (~(~|(wire436 ~^ reg455))))};
          reg469 = {($signed(((|reg459) ? {reg455} : (~&wire436))) << reg455),
              reg463};
        end
      else
        begin
          for (forvar462 = (1'h0); (forvar462 < (2'h3)); forvar462 = (forvar462 + (1'h1)))
            begin
              reg463 <= ((reg453 * reg463[(4'ha):(3'h5)]) ?
                  reg451 : {(wire437[(1'h0):(1'h0)] < (wire439[(4'hc):(3'h5)] ?
                          (8'hab) : wire439))});
              reg466 <= reg468[(4'h9):(3'h7)];
              reg467 <= ($signed(reg457[(5'h10):(2'h3)]) ?
                  reg457 : $signed(($unsigned((7'h48)) ?
                      ($unsigned(reg450) ?
                          $unsigned(reg451) : $unsigned(reg442)) : $unsigned((forvar462 ?
                          reg448 : wire439)))));
            end
          reg469 = (reg468[(1'h1):(1'h0)] << $unsigned($unsigned(reg456)));
          reg470 <= reg466;
          reg471 = ({wire436} ?
              $unsigned({((reg465 ? wire437 : reg448) >= (wire441 ?
                      wire436 : (8'hb8)))}) : wire440);
        end
      reg472 = $unsigned((+((~(8'hbb)) <= ({wire436} * $unsigned(wire445)))));
      if (reg448)
        begin
          for (forvar473 = (1'h0); (forvar473 < (2'h2)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 <= ({reg455, reg450} ?
                  $signed($unsigned(reg472[(2'h3):(2'h2)])) : reg461);
              reg475 = ($signed($unsigned((reg467[(4'h9):(1'h1)] ?
                      $unsigned(forvar447) : reg461[(3'h4):(1'h0)]))) ?
                  $unsigned($unsigned(reg468)) : {(^$signed({reg461, reg455})),
                      ({$unsigned(reg464), (-reg474)} ?
                          (~^$unsigned(reg454)) : $unsigned({wire439,
                              reg454}))});
              reg476 <= forvar473[(1'h0):(1'h0)];
              reg477 <= ((($unsigned(forvar447) > $unsigned($signed(reg459))) | $unsigned(reg468[(1'h0):(1'h0)])) < wire440);
              reg478 <= reg450[(1'h1):(1'h0)];
            end
          reg479 = $unsigned($unsigned(({$signed(wire438),
              $signed((8'hb6))} != reg459)));
          if ($unsigned(reg471[(4'ha):(3'h4)]))
            begin
              reg480 = ($signed(reg453) ?
                  (&{$signed(reg454), (!$unsigned(reg451))}) : {{reg453}});
              reg481 = $signed(reg442[(4'h9):(3'h5)]);
              reg482 = $signed(reg463);
              reg483 = {(!$signed(($signed(reg443) ? (~^(7'h41)) : reg463))),
                  ($signed(($unsigned((7'h49)) > (reg450 ?
                      reg469 : reg450))) ^~ (^{(~&reg476)}))};
            end
          else
            begin
              reg484 <= reg471[(5'h16):(1'h0)];
              reg485 = ($unsigned($unsigned($signed(((7'h49) == (8'had))))) & $unsigned((|$signed((forvar462 | reg448)))));
              reg486 <= $unsigned((~&{((reg463 && reg454) << reg458),
                  $unsigned((!forvar462))}));
              reg487 = $signed($unsigned(reg477[(4'he):(4'hc)]));
            end
          if (reg477)
            begin
              reg488 <= reg480;
              reg489 <= reg475;
            end
          else
            begin
              reg488 <= reg472;
              reg489 <= $signed((~(reg458 ~^ reg442[(2'h3):(1'h1)])));
              reg490 = {(((~^$signed(reg486)) ?
                      (reg481 ?
                          (wire440 ? reg476 : wire440) : ((7'h44) ?
                              reg468 : wire441)) : reg457[(3'h4):(1'h1)]) - forvar473)};
            end
          if ((!(($unsigned($unsigned(wire441)) ?
              $unsigned((wire438 ?
                  reg478 : (8'haa))) : reg443) * $unsigned((+reg466[(1'h0):(1'h0)])))))
            begin
              reg491 = reg480;
              reg492 = ({{$signed((~&reg484)),
                      ($signed(reg491) ?
                          ((8'hac) ?
                              reg466 : reg470) : {wire439})}} < reg468[(2'h2):(1'h1)]);
              reg493 <= ($unsigned((^((reg449 > reg469) || (reg481 != (7'h45))))) ?
                  (($unsigned((reg470 < reg456)) * (+((8'hbe) ~^ (7'h43)))) | ((8'hb8) ?
                      (~^(^~(8'h9e))) : (~^(wire436 < reg460)))) : ($unsigned($signed((!(7'h46)))) ?
                      ((&(reg474 ?
                          reg453 : reg470)) ^~ reg465) : $unsigned((reg488 < reg452[(1'h1):(1'h0)]))));
            end
          else
            begin
              reg493 <= $unsigned(reg458[(3'h7):(3'h7)]);
              reg494 = reg466;
              reg495 = (reg453[(1'h0):(1'h0)] & $unsigned((7'h41)));
              reg496 <= reg488[(3'h6):(2'h2)];
            end
        end
      else
        begin
          if ($signed((~((~^$signed(reg466)) | {reg465, reg451}))))
            begin
              reg473 = {(~|($signed($unsigned(forvar462)) << (~|((7'h48) ?
                      reg464 : reg468))))};
              reg475 = {(($signed($signed(reg488)) ?
                      reg463[(4'h8):(1'h1)] : $unsigned(reg452[(1'h1):(1'h0)])) >= {((|reg478) << wire438)}),
                  $signed(((^~$signed(wire439)) & $unsigned({(8'ha1),
                      reg490})))};
              reg476 <= $unsigned((8'hb3));
              reg479 = ($unsigned({{wire437},
                  reg471}) < (($unsigned(reg452[(2'h2):(1'h0)]) ?
                      wire437[(1'h0):(1'h0)] : (reg448[(4'ha):(1'h1)] ?
                          (reg449 ? reg486 : reg462) : reg479[(3'h5):(1'h1)])) ?
                  reg488[(1'h1):(1'h1)] : $signed(((reg481 ?
                      reg474 : wire438) & reg474[(4'he):(4'hd)]))));
              reg484 <= reg475;
            end
          else
            begin
              reg474 <= reg494[(4'hc):(1'h0)];
              reg475 = ($unsigned(($unsigned((!(8'h9c))) ?
                  reg463[(4'h9):(4'h9)] : {$unsigned(reg477),
                      (~reg457)})) != $unsigned($unsigned((7'h48))));
              reg476 <= $signed(reg488[(3'h7):(2'h3)]);
              reg477 <= $unsigned(reg454[(1'h1):(1'h0)]);
              reg478 <= wire437;
            end
        end
    end
  assign wire497 = {((~&reg477) > reg460[(2'h3):(2'h2)])};
  assign wire498 = (reg466 ~^ (reg460[(4'he):(3'h6)] * (^reg462)));
  always
    @(posedge clk) begin
      reg499 = $unsigned(((|reg496[(1'h0):(1'h0)]) ?
          (-$unsigned(((8'hb0) ~^ reg461))) : (~^(|$unsigned((8'hbf))))));
      for (forvar500 = (1'h0); (forvar500 < (1'h1)); forvar500 = (forvar500 + (1'h1)))
        begin
          reg501 <= $unsigned({reg470[(3'h4):(3'h4)], (8'ha3)});
          reg502 <= (|$signed((8'hab)));
          reg503 = reg476;
          for (forvar504 = (1'h0); (forvar504 < (3'h4)); forvar504 = (forvar504 + (1'h1)))
            begin
              reg505 <= {(~|$unsigned(((^reg460) < {reg442, wire438}))),
                  ($unsigned(reg463[(1'h1):(1'h0)]) ?
                      ((|$signed(reg466)) ?
                          wire441[(1'h0):(1'h0)] : $unsigned(reg456)) : (($unsigned(reg459) >= $unsigned(reg477)) ?
                          {(reg442 ? (7'h40) : reg493)} : ({reg453} ?
                              forvar500 : $unsigned(reg484))))};
              reg506 <= reg456;
            end
        end
      reg507 <= {($unsigned((reg449[(4'h8):(3'h6)] ?
                  (reg466 <<< wire497) : (+forvar500))) ?
              (&(~$unsigned(reg499))) : $unsigned(($signed((8'h9e)) ~^ (reg450 ?
                  reg443 : reg460)))),
          (~(~&($unsigned((7'h42)) >> (!reg468))))};
      if ((((reg443 ?
                  ((-reg443) ? {wire439, wire445} : (&reg503)) : ({reg461} ?
                      reg459 : (reg503 ? wire445 : reg442))) ?
              reg461 : ($signed(reg488[(2'h2):(1'h1)]) ?
                  {$unsigned(reg474),
                      (reg470 ? (7'h43) : wire436)} : ((!reg456) + (8'ha0)))) ?
          reg460[(4'hc):(3'h4)] : (({(reg466 ^~ reg451)} >>> $unsigned($unsigned(wire441))) * (~&{wire436[(4'h9):(4'h9)],
              (reg503 ? reg486 : (8'h9c))}))))
        begin
          reg508 <= ($signed((($signed(reg466) != {reg488, reg448}) ?
              $signed(reg459) : wire440[(4'hf):(4'hd)])) ^~ wire437);
          reg509 = $signed(({(8'hbc)} <= wire438));
          for (forvar510 = (1'h0); (forvar510 < (1'h0)); forvar510 = (forvar510 + (1'h1)))
            begin
              reg511 <= (reg453 ?
                  $signed((reg493 ?
                      $unsigned((~&wire439)) : $signed(wire445[(3'h6):(1'h0)]))) : $unsigned(reg476[(1'h0):(1'h0)]));
              reg512 = ($unsigned((-(reg501[(1'h0):(1'h0)] ?
                  $signed(reg442) : $unsigned(reg470)))) && ((wire441[(2'h3):(2'h2)] >> ((reg489 | reg466) > (reg474 < (8'had)))) ?
                  ($signed((reg463 >> reg459)) * ((-forvar500) && (wire498 ?
                      reg489 : reg468))) : reg484));
              reg513 <= $unsigned(wire497);
            end
          if (reg470[(3'h4):(3'h4)])
            begin
              reg514 = ((7'h44) ? (~^reg476[(1'h0):(1'h0)]) : wire438);
              reg515 <= $signed((~^$unsigned({$signed(reg456)})));
              reg516 <= $unsigned((((reg474[(1'h0):(1'h0)] ?
                      {reg505} : (!reg509)) & ((forvar500 ?
                      forvar510 : reg513) || (reg496 >> reg443))) ?
                  (^~reg512[(1'h0):(1'h0)]) : reg484[(4'h8):(3'h6)]));
            end
          else
            begin
              reg515 <= ({(($unsigned(reg459) <<< (forvar510 ?
                      reg505 : wire439)) << $unsigned($unsigned(reg489))),
                  ((~^(~^(8'hb6))) ?
                      reg466[(2'h3):(1'h1)] : reg493)} > $signed(reg507));
            end
          for (forvar517 = (1'h0); (forvar517 < (2'h2)); forvar517 = (forvar517 + (1'h1)))
            begin
              reg518 = (&$unsigned((|$signed((!reg484)))));
              reg519 = $signed($unsigned(reg499[(4'hf):(1'h0)]));
              reg520 <= (7'h42);
            end
        end
      else
        begin
          reg508 <= reg518;
        end
    end
  assign wire521 = ((($signed((7'h41)) ?
                           reg511[(3'h4):(3'h4)] : ((reg515 || (8'ha5)) && (7'h49))) ?
                       (({(8'ha8), reg461} ?
                           $unsigned(reg477) : {reg484,
                               reg477}) ^ reg462) : (((reg516 ?
                               (8'hab) : reg513) ~^ reg516[(5'h11):(4'he)]) ?
                           reg513 : (reg520[(1'h0):(1'h0)] ?
                               (7'h43) : $signed((8'haa))))) >= $unsigned((~|((~^reg513) ?
                       (reg451 * (8'ha8)) : $signed((8'hab))))));
  assign wire522 = wire440[(4'hb):(4'h9)];
  assign wire523 = ((^~wire440[(4'hd):(2'h3)]) ?
                       $unsigned($unsigned(($unsigned(reg493) ?
                           wire436[(1'h1):(1'h1)] : reg508[(3'h4):(2'h2)]))) : {($unsigned(((8'ha7) ?
                               reg507 : wire498)) >= reg496[(4'h9):(4'h8)]),
                           $unsigned(wire521[(4'hd):(4'h9)])});
  always
    @(posedge clk) begin
      reg524 <= $unsigned((reg513 >>> (8'had)));
      for (forvar525 = (1'h0); (forvar525 < (3'h4)); forvar525 = (forvar525 + (1'h1)))
        begin
          reg526 <= (((reg496[(4'h9):(3'h5)] | ($unsigned(reg502) ?
                      (reg484 >= (7'h43)) : (!reg524))) ?
                  (|$unsigned((reg463 == reg484))) : (^reg496[(1'h1):(1'h1)])) ?
              $unsigned(($signed($unsigned(reg511)) ?
                  (&(8'h9f)) : (~(~^reg453)))) : ((~$unsigned((reg450 <<< wire522))) == (&((|reg515) ?
                  (wire440 <<< reg516) : wire438))));
          reg527 = reg489[(1'h0):(1'h0)];
        end
      for (forvar528 = (1'h0); (forvar528 < (1'h1)); forvar528 = (forvar528 + (1'h1)))
        begin
          for (forvar529 = (1'h0); (forvar529 < (2'h2)); forvar529 = (forvar529 + (1'h1)))
            begin
              reg530 <= forvar525[(2'h2):(1'h1)];
              reg531 = (wire441[(2'h2):(1'h0)] ?
                  (wire437 ?
                      (reg477[(4'ha):(4'ha)] ?
                          $signed(wire438[(4'hf):(1'h0)]) : wire437[(2'h3):(1'h0)]) : {reg526[(4'hb):(3'h6)]}) : {(($signed(reg496) ?
                              $unsigned(reg527) : (reg524 ? reg463 : reg515)) ?
                          wire437 : $unsigned({(7'h46)})),
                      reg506});
              reg532 <= reg506;
              reg533 <= (8'hb2);
              reg534 = wire441;
            end
          reg535 <= $signed({(({(7'h49),
                  wire497} ^ reg532) == (&reg455[(5'h12):(4'h9)])),
              {wire521, ({wire437} ? $signed(reg448) : $signed((8'hb8)))}});
          reg536 = (!reg507[(1'h1):(1'h1)]);
        end
      for (forvar537 = (1'h0); (forvar537 < (1'h1)); forvar537 = (forvar537 + (1'h1)))
        begin
          reg538 = (wire441[(1'h1):(1'h1)] ?
              (reg524 ?
                  $unsigned(((|forvar529) >> ((7'h48) * reg501))) : $unsigned(wire523[(2'h2):(1'h0)])) : $unsigned($signed(reg450)));
        end
    end
  assign wire539 = {reg511,
                       ((reg448 ?
                               ($unsigned(reg524) ?
                                   reg488[(3'h4):(2'h3)] : $unsigned(wire498)) : reg489) ?
                           ($unsigned((~&wire523)) >> reg443[(1'h0):(1'h0)]) : reg463)};
  assign wire540 = ($signed((8'hae)) ?
                       $signed($signed($unsigned(reg459))) : reg455[(4'h9):(1'h1)]);
  always
    @(posedge clk) begin
      if ($unsigned($signed(reg443[(3'h5):(1'h1)])))
        begin
          if (((~&{reg456}) ?
              $signed((reg532[(4'ha):(4'ha)] ~^ $signed(reg535))) : (-reg515)))
            begin
              reg541 <= (^$unsigned($signed($unsigned(wire438))));
              reg542 = wire540[(5'h16):(3'h7)];
              reg543 = $signed(reg524);
              reg544 = $unsigned(({reg467, {(wire540 ? reg443 : reg532)}} ?
                  ((~^reg451[(4'h8):(4'h8)]) ?
                      {reg516[(3'h7):(3'h6)]} : $signed($signed(reg459))) : ($unsigned(reg462[(4'ha):(2'h3)]) != ($signed(wire445) ?
                      (reg462 ? wire497 : reg453) : $signed((8'hb5))))));
            end
          else
            begin
              reg542 = reg476;
            end
          if ($unsigned((reg511[(2'h3):(1'h1)] ?
              (reg486 ?
                  ((wire521 ~^ reg541) ^~ $signed(reg520)) : $unsigned({reg477,
                      (8'h9c)})) : (8'hba))))
            begin
              reg545 = $unsigned((wire540 ? reg526 : (~|reg463)));
            end
          else
            begin
              reg546 <= $signed(((!reg533[(4'hd):(4'h9)]) ?
                  $unsigned(wire437) : (!(~^(reg507 ? reg462 : reg526)))));
              reg547 <= (wire540[(4'h8):(4'h8)] ?
                  (~^$unsigned(($unsigned(reg515) <<< $signed(reg489)))) : (reg493 ?
                      (8'hb5) : reg544[(4'hf):(4'hb)]));
              reg548 = (^~wire522);
            end
          for (forvar549 = (1'h0); (forvar549 < (2'h3)); forvar549 = (forvar549 + (1'h1)))
            begin
              reg550 <= $unsigned(((reg520[(3'h6):(1'h1)] ?
                      $signed(reg478) : (8'hb1)) ?
                  reg505[(2'h3):(1'h0)] : $signed($unsigned((reg453 <= wire438)))));
              reg551 <= $signed(((reg526 < {{reg530}}) ?
                  $signed(reg526) : $unsigned((reg493[(3'h4):(1'h1)] >= (^~reg507)))));
              reg552 <= wire445;
            end
        end
      else
        begin
          reg542 = {((reg508 ?
                  ((forvar549 <<< wire539) ^ (reg496 ^ reg547)) : $signed(reg486[(2'h2):(2'h2)])) <<< $unsigned(wire522[(3'h5):(3'h4)]))};
          if ((-(-reg541[(2'h3):(2'h3)])))
            begin
              reg546 <= reg477[(1'h1):(1'h0)];
            end
          else
            begin
              reg546 <= reg474[(4'ha):(3'h4)];
              reg547 <= ((~^$signed((+(-(8'hb7))))) ?
                  ((^(wire438 ?
                      (wire439 ?
                          wire438 : reg515) : reg477[(4'h8):(4'h8)])) ^ $signed(($unsigned(reg459) ?
                      $unsigned((8'hac)) : (reg551 ?
                          reg508 : reg470)))) : reg476[(1'h1):(1'h0)]);
              reg549 <= $signed(($unsigned(wire522[(1'h0):(1'h0)]) ^~ {((reg508 ?
                          reg477 : reg548) ?
                      {wire441} : reg449)}));
            end
          if (((((&(reg513 == reg462)) || reg466) ?
                  (reg453[(2'h2):(1'h0)] ?
                      reg511[(3'h4):(1'h0)] : $unsigned($unsigned(reg449))) : reg468[(5'h10):(2'h2)]) ?
              $signed((~&(8'hb6))) : (^~$unsigned(reg449))))
            begin
              reg553 = reg502[(4'h8):(3'h4)];
              reg554 <= (^({$unsigned($signed(reg486)),
                  $signed(reg486)} >> (!{(reg466 && reg549),
                  (reg477 ? forvar549 : reg547)})));
            end
          else
            begin
              reg550 <= $signed((-reg477[(3'h7):(2'h3)]));
              reg553 = (wire498[(3'h4):(1'h0)] ?
                  {{(~&{reg530, reg541}),
                          $unsigned($signed(reg541))}} : (reg478[(1'h1):(1'h0)] ?
                      $signed(({wire440} ?
                          wire521[(1'h0):(1'h0)] : reg476[(1'h0):(1'h0)])) : $unsigned(reg496)));
              reg554 <= ((^reg450[(3'h6):(1'h0)]) ?
                  ((reg468[(4'h9):(3'h7)] ^~ ((reg449 ?
                          reg552 : (7'h4a)) >>> $signed(reg511))) ?
                      (-$signed(reg455)) : ($unsigned(wire522) >>> ($unsigned(wire497) ?
                          (reg451 << reg516) : (~^reg532)))) : (!$signed(reg486)));
              reg555 = (((wire497 ?
                      (~&reg532) : (&reg545)) <<< ($unsigned(wire540[(4'h8):(2'h3)]) != ((|reg489) ?
                      reg526[(4'ha):(3'h4)] : reg489[(3'h4):(2'h3)]))) ?
                  $signed(wire522[(1'h1):(1'h1)]) : reg443);
              reg556 = wire441;
            end
        end
      for (forvar557 = (1'h0); (forvar557 < (3'h4)); forvar557 = (forvar557 + (1'h1)))
        begin
          reg558 <= {(~^(!reg477[(4'ha):(3'h4)]))};
          reg559 <= ((^~$signed(($unsigned(reg553) ?
              $signed(reg488) : (reg513 ?
                  (8'hb2) : reg547)))) <<< $unsigned((($signed((7'h41)) ?
                  (|reg511) : $signed(reg555)) ?
              $unsigned({wire498}) : $unsigned(reg524))));
        end
      for (forvar560 = (1'h0); (forvar560 < (2'h3)); forvar560 = (forvar560 + (1'h1)))
        begin
          reg561 <= $signed({{$unsigned((reg477 ? reg549 : reg547))},
              reg555[(3'h5):(3'h4)]});
        end
      reg562 <= $unsigned(wire540[(4'he):(1'h0)]);
      if ($unsigned($signed(forvar560)))
        begin
          reg563 = (~&reg449);
          for (forvar564 = (1'h0); (forvar564 < (1'h1)); forvar564 = (forvar564 + (1'h1)))
            begin
              reg565 <= $unsigned((($signed((^~(8'hb4))) ~^ $signed(reg555[(3'h7):(3'h6)])) ?
                  (((8'h9c) | {reg486}) ?
                      $signed(reg460) : reg549) : $signed({$unsigned((7'h43)),
                      $signed(reg543)})));
            end
          reg566 = $signed($unsigned(($signed($signed(reg455)) >> (&$unsigned(wire522)))));
          for (forvar567 = (1'h0); (forvar567 < (1'h0)); forvar567 = (forvar567 + (1'h1)))
            begin
              reg568 = ((8'hb5) >= {(8'hb5), (~|reg453[(1'h0):(1'h0)])});
              reg569 <= $unsigned((7'h47));
              reg570 <= (reg563 || (({$unsigned(reg449)} ?
                      reg566[(5'h15):(4'ha)] : ((wire497 >> (8'haa)) <<< $signed(reg462))) ?
                  reg442[(4'h9):(4'h9)] : wire540[(5'h13):(2'h3)]));
              reg571 = (~^forvar560);
              reg572 = $unsigned($signed(forvar564[(4'ha):(4'ha)]));
            end
          if (reg493[(4'h8):(2'h3)])
            begin
              reg573 <= $unsigned(reg484[(1'h1):(1'h1)]);
              reg574 <= {{reg463[(1'h1):(1'h0)],
                      (($signed(reg551) | ((8'ha0) ? reg507 : reg535)) ?
                          $unsigned((-reg568)) : reg477)}};
            end
          else
            begin
              reg575 = reg493[(3'h6):(1'h0)];
              reg576 <= $unsigned(({$signed((|wire540))} ?
                  $unsigned(($signed(reg507) ?
                      reg549[(1'h1):(1'h1)] : reg559)) : {(~^{reg488})}));
            end
        end
      else
        begin
          for (forvar563 = (1'h0); (forvar563 < (1'h0)); forvar563 = (forvar563 + (1'h1)))
            begin
              reg564 = reg575[(3'h5):(3'h5)];
              reg566 = (((~|{(&reg544), (reg466 > wire445)}) ?
                  (8'ha3) : (wire539 != ((reg556 != (7'h43)) > $unsigned((8'ha2))))) || {(7'h41)});
              reg567 = $signed({$unsigned(reg448[(2'h2):(2'h2)])});
              reg569 <= (($unsigned((reg451[(4'hf):(4'ha)] > $unsigned((8'haf)))) + $unsigned({reg442,
                      $signed(wire440)})) ?
                  (8'ha5) : reg565[(4'h8):(1'h0)]);
              reg571 = ($unsigned((reg443[(2'h3):(1'h1)] ?
                      (~reg478) : $signed($unsigned(reg484)))) ?
                  ($signed($signed((reg501 - wire441))) & reg542[(3'h4):(2'h2)]) : ($signed($unsigned(reg449[(3'h4):(1'h0)])) ?
                      reg508 : reg550[(5'h11):(4'he)]));
            end
          reg573 <= ((~|$unsigned($unsigned(wire445[(1'h0):(1'h0)]))) ?
              reg541[(4'ha):(1'h0)] : reg460[(3'h4):(2'h3)]);
          for (forvar574 = (1'h0); (forvar574 < (2'h2)); forvar574 = (forvar574 + (1'h1)))
            begin
              reg575 = (~reg453);
              reg576 <= $unsigned((($unsigned($signed((8'haf))) != $unsigned($unsigned((8'hbc)))) <<< (~reg451[(3'h7):(3'h7)])));
              reg577 <= {reg507[(1'h1):(1'h1)],
                  ((^(reg463[(4'hb):(1'h0)] ? $unsigned(reg563) : wire522)) ?
                      $unsigned($signed(wire445)) : {wire438})};
              reg578 = {reg577[(1'h1):(1'h0)]};
            end
          if ((8'hb8))
            begin
              reg579 = $unsigned({{(&(reg543 >> (7'h4a)))}});
            end
          else
            begin
              reg580 <= wire522;
              reg581 = $unsigned($unsigned($unsigned(({(7'h45)} <<< (~&(8'haf))))));
              reg582 <= ($unsigned((~&reg573[(1'h0):(1'h0)])) - (^($unsigned({reg493,
                      reg449}) ?
                  reg513 : ($unsigned(wire539) && $unsigned(wire436)))));
              reg583 = (reg442 ? $unsigned(reg547) : reg533);
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed((reg573 ?
          (~|reg496[(2'h2):(1'h1)]) : ($signed({reg515}) ?
              ((reg577 << reg530) <<< (reg463 ?
                  reg565 : reg535)) : $signed(reg449)))))
        begin
          for (forvar584 = (1'h0); (forvar584 < (1'h0)); forvar584 = (forvar584 + (1'h1)))
            begin
              reg585 = ((reg562[(4'hd):(2'h3)] == $signed($signed((8'hae)))) ?
                  $signed(reg453[(1'h1):(1'h1)]) : $unsigned($unsigned(reg477[(4'hd):(3'h4)])));
            end
          if ((^~wire540))
            begin
              reg586 = ((({reg533[(4'ha):(1'h1)], reg535} ?
                      $unsigned(reg546[(5'h10):(4'hc)]) : $unsigned((-reg526))) ?
                  ({(reg552 ^ wire439)} ?
                      $signed((reg443 | reg582)) : reg507[(2'h2):(1'h1)]) : (((reg468 <<< reg455) ?
                      {wire498} : (reg532 ?
                          reg577 : reg467)) ^~ reg550)) >= (+($unsigned((reg580 || reg585)) ?
                  (reg565[(4'hb):(4'ha)] ?
                      $signed(reg493) : $unsigned(wire497)) : (+$signed(reg549)))));
              reg587 <= reg574[(4'ha):(1'h1)];
              reg588 <= $signed($signed((~|reg532[(4'ha):(3'h4)])));
            end
          else
            begin
              reg586 = {((~$signed((reg532 ~^ (8'hae)))) & ($unsigned(reg569[(4'hc):(4'ha)]) ?
                      reg456[(5'h11):(5'h10)] : forvar584[(2'h2):(1'h0)])),
                  reg511[(1'h1):(1'h0)]};
              reg587 <= reg459[(2'h2):(1'h0)];
              reg588 <= $unsigned({$unsigned((reg533 ?
                      (~&reg476) : reg574[(4'hc):(3'h5)]))});
              reg589 = (($signed((reg573[(3'h7):(1'h1)] ?
                          $signed(reg577) : (reg587 ? reg456 : (7'h43)))) ?
                      wire498 : reg535) ?
                  {(((&reg453) || ((7'h41) << reg443)) ?
                          (((8'ha7) > reg467) && (forvar584 ?
                              reg496 : reg587)) : wire540),
                      $unsigned((~&(^wire523)))} : (reg508 ?
                      (reg456[(2'h2):(1'h0)] ?
                          ((~^reg580) ?
                              $unsigned((8'haf)) : reg513[(2'h2):(2'h2)]) : reg569) : {{(reg459 ?
                                  reg577 : wire498)}}));
            end
        end
      else
        begin
          reg584 = (~$unsigned((+((wire523 ? reg520 : (8'ha3)) ?
              (reg467 ? (8'hb2) : reg552) : {reg476, reg526}))));
          reg587 <= {(((~(|reg461)) ?
                  (reg461 ^~ $unsigned(reg573)) : (~reg489)) >> $unsigned((+(reg576 | (7'h46)))))};
          if ($signed((^(($unsigned(reg516) ?
                  $unsigned(reg484) : (reg508 <<< (8'h9d))) ?
              wire497[(2'h2):(1'h0)] : $unsigned({reg450})))))
            begin
              reg588 <= reg588;
              reg590 <= {$signed(({$signed(reg526),
                      {reg470, wire498}} <<< wire441)),
                  reg532};
              reg591 <= {wire540};
              reg592 <= ($unsigned((reg484[(2'h2):(2'h2)] ?
                  $unsigned(wire445) : $signed((^~wire441)))) + reg508);
            end
          else
            begin
              reg588 <= $signed(reg547);
              reg589 = ((reg587[(2'h2):(1'h1)] ?
                  (~|(reg459[(2'h3):(2'h2)] <<< (reg573 ?
                      reg443 : (8'ha0)))) : (((forvar584 ? reg558 : reg588) ?
                      reg461 : $signed(wire497)) - ((-wire437) ?
                      (reg488 <= wire523) : reg507[(1'h1):(1'h1)]))) == reg461[(4'hb):(2'h3)]);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar593 = (1'h0); (forvar593 < (2'h3)); forvar593 = (forvar593 + (1'h1)))
        begin
          if ((~$unsigned(($signed(((8'hbd) ? reg453 : wire445)) ?
              reg463 : {$signed((7'h48)), $unsigned(reg549)}))))
            begin
              reg594 = reg561[(2'h2):(1'h0)];
              reg595 = $signed($signed((!$signed(wire540[(1'h1):(1'h0)]))));
              reg596 <= $signed({reg576[(4'hf):(4'ha)],
                  ($unsigned((7'h49)) - ((8'ha1) ?
                      $unsigned(reg547) : {reg551}))});
              reg597 <= (7'h47);
            end
          else
            begin
              reg594 = reg442;
              reg595 = reg502;
              reg598 = ((8'h9f) | $unsigned($unsigned(reg506)));
              reg599 <= reg561[(2'h2):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar600 = (1'h0); (forvar600 < (2'h3)); forvar600 = (forvar600 + (1'h1)))
        begin
          reg601 <= (^reg468[(4'h8):(3'h5)]);
          reg602 = (($signed(reg550[(4'ha):(3'h5)]) < (|(reg524[(4'hd):(4'hc)] ?
              reg460 : (reg501 * reg597)))) * wire438[(3'h7):(1'h1)]);
          for (forvar603 = (1'h0); (forvar603 < (2'h3)); forvar603 = (forvar603 + (1'h1)))
            begin
              reg604 <= reg460;
              reg605 = (&(+(~&$unsigned(reg459[(2'h2):(1'h1)]))));
              reg606 = $signed({$signed((~^(8'hae)))});
            end
          reg607 = ((~^reg462) << (~reg459[(2'h3):(2'h3)]));
        end
      for (forvar608 = (1'h0); (forvar608 < (3'h4)); forvar608 = (forvar608 + (1'h1)))
        begin
          reg609 <= $unsigned(reg460);
          reg610 <= $unsigned((!$unsigned({{(7'h45), reg609}})));
        end
      for (forvar611 = (1'h0); (forvar611 < (1'h0)); forvar611 = (forvar611 + (1'h1)))
        begin
          reg612 = reg496;
        end
      if ((reg459[(1'h1):(1'h1)] ?
          (($unsigned((reg577 ? wire523 : wire440)) ?
                  ((8'hab) ^ $signed((7'h47))) : $unsigned($signed(reg476))) ?
              wire540[(4'h9):(4'h9)] : $unsigned($unsigned(((8'hbf) >> reg587)))) : $unsigned(((7'h41) ?
              {$unsigned(reg459)} : ({reg573, (8'h9c)} ?
                  reg587 : $signed(reg607))))))
        begin
          for (forvar613 = (1'h0); (forvar613 < (2'h3)); forvar613 = (forvar613 + (1'h1)))
            begin
              reg614 <= ($signed({$unsigned({reg541, reg459}),
                  $unsigned($signed(wire539))}) != $signed(reg455));
            end
          reg615 = ((reg526[(3'h4):(1'h0)] ?
                  (($signed(wire498) ?
                      (+reg550) : (8'hbb)) & ($signed(reg558) - $signed(reg552))) : $unsigned(({wire498} <= reg562[(4'h9):(3'h6)]))) ?
              (reg488[(3'h5):(1'h0)] * $signed((reg496 ?
                  {reg460} : $unsigned(reg614)))) : reg602[(2'h3):(1'h0)]);
          reg616 = (7'h44);
          for (forvar617 = (1'h0); (forvar617 < (2'h3)); forvar617 = (forvar617 + (1'h1)))
            begin
              reg618 <= reg515[(4'hc):(3'h7)];
              reg619 = reg484[(5'h16):(4'he)];
              reg620 <= reg463[(4'hb):(3'h7)];
            end
        end
      else
        begin
          reg613 <= (reg552[(2'h3):(1'h1)] ?
              $unsigned((wire439 << reg486[(2'h3):(2'h3)])) : $unsigned(wire521));
          reg614 <= reg524;
          if ($signed({reg451[(4'hb):(1'h1)]}))
            begin
              reg617 <= (~&reg484[(4'h8):(3'h5)]);
              reg618 <= $unsigned(reg486[(1'h1):(1'h0)]);
              reg620 <= {((reg535 || ((-(8'hbe)) - (reg552 && reg559))) >>> {$unsigned((reg617 * forvar613))}),
                  {{((reg486 << reg546) + reg488[(2'h3):(1'h0)])},
                      $signed(($unsigned(forvar608) ?
                          reg558 : $signed(reg450)))}};
              reg621 <= ((($signed($unsigned(reg533)) && {$signed(reg466)}) ?
                      (+wire445) : wire521) ?
                  wire439 : (~^reg468));
            end
          else
            begin
              reg617 <= (|((!$unsigned((reg612 ?
                  (8'hb3) : forvar603))) <<< reg615));
              reg618 <= (reg489 ?
                  {(~&(reg621[(2'h2):(1'h1)] ?
                          ((7'h46) | reg459) : $signed(reg496))),
                      forvar611} : $unsigned($signed(reg496[(2'h2):(2'h2)])));
              reg619 = (!reg442[(1'h0):(1'h0)]);
              reg620 <= forvar608[(4'hf):(2'h2)];
              reg621 <= reg574[(3'h4):(1'h0)];
            end
          for (forvar622 = (1'h0); (forvar622 < (1'h0)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 = ({((~^(wire539 == (8'had))) ^~ $signed(((8'hb1) ?
                          reg596 : reg530)))} ?
                  $signed({reg559[(3'h7):(1'h1)],
                      $unsigned($signed(reg554))}) : wire497);
              reg624 = $signed((reg466 ?
                  reg588 : {$signed((~&reg573)),
                      $unsigned(((8'hae) ? reg547 : reg448))}));
              reg625 = reg489;
            end
          if (reg449[(4'h9):(3'h7)])
            begin
              reg626 = $unsigned($unsigned($unsigned(({reg554, reg466} ?
                  reg573 : {reg486, forvar622}))));
            end
          else
            begin
              reg626 = (($unsigned($unsigned((reg559 ?
                  (8'h9f) : reg591))) ^~ reg530) * ($unsigned($signed(reg624)) <= (8'hbd)));
            end
        end
    end
  assign wire627 = (-wire439[(4'hc):(1'h1)]);
  always
    @(posedge clk) begin
      reg628 <= $signed(reg453[(2'h2):(1'h1)]);
      for (forvar629 = (1'h0); (forvar629 < (2'h3)); forvar629 = (forvar629 + (1'h1)))
        begin
          if (reg591[(4'hb):(4'h8)])
            begin
              reg630 = {$signed(reg601[(1'h1):(1'h1)]),
                  $signed($unsigned({$signed(reg502), reg561[(1'h0):(1'h0)]}))};
            end
          else
            begin
              reg631 <= $signed($unsigned(reg569[(4'h9):(1'h0)]));
            end
          if (wire438)
            begin
              reg632 = (reg588[(2'h2):(1'h1)] <= reg459[(1'h0):(1'h0)]);
              reg633 = $signed((8'hb3));
              reg634 <= (+(7'h4a));
              reg635 = $unsigned((|(|{$unsigned(reg541), $unsigned(reg552)})));
            end
          else
            begin
              reg634 <= (~&(^~((&$unsigned(reg466)) >= reg453[(1'h1):(1'h0)])));
              reg636 <= ($unsigned((reg634 ?
                      reg565[(4'hb):(2'h3)] : {reg633[(5'h13):(4'hb)]})) ?
                  (wire521 ? reg609 : reg461) : (-$signed(reg632)));
            end
        end
      reg637 = reg577[(1'h0):(1'h0)];
      if ((((((~wire436) - (reg448 & reg552)) + $signed(wire437)) ?
          (~&$unsigned((reg449 ? reg502 : reg549))) : reg541) < reg580))
        begin
          reg638 = (-{$unsigned($unsigned(((8'hbe) ? wire438 : (8'hbd)))),
              (-{$signed(reg632)})});
          reg639 = ($signed(reg489) > reg484[(3'h6):(2'h2)]);
          for (forvar640 = (1'h0); (forvar640 < (3'h4)); forvar640 = (forvar640 + (1'h1)))
            begin
              reg641 = $signed($signed({reg541[(3'h5):(3'h4)]}));
              reg642 = $signed(forvar640[(4'he):(3'h7)]);
              reg643 <= $signed({reg596});
            end
          for (forvar644 = (1'h0); (forvar644 < (3'h4)); forvar644 = (forvar644 + (1'h1)))
            begin
              reg645 = wire498[(3'h7):(3'h7)];
              reg646 <= $unsigned($unsigned((reg453 >>> ($signed(reg632) < (reg633 != reg461)))));
            end
          for (forvar647 = (1'h0); (forvar647 < (1'h0)); forvar647 = (forvar647 + (1'h1)))
            begin
              reg648 = reg577[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg640 <= reg532[(4'ha):(4'h9)];
          reg641 = $unsigned(wire498);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module266  (y, clk, wire271, wire270, wire269, wire268, wire267);
  output wire [(32'h7ef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h16):(1'h0)] wire271;
  input wire [(5'h13):(1'h0)] wire270;
  input wire signed [(4'h9):(1'h0)] wire269;
  input wire [(2'h2):(1'h0)] wire268;
  input wire signed [(4'hd):(1'h0)] wire267;
  wire [(5'h10):(1'h0)] wire430;
  wire [(4'h8):(1'h0)] wire338;
  wire [(5'h15):(1'h0)] wire337;
  wire signed [(5'h17):(1'h0)] wire336;
  wire [(4'hf):(1'h0)] wire335;
  wire [(3'h7):(1'h0)] wire334;
  wire signed [(5'h15):(1'h0)] wire333;
  wire signed [(3'h4):(1'h0)] wire332;
  reg signed [(2'h3):(1'h0)] reg429 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg426 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg425 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg423 = (1'h0);
  reg signed [(4'he):(1'h0)] reg421 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg420 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg419 = (1'h0);
  reg [(3'h6):(1'h0)] reg418 = (1'h0);
  reg signed [(4'he):(1'h0)] reg414 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg412 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg411 = (1'h0);
  reg [(2'h3):(1'h0)] reg410 = (1'h0);
  reg [(2'h3):(1'h0)] reg407 = (1'h0);
  reg [(5'h13):(1'h0)] reg406 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg404 = (1'h0);
  reg [(5'h15):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg402 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg398 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg397 = (1'h0);
  reg [(4'hd):(1'h0)] reg394 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg392 = (1'h0);
  reg [(5'h12):(1'h0)] reg391 = (1'h0);
  reg [(4'hd):(1'h0)] reg388 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg385 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg383 = (1'h0);
  reg [(4'h9):(1'h0)] reg382 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg380 = (1'h0);
  reg [(5'h12):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg378 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg377 = (1'h0);
  reg [(5'h14):(1'h0)] reg376 = (1'h0);
  reg [(3'h7):(1'h0)] reg375 = (1'h0);
  reg [(5'h14):(1'h0)] reg369 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg368 = (1'h0);
  reg [(4'h8):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg365 = (1'h0);
  reg [(5'h15):(1'h0)] reg364 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg363 = (1'h0);
  reg [(4'ha):(1'h0)] reg362 = (1'h0);
  reg [(5'h17):(1'h0)] reg361 = (1'h0);
  reg [(4'he):(1'h0)] reg359 = (1'h0);
  reg [(5'h16):(1'h0)] reg357 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg356 = (1'h0);
  reg [(2'h3):(1'h0)] reg355 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg352 = (1'h0);
  reg [(4'he):(1'h0)] reg351 = (1'h0);
  reg [(4'ha):(1'h0)] reg349 = (1'h0);
  reg [(3'h5):(1'h0)] reg348 = (1'h0);
  reg [(2'h2):(1'h0)] reg346 = (1'h0);
  reg [(4'hd):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg341 = (1'h0);
  reg [(3'h4):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg326 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg320 = (1'h0);
  reg [(5'h18):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg315 = (1'h0);
  reg [(3'h7):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg311 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg310 = (1'h0);
  reg [(3'h4):(1'h0)] reg309 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg306 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg305 = (1'h0);
  reg [(3'h4):(1'h0)] reg303 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg302 = (1'h0);
  reg [(4'hc):(1'h0)] reg301 = (1'h0);
  reg [(5'h12):(1'h0)] reg300 = (1'h0);
  reg [(3'h5):(1'h0)] reg299 = (1'h0);
  reg [(4'h9):(1'h0)] reg298 = (1'h0);
  reg [(5'h17):(1'h0)] reg295 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg294 = (1'h0);
  reg [(4'he):(1'h0)] reg293 = (1'h0);
  reg [(5'h15):(1'h0)] reg291 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg290 = (1'h0);
  reg [(4'h8):(1'h0)] reg289 = (1'h0);
  reg [(4'hb):(1'h0)] reg288 = (1'h0);
  reg [(5'h17):(1'h0)] reg287 = (1'h0);
  reg [(5'h10):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg282 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg280 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg279 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg276 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg275 = (1'h0);
  reg [(3'h4):(1'h0)] reg428 = (1'h0);
  reg [(3'h4):(1'h0)] reg427 = (1'h0);
  reg [(4'ha):(1'h0)] reg424 = (1'h0);
  reg [(3'h6):(1'h0)] forvar422 = (1'h0);
  reg [(5'h13):(1'h0)] reg417 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg415 = (1'h0);
  reg [(5'h17):(1'h0)] reg413 = (1'h0);
  reg [(5'h11):(1'h0)] forvar409 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg408 = (1'h0);
  reg [(4'h9):(1'h0)] reg405 = (1'h0);
  reg [(4'h9):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg400 = (1'h0);
  reg [(5'h12):(1'h0)] forvar399 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar396 = (1'h0);
  reg [(5'h17):(1'h0)] reg395 = (1'h0);
  reg [(4'hb):(1'h0)] reg393 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg390 = (1'h0);
  reg [(3'h6):(1'h0)] reg389 = (1'h0);
  reg [(5'h10):(1'h0)] reg387 = (1'h0);
  reg [(3'h7):(1'h0)] forvar386 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg384 = (1'h0);
  reg [(5'h11):(1'h0)] forvar372 = (1'h0);
  reg [(5'h17):(1'h0)] forvar359 = (1'h0);
  reg [(4'h9):(1'h0)] reg381 = (1'h0);
  reg [(5'h15):(1'h0)] reg374 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg373 = (1'h0);
  reg [(2'h2):(1'h0)] reg372 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg371 = (1'h0);
  reg [(4'h9):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg366 = (1'h0);
  reg [(4'hc):(1'h0)] reg360 = (1'h0);
  reg [(5'h14):(1'h0)] reg358 = (1'h0);
  reg [(3'h4):(1'h0)] reg354 = (1'h0);
  reg [(2'h2):(1'h0)] reg353 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg350 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg347 = (1'h0);
  reg [(5'h10):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg343 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar342 = (1'h0);
  reg [(5'h10):(1'h0)] forvar340 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg339 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg331 = (1'h0);
  reg signed [(4'he):(1'h0)] reg330 = (1'h0);
  reg [(4'ha):(1'h0)] reg329 = (1'h0);
  reg [(4'hc):(1'h0)] forvar327 = (1'h0);
  reg [(5'h16):(1'h0)] reg325 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg324 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar322 = (1'h0);
  reg [(5'h11):(1'h0)] reg321 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg319 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg317 = (1'h0);
  reg [(3'h4):(1'h0)] forvar316 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg313 = (1'h0);
  reg [(3'h4):(1'h0)] reg308 = (1'h0);
  reg [(3'h6):(1'h0)] reg307 = (1'h0);
  reg [(5'h16):(1'h0)] reg304 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg297 = (1'h0);
  reg [(5'h16):(1'h0)] forvar296 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar292 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar286 = (1'h0);
  reg [(4'hd):(1'h0)] reg285 = (1'h0);
  reg [(2'h3):(1'h0)] reg284 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar281 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg277 = (1'h0);
  reg signed [(4'he):(1'h0)] reg274 = (1'h0);
  reg [(3'h7):(1'h0)] forvar273 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg272 = (1'h0);
  assign y = {wire430,
                 wire338,
                 wire337,
                 wire336,
                 wire335,
                 wire334,
                 wire333,
                 wire332,
                 reg429,
                 reg426,
                 reg425,
                 reg423,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg414,
                 reg412,
                 reg411,
                 reg410,
                 reg407,
                 reg406,
                 reg404,
                 reg403,
                 reg402,
                 reg398,
                 reg397,
                 reg394,
                 reg392,
                 reg391,
                 reg388,
                 reg385,
                 reg383,
                 reg382,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg369,
                 reg368,
                 reg367,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg359,
                 reg357,
                 reg356,
                 reg355,
                 reg352,
                 reg351,
                 reg349,
                 reg348,
                 reg346,
                 reg345,
                 reg341,
                 reg328,
                 reg326,
                 reg323,
                 reg320,
                 reg318,
                 reg315,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg306,
                 reg305,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg295,
                 reg294,
                 reg293,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg283,
                 reg282,
                 reg280,
                 reg279,
                 reg278,
                 reg276,
                 reg275,
                 reg428,
                 reg427,
                 reg424,
                 forvar422,
                 reg417,
                 reg416,
                 reg415,
                 reg413,
                 forvar409,
                 reg408,
                 reg405,
                 reg401,
                 reg400,
                 forvar399,
                 forvar396,
                 reg395,
                 reg393,
                 reg390,
                 reg389,
                 reg387,
                 forvar386,
                 reg384,
                 forvar372,
                 forvar359,
                 reg381,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg366,
                 reg360,
                 reg358,
                 reg354,
                 reg353,
                 reg350,
                 reg347,
                 reg344,
                 reg343,
                 forvar342,
                 forvar340,
                 reg339,
                 reg331,
                 reg330,
                 reg329,
                 forvar327,
                 reg325,
                 reg324,
                 forvar322,
                 reg321,
                 reg319,
                 reg317,
                 forvar316,
                 reg314,
                 reg313,
                 reg308,
                 reg307,
                 reg304,
                 reg297,
                 forvar296,
                 forvar292,
                 forvar286,
                 reg285,
                 reg284,
                 forvar281,
                 reg277,
                 reg274,
                 forvar273,
                 reg272,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg272 = (wire271 * $unsigned($signed((wire268 ?
          (8'ha9) : wire270[(5'h10):(4'hd)]))));
      for (forvar273 = (1'h0); (forvar273 < (1'h1)); forvar273 = (forvar273 + (1'h1)))
        begin
          reg274 = forvar273;
          if (reg272[(5'h18):(5'h14)])
            begin
              reg275 <= $unsigned({((~|$signed((8'h9f))) ?
                      (~&$signed(wire269)) : $unsigned(reg272[(1'h1):(1'h1)])),
                  {wire269}});
              reg276 <= $signed(($signed($unsigned(wire268)) ?
                  forvar273[(2'h2):(1'h1)] : (($signed(wire269) ^~ wire267) ?
                      (wire271[(4'hd):(1'h1)] ?
                          $unsigned(wire270) : (wire270 | reg272)) : ((reg274 == reg272) ?
                          reg272 : (|wire267)))));
            end
          else
            begin
              reg277 = reg272;
              reg278 <= reg276[(1'h1):(1'h0)];
              reg279 <= $signed($unsigned((8'hbe)));
              reg280 <= (wire269 ?
                  reg276 : ({{$signed(reg277)}, reg274} < (+(^(-reg275)))));
            end
          for (forvar281 = (1'h0); (forvar281 < (1'h0)); forvar281 = (forvar281 + (1'h1)))
            begin
              reg282 <= reg275[(1'h0):(1'h0)];
              reg283 <= reg277[(4'h8):(2'h2)];
              reg284 = (~|(reg283 ?
                  (|(wire267[(3'h4):(3'h4)] ^ (reg278 ?
                      forvar281 : (8'hb9)))) : reg275[(2'h3):(2'h2)]));
            end
        end
      if (((|((-$signed(wire271)) ?
          $unsigned((8'hac)) : reg283)) << ((wire269[(3'h6):(2'h2)] ?
          ((~forvar273) | (reg280 ?
              reg284 : (8'hbe))) : wire267[(4'hb):(4'h8)]) ^~ reg277)))
        begin
          reg285 = (&wire268);
        end
      else
        begin
          if (wire271)
            begin
              reg285 = {wire267[(4'ha):(1'h1)], reg282};
            end
          else
            begin
              reg285 = reg284[(1'h1):(1'h0)];
            end
          for (forvar286 = (1'h0); (forvar286 < (1'h1)); forvar286 = (forvar286 + (1'h1)))
            begin
              reg287 <= (~&($signed($unsigned(reg280[(3'h5):(1'h1)])) ?
                  $signed($signed($unsigned(reg277))) : (wire267 ?
                      $signed($unsigned(forvar281)) : reg274[(4'hd):(1'h0)])));
              reg288 <= $unsigned((reg280[(3'h4):(1'h0)] & reg284[(2'h2):(1'h1)]));
              reg289 <= $signed($unsigned($unsigned(reg272[(4'hc):(2'h2)])));
              reg290 <= (^{$unsigned({wire269[(3'h4):(2'h3)],
                      $signed(reg278)})});
              reg291 <= $signed(reg283);
            end
          for (forvar292 = (1'h0); (forvar292 < (1'h0)); forvar292 = (forvar292 + (1'h1)))
            begin
              reg293 <= $signed(($unsigned(($unsigned((8'ha5)) || $unsigned(reg280))) ?
                  wire271[(4'ha):(3'h6)] : $signed(reg275[(3'h5):(1'h0)])));
              reg294 <= $unsigned((reg291[(3'h7):(2'h2)] ^~ (8'hba)));
              reg295 <= ((!(reg275 ? $signed(wire268) : $unsigned(wire268))) ?
                  (($signed($unsigned(forvar286)) ?
                          ((forvar292 ? reg282 : forvar281) >= (reg287 ?
                              forvar292 : reg294)) : (forvar281[(4'hb):(3'h5)] != $signed(reg280))) ?
                      reg274[(1'h0):(1'h0)] : reg275) : reg291);
            end
        end
      for (forvar296 = (1'h0); (forvar296 < (3'h4)); forvar296 = (forvar296 + (1'h1)))
        begin
          reg297 = {(!$signed(reg282[(4'ha):(4'h9)])), {reg277[(1'h0):(1'h0)]}};
          reg298 <= ((reg279 * wire270[(1'h1):(1'h1)]) ?
              reg275 : (reg284[(1'h1):(1'h0)] && $signed(((~|wire271) ^~ (reg295 <= (8'hba))))));
          if ((wire267[(4'hd):(4'ha)] << $unsigned($unsigned(({wire268} ?
              $signed(reg297) : (reg293 ~^ (8'hbd)))))))
            begin
              reg299 <= (reg288[(2'h3):(1'h0)] - reg284[(2'h3):(1'h0)]);
              reg300 <= reg298[(2'h3):(1'h1)];
            end
          else
            begin
              reg299 <= (&wire269[(3'h4):(1'h1)]);
              reg300 <= reg272[(4'h8):(3'h4)];
              reg301 <= reg285[(3'h6):(2'h3)];
              reg302 <= reg284;
            end
          if (forvar296)
            begin
              reg303 <= $unsigned($unsigned(($signed((wire270 ?
                      forvar281 : reg295)) ?
                  reg293 : $signed((reg288 ? (8'hbc) : (8'ha7))))));
            end
          else
            begin
              reg304 = ($signed($signed(forvar296[(3'h6):(1'h0)])) ?
                  (&$signed(reg290[(1'h1):(1'h1)])) : $unsigned($signed((forvar286[(3'h5):(3'h5)] ?
                      (reg291 >>> wire268) : $signed(forvar281)))));
              reg305 <= reg279;
              reg306 <= $signed(wire268);
            end
          if ($signed(reg306[(3'h7):(1'h0)]))
            begin
              reg307 = ((8'h9f) >= ($signed(reg306[(3'h6):(3'h5)]) > (($signed(forvar273) - $signed(reg295)) - (reg277[(3'h6):(1'h1)] == wire270))));
              reg308 = reg304;
            end
          else
            begin
              reg309 <= (&reg308);
              reg310 <= (((reg277 == $unsigned($unsigned(forvar286))) ?
                  (wire270 > $unsigned((reg307 && reg308))) : (8'hab)) && (~|$unsigned((wire271[(4'hc):(3'h4)] == $signed(reg294)))));
              reg311 <= $signed(({reg293[(4'ha):(2'h3)],
                  reg287[(4'hd):(4'hb)]} + ((&(^wire269)) ?
                  (reg297[(2'h2):(2'h2)] != (~^(8'hb5))) : {(wire267 ~^ reg300)})));
              reg312 <= (8'h9e);
            end
        end
      if ({$signed(reg302)})
        begin
          reg313 = $unsigned(reg311[(5'h11):(5'h11)]);
          reg314 = ($unsigned({(wire271[(3'h6):(1'h1)] ?
                  (wire267 ?
                      reg291 : (8'hb7)) : $unsigned(reg293))}) + $signed(((forvar286[(3'h7):(2'h2)] ?
                  (reg291 - forvar286) : reg289[(1'h1):(1'h0)]) ?
              reg308 : ((forvar292 ? reg293 : reg308) - $unsigned((7'h48))))));
          reg315 <= reg312;
          for (forvar316 = (1'h0); (forvar316 < (2'h2)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg317 = reg294[(3'h7):(3'h4)];
              reg318 <= reg309[(2'h2):(1'h0)];
              reg319 = (8'hbb);
            end
          reg320 <= (^~(({reg319} ?
              (reg279 != reg279[(3'h6):(3'h4)]) : {(reg304 << (7'h48)),
                  ((8'hb6) >>> wire269)}) ~^ reg306[(3'h4):(2'h3)]));
        end
      else
        begin
          reg315 <= (reg279[(3'h5):(2'h2)] ?
              (~^(^~$unsigned((reg283 < forvar281)))) : reg302);
          for (forvar316 = (1'h0); (forvar316 < (1'h0)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg318 <= (|$signed(($signed(reg315[(5'h13):(5'h11)]) - $unsigned({reg284,
                  (8'hbc)}))));
              reg320 <= ($signed(($unsigned((reg277 - forvar292)) > forvar286)) | $unsigned(($signed(reg293[(3'h5):(3'h4)]) ?
                  (reg284[(2'h2):(1'h1)] ?
                      $unsigned(reg287) : (reg300 ?
                          reg303 : (8'hb9))) : reg302[(1'h0):(1'h0)])));
              reg321 = (|($unsigned($signed((|reg311))) ?
                  (reg308 ?
                      ((reg294 >>> forvar292) != $unsigned(reg312)) : ((^~reg306) ?
                          reg301[(4'hc):(4'hc)] : $unsigned(reg318))) : {((reg276 ^~ reg278) ?
                          (+reg317) : wire267),
                      $unsigned((reg302 == reg277))}));
            end
          for (forvar322 = (1'h0); (forvar322 < (2'h2)); forvar322 = (forvar322 + (1'h1)))
            begin
              reg323 <= forvar322;
              reg324 = {{forvar322[(3'h4):(1'h1)]},
                  $unsigned((^$unsigned(reg282[(2'h3):(2'h2)])))};
              reg325 = {$unsigned($signed(((8'h9c) ? wire268 : (~(8'hba)))))};
            end
          reg326 <= $signed($signed(reg319));
          for (forvar327 = (1'h0); (forvar327 < (1'h0)); forvar327 = (forvar327 + (1'h1)))
            begin
              reg328 <= (8'hb6);
              reg329 = (~&$unsigned(reg323[(3'h4):(2'h3)]));
              reg330 = ((((^$signed(reg305)) ?
                  $unsigned({reg326}) : ($unsigned(reg301) ^~ (forvar316 ?
                      forvar281 : reg325))) != reg329) != (^reg289[(3'h7):(3'h7)]));
              reg331 = (^(^~($unsigned($unsigned(forvar316)) ?
                  $signed((reg274 <<< reg313)) : $signed((reg328 ?
                      reg312 : (8'hb1))))));
            end
        end
    end
  assign wire332 = reg291;
  assign wire333 = (^~reg276[(1'h1):(1'h1)]);
  assign wire334 = (reg320 ^~ ((~|(~^(wire332 != reg279))) && reg290));
  assign wire335 = (((reg287 ~^ $signed((reg323 ?
                           reg318 : wire268))) < (($signed(reg298) ?
                               reg310 : wire268) ?
                           ((reg299 == wire270) ^ reg282) : ($signed(reg288) ?
                               reg311[(4'hc):(1'h0)] : (reg288 ?
                                   reg301 : wire269)))) ?
                       (^~reg291[(1'h0):(1'h0)]) : reg311);
  assign wire336 = reg309[(3'h4):(3'h4)];
  assign wire337 = $unsigned($unsigned((|$signed($unsigned(wire270)))));
  assign wire338 = $unsigned($signed(((reg299[(2'h2):(2'h2)] > {reg302}) ?
                       (!(~reg309)) : reg283[(4'he):(3'h4)])));
  always
    @(posedge clk) begin
      reg339 = $unsigned((reg315[(3'h6):(3'h6)] << (+$signed((reg275 ?
          reg293 : reg295)))));
      for (forvar340 = (1'h0); (forvar340 < (2'h3)); forvar340 = (forvar340 + (1'h1)))
        begin
          reg341 <= (reg278[(2'h2):(2'h2)] ?
              $unsigned((&(^(8'ha1)))) : $unsigned(reg328[(2'h3):(2'h2)]));
          for (forvar342 = (1'h0); (forvar342 < (2'h3)); forvar342 = (forvar342 + (1'h1)))
            begin
              reg343 = ((reg306 ?
                  $signed(({reg301} ~^ {(8'hb6)})) : ($signed((-reg294)) ?
                      $unsigned((reg300 ?
                          reg276 : (8'ha8))) : ($unsigned(reg305) || $unsigned(reg275)))) >> reg315[(4'hb):(1'h1)]);
              reg344 = (~(reg343[(4'hd):(3'h4)] >= reg343));
              reg345 <= (+reg302);
              reg346 <= ($signed({{reg341[(5'h18):(2'h3)], {reg301}}}) ?
                  reg301[(2'h2):(1'h1)] : (+$signed((((8'h9d) != reg280) < (wire333 ?
                      reg290 : reg344)))));
              reg347 = (($signed(wire270) <<< $signed(reg326[(3'h5):(2'h2)])) >>> reg346[(1'h0):(1'h0)]);
            end
          if ($unsigned($signed($signed(reg289[(3'h6):(2'h2)]))))
            begin
              reg348 <= reg291;
              reg349 <= (8'hbd);
              reg350 = {($unsigned((forvar340[(4'hd):(4'h9)] ?
                      $signed((8'ha5)) : wire336)) + reg309[(3'h4):(2'h2)]),
                  $unsigned($signed((8'ha6)))};
              reg351 <= $unsigned(reg287);
            end
          else
            begin
              reg348 <= {({$unsigned((wire334 <= reg341))} ?
                      $unsigned(reg311) : {(+reg299),
                          $signed({wire271, (8'ha9)})})};
            end
          reg352 <= $signed((~|reg349));
          if ($unsigned((-(~&($signed(reg288) ?
              (reg343 <<< wire338) : {reg347, (7'h47)})))))
            begin
              reg353 = reg323[(2'h3):(2'h3)];
              reg354 = reg293[(1'h0):(1'h0)];
              reg355 <= wire333[(3'h6):(3'h6)];
              reg356 <= reg328;
              reg357 <= reg310[(3'h5):(2'h2)];
            end
          else
            begin
              reg353 = $signed(reg315[(5'h12):(2'h2)]);
              reg354 = ((~&($unsigned($unsigned(reg300)) ?
                      {reg290, (reg278 && reg294)} : {(!reg310), reg349})) ?
                  $unsigned((8'h9c)) : {((8'hbb) != reg298)});
              reg358 = $unsigned((wire270[(3'h4):(1'h1)] >> wire335[(4'hd):(2'h2)]));
            end
        end
      if (reg356)
        begin
          reg359 <= $signed(reg302);
          if ($unsigned((((-(reg349 ~^ reg299)) ?
              $signed(wire334) : (^$unsigned(reg347))) * $signed((reg345 ^~ (reg280 ?
              reg303 : reg289))))))
            begin
              reg360 = (~(^((reg355 ? $signed(reg350) : ((8'hbe) + reg345)) ?
                  (+reg291) : reg354[(2'h2):(1'h0)])));
            end
          else
            begin
              reg361 <= $unsigned(reg291[(4'ha):(3'h5)]);
              reg362 <= {reg355};
            end
          if ($unsigned($unsigned((~|((8'hb0) ?
              (reg320 ? wire271 : reg350) : {wire335})))))
            begin
              reg363 <= $unsigned(((~($signed(reg280) ?
                  $unsigned(reg291) : (reg293 ?
                      reg344 : wire334))) ^ reg345[(4'hb):(4'ha)]));
              reg364 <= $unsigned((~^wire271[(3'h5):(3'h5)]));
              reg365 <= wire337;
            end
          else
            begin
              reg366 = $unsigned(($unsigned((reg305 ?
                  $signed(reg289) : $signed(reg365))) - {$signed($signed(reg300)),
                  reg361[(4'h8):(3'h4)]}));
              reg367 <= ($signed(((^(8'hb0)) >> reg341[(4'hd):(4'hb)])) >>> reg341[(3'h4):(1'h1)]);
              reg368 <= (7'h45);
              reg369 <= (reg365 ?
                  ($unsigned(reg289[(1'h1):(1'h1)]) * $unsigned($signed($signed(reg301)))) : $unsigned($signed((!reg306))));
            end
          if ((wire337 >>> $unsigned((8'hbf))))
            begin
              reg370 = ($signed((~$signed(reg283[(4'hd):(4'hd)]))) ?
                  {(^~(|reg366[(1'h0):(1'h0)])),
                      {(!(reg293 + forvar340)),
                          $unsigned($unsigned(reg346))}} : reg362[(4'ha):(4'h8)]);
              reg371 = ((-reg345) >= reg295);
              reg372 = (($signed($unsigned($signed(reg364))) ?
                      reg371 : reg359[(4'h8):(3'h5)]) ?
                  (wire332[(2'h3):(1'h0)] * reg349) : reg289);
              reg373 = ($unsigned((-(|(reg359 ?
                  (8'h9c) : (8'hbd))))) ^ (8'hba));
              reg374 = reg326;
            end
          else
            begin
              reg375 <= ($signed($unsigned((8'hb6))) | $unsigned(wire271[(4'ha):(3'h4)]));
              reg376 <= (8'ha6);
              reg377 <= (((reg294[(3'h6):(3'h4)] && (~|reg371)) ?
                  wire335[(4'hd):(2'h2)] : reg355[(1'h1):(1'h0)]) != $unsigned($unsigned($signed((&(7'h49))))));
            end
          if ({wire268[(2'h2):(2'h2)]})
            begin
              reg378 <= (((($unsigned(reg301) ? (8'hb7) : $signed(reg361)) ?
                      reg295[(5'h11):(3'h6)] : {forvar340[(3'h7):(2'h2)],
                          $unsigned(reg357)}) ~^ reg300[(3'h6):(2'h3)]) ?
                  $signed(((reg339[(4'h9):(3'h7)] <= $signed((8'h9e))) ?
                      reg364[(3'h5):(2'h3)] : {{reg351, reg361},
                          reg288})) : $unsigned(($unsigned(((8'ha0) ?
                          (7'h49) : wire270)) ?
                      ({reg278, reg276} ?
                          reg278[(3'h4):(2'h3)] : (~^(7'h42))) : (-(reg275 && reg377)))));
              reg379 <= ({{((+reg359) < (reg378 == reg355)),
                          $unsigned((&reg362))},
                      reg311} ?
                  (^~(~^($unsigned(reg378) ?
                      reg364[(4'hd):(3'h4)] : (reg310 ?
                          reg315 : (8'ha6))))) : ($unsigned($unsigned(reg368[(4'h8):(3'h6)])) + $unsigned(($unsigned(reg300) >= reg298[(3'h4):(2'h3)]))));
              reg380 <= (($signed($unsigned(reg343[(4'ha):(3'h4)])) ?
                      (((reg358 ? reg366 : reg358) & reg300[(5'h11):(5'h11)]) ?
                          ((&reg354) + (wire338 ?
                              reg375 : (8'hae))) : {$signed(wire267)}) : ({(reg377 ?
                                  wire336 : (8'ha9)),
                              (^reg320)} ?
                          ({reg349} ?
                              (~&reg275) : (wire270 == wire267)) : (~&wire269[(3'h5):(1'h1)]))) ?
                  (~{$unsigned(((8'hb0) ? wire337 : reg312)),
                      ((8'ha4) ^~ reg279)}) : (reg377[(2'h3):(2'h2)] ?
                      $signed((+(8'hab))) : ($signed($signed(reg374)) >= $unsigned($unsigned(reg290)))));
            end
          else
            begin
              reg381 = reg339[(4'hd):(2'h2)];
              reg382 <= reg348;
              reg383 <= {$unsigned(((+reg306) ?
                      $signed((8'hb7)) : $signed(wire337))),
                  (&((~&reg354) < $signed((~|reg301))))};
            end
        end
      else
        begin
          for (forvar359 = (1'h0); (forvar359 < (1'h0)); forvar359 = (forvar359 + (1'h1)))
            begin
              reg361 <= $signed($signed(((^~$unsigned(reg377)) || {$unsigned(forvar342),
                  $unsigned(reg372)})));
              reg366 = $unsigned({$signed((^~(reg339 ? reg328 : reg377))),
                  $unsigned($signed($signed(reg290)))});
              reg367 <= reg339[(5'h16):(1'h0)];
              reg370 = reg345;
              reg371 = $unsigned(wire334);
            end
          for (forvar372 = (1'h0); (forvar372 < (1'h0)); forvar372 = (forvar372 + (1'h1)))
            begin
              reg373 = $signed(reg326[(5'h17):(4'ha)]);
              reg374 = $signed(((+((~&(8'ha2)) ?
                  forvar342 : reg372)) < wire338));
            end
          reg381 = wire333[(5'h12):(1'h0)];
        end
      if (reg287[(1'h1):(1'h0)])
        begin
          reg384 = reg360[(2'h2):(1'h0)];
          reg385 <= (^~((reg370[(1'h1):(1'h0)] ?
              (reg379[(4'he):(3'h4)] ?
                  (~^wire271) : (reg350 * wire334)) : reg310[(3'h6):(2'h2)]) >> reg306[(3'h5):(3'h4)]));
          for (forvar386 = (1'h0); (forvar386 < (2'h2)); forvar386 = (forvar386 + (1'h1)))
            begin
              reg387 = $signed((~(8'ha9)));
              reg388 <= (({$signed((~(7'h44)))} >= {(8'h9d)}) ?
                  (reg318 ? reg289 : $unsigned(forvar359)) : wire337);
            end
          if ((($unsigned($unsigned(reg357)) != (($unsigned(reg283) <<< (|reg276)) ?
              ((|reg294) ^~ (&forvar340)) : $unsigned($unsigned(reg381)))) == $signed($unsigned((7'h44)))))
            begin
              reg389 = $signed({$signed($unsigned(reg375[(2'h2):(1'h1)])),
                  $unsigned($unsigned($unsigned(reg351)))});
              reg390 = (8'hbc);
            end
          else
            begin
              reg391 <= $unsigned(reg345[(1'h0):(1'h0)]);
              reg392 <= (((((~&reg364) | $unsigned(reg361)) != (~|$unsigned(reg299))) ?
                      $signed($unsigned({forvar386,
                          reg344})) : reg390[(4'hb):(3'h5)]) ?
                  $signed((~|forvar386)) : ({(reg344[(5'h10):(4'h8)] && $signed(reg381))} ?
                      (~|({reg379, reg383} ?
                          $signed((8'had)) : (reg389 << reg339))) : (forvar372[(4'hb):(1'h0)] && (8'h9c))));
              reg393 = reg283[(4'hd):(2'h3)];
              reg394 <= (-$unsigned((~^reg326[(3'h4):(3'h4)])));
            end
        end
      else
        begin
          reg385 <= reg291;
        end
      reg395 = reg368;
    end
  always
    @(posedge clk) begin
      for (forvar396 = (1'h0); (forvar396 < (2'h3)); forvar396 = (forvar396 + (1'h1)))
        begin
          reg397 <= wire334;
          reg398 <= (wire333[(3'h4):(2'h2)] ?
              reg323[(2'h2):(2'h2)] : (+(|reg315)));
        end
      if ({{(~^$signed($signed(reg368))), reg383[(4'h9):(2'h3)]}, reg305})
        begin
          for (forvar399 = (1'h0); (forvar399 < (2'h2)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg400 = ($unsigned(((reg378 ?
                      {wire335} : reg295[(5'h17):(4'hb)]) >>> $unsigned(reg294[(3'h4):(3'h4)]))) ?
                  $signed($signed(reg369[(5'h14):(1'h0)])) : reg298[(3'h6):(3'h6)]);
              reg401 = $unsigned(wire269);
              reg402 <= reg345;
            end
          reg403 <= {$signed($unsigned(({reg355} ^ (^reg364))))};
          reg404 <= (~|reg378);
        end
      else
        begin
          for (forvar399 = (1'h0); (forvar399 < (3'h4)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg402 <= (({$signed((~(8'ha2)))} <= {wire333,
                  $unsigned(reg388[(4'hb):(2'h2)])}) == (7'h40));
              reg403 <= reg404[(1'h0):(1'h0)];
              reg405 = reg397[(1'h1):(1'h0)];
              reg406 <= ((~&$unsigned(reg312[(1'h1):(1'h0)])) <<< (^((reg326 ~^ reg289) <= (+(forvar396 ?
                  reg351 : reg283)))));
            end
          reg407 <= (reg359 ?
              (((~&(-reg341)) < reg280) ?
                  $unsigned((reg294[(3'h6):(3'h5)] ^ reg375)) : wire271) : reg388[(1'h1):(1'h1)]);
          reg408 = $signed(wire270);
        end
      for (forvar409 = (1'h0); (forvar409 < (2'h3)); forvar409 = (forvar409 + (1'h1)))
        begin
          if (((8'hae) ?
              (^~($signed($unsigned(reg306)) ?
                  reg378[(4'hc):(4'h8)] : wire333[(5'h12):(2'h2)])) : wire336[(5'h14):(2'h3)]))
            begin
              reg410 <= $signed($unsigned($signed(($unsigned(reg408) ?
                  {reg276, reg356} : reg293))));
              reg411 <= $signed({((reg391[(2'h2):(1'h0)] ?
                      $unsigned(forvar409) : $signed(reg404)) == reg382[(4'h9):(3'h7)])});
              reg412 <= ((!(8'hb8)) ?
                  (reg385[(1'h1):(1'h1)] << reg356[(2'h3):(1'h1)]) : ((reg410 ?
                      (-$signed(reg363)) : reg310[(3'h4):(1'h0)]) | $signed(reg288[(3'h7):(3'h5)])));
              reg413 = {$signed(reg365), (&(!{reg364}))};
              reg414 <= reg318;
            end
          else
            begin
              reg410 <= {reg288[(4'hb):(2'h2)],
                  (^(((~&reg291) * (+(8'ha8))) ?
                      (reg311 ?
                          $signed(reg341) : reg346[(2'h2):(2'h2)]) : ((reg402 >>> wire336) >= (reg357 ?
                          reg315 : reg364))))};
              reg413 = reg383[(2'h3):(2'h3)];
              reg415 = $unsigned((reg378[(3'h7):(1'h1)] ?
                  reg326 : $unsigned($signed($signed(reg368)))));
              reg416 = reg352;
            end
          if ((($unsigned((8'hb6)) << ((reg290[(2'h2):(2'h2)] ?
                  $signed(wire333) : $unsigned(reg311)) + ((8'hbf) | (reg388 ?
                  reg302 : reg355)))) ?
              (($signed($signed((8'h9d))) ^~ $unsigned((reg377 ?
                  reg406 : (7'h47)))) || $unsigned(reg415[(5'h15):(4'hd)])) : $unsigned(reg398)))
            begin
              reg417 = (~^$unsigned($signed({reg315[(5'h10):(4'hc)]})));
              reg418 <= reg299[(1'h1):(1'h0)];
              reg419 <= reg378;
              reg420 <= $signed(($unsigned((^reg361)) ~^ reg352));
              reg421 <= reg385;
            end
          else
            begin
              reg418 <= reg287;
            end
        end
      for (forvar422 = (1'h0); (forvar422 < (1'h0)); forvar422 = (forvar422 + (1'h1)))
        begin
          reg423 <= reg412[(2'h2):(2'h2)];
          if (($unsigned(({(wire332 ?
                      reg394 : reg309)} <<< reg383[(2'h3):(1'h1)])) ?
              $unsigned((+reg289[(3'h7):(2'h3)])) : (reg359 ?
                  (^~reg368) : (-wire338[(1'h0):(1'h0)]))))
            begin
              reg424 = (|$signed(reg362));
            end
          else
            begin
              reg424 = $unsigned(((((reg295 >= reg278) ?
                  wire337[(3'h4):(1'h0)] : $signed(reg376)) & $unsigned(((8'hbb) <= reg311))) - (+$signed((~reg295)))));
              reg425 <= reg410[(2'h2):(1'h0)];
              reg426 <= (^(&(|$signed($unsigned(wire269)))));
              reg427 = (^$signed($signed(($unsigned(reg375) ?
                  $unsigned(reg415) : (8'hb7)))));
            end
          reg428 = (!$signed({reg382, reg309}));
          reg429 <= {(reg356[(3'h6):(3'h4)] ? wire338 : reg359)};
        end
    end
  assign wire430 = (reg287 ?
                       $unsigned(((reg318 > wire332) >= reg282[(4'hb):(3'h4)])) : (reg318[(1'h0):(1'h0)] >= (~^((wire335 > reg287) ?
                           $unsigned(reg365) : (&reg380)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module127  (y, clk, wire132, wire131, wire130, wire129, wire128);
  output wire [(32'h413):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire132;
  input wire signed [(5'h16):(1'h0)] wire131;
  input wire [(5'h16):(1'h0)] wire130;
  input wire signed [(5'h11):(1'h0)] wire129;
  input wire signed [(5'h11):(1'h0)] wire128;
  wire [(3'h7):(1'h0)] wire204;
  wire signed [(4'hb):(1'h0)] wire179;
  wire [(2'h2):(1'h0)] wire178;
  wire [(2'h3):(1'h0)] wire177;
  wire [(5'h18):(1'h0)] wire176;
  wire [(3'h5):(1'h0)] wire133;
  reg [(5'h15):(1'h0)] reg213 = (1'h0);
  reg signed [(4'he):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg206 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg205 = (1'h0);
  reg [(5'h15):(1'h0)] reg203 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg202 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg201 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg189 = (1'h0);
  reg signed [(4'he):(1'h0)] reg183 = (1'h0);
  reg [(4'h8):(1'h0)] reg182 = (1'h0);
  reg [(4'h8):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg169 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg166 = (1'h0);
  reg [(4'h9):(1'h0)] reg165 = (1'h0);
  reg [(2'h2):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg162 = (1'h0);
  reg [(4'hd):(1'h0)] reg159 = (1'h0);
  reg [(3'h5):(1'h0)] reg158 = (1'h0);
  reg [(3'h6):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg156 = (1'h0);
  reg [(3'h5):(1'h0)] reg154 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg150 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg149 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg148 = (1'h0);
  reg [(3'h6):(1'h0)] reg147 = (1'h0);
  reg [(3'h5):(1'h0)] reg145 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg143 = (1'h0);
  reg [(5'h15):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg139 = (1'h0);
  reg [(3'h6):(1'h0)] reg138 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg137 = (1'h0);
  reg [(3'h4):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg215 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar214 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar211 = (1'h0);
  reg [(4'hb):(1'h0)] reg210 = (1'h0);
  reg [(2'h2):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg207 = (1'h0);
  reg [(4'hd):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar199 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg197 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg196 = (1'h0);
  reg [(5'h17):(1'h0)] reg195 = (1'h0);
  reg [(5'h14):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar192 = (1'h0);
  reg [(4'hf):(1'h0)] reg191 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar190 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg188 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg187 = (1'h0);
  reg [(5'h18):(1'h0)] forvar186 = (1'h0);
  reg [(2'h3):(1'h0)] reg185 = (1'h0);
  reg [(4'hd):(1'h0)] reg184 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar181 = (1'h0);
  reg [(4'h8):(1'h0)] forvar180 = (1'h0);
  reg [(4'he):(1'h0)] reg175 = (1'h0);
  reg [(5'h17):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg171 = (1'h0);
  reg [(5'h14):(1'h0)] reg170 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg168 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar163 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg161 = (1'h0);
  reg [(2'h2):(1'h0)] reg160 = (1'h0);
  reg [(4'hb):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg153 = (1'h0);
  reg [(3'h6):(1'h0)] forvar152 = (1'h0);
  reg [(3'h7):(1'h0)] forvar151 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar142 = (1'h0);
  reg [(4'he):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar135 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar134 = (1'h0);
  assign y = {wire204,
                 wire179,
                 wire178,
                 wire177,
                 wire176,
                 wire133,
                 reg213,
                 reg212,
                 reg208,
                 reg206,
                 reg205,
                 reg203,
                 reg202,
                 reg201,
                 reg198,
                 reg193,
                 reg189,
                 reg183,
                 reg182,
                 reg174,
                 reg172,
                 reg169,
                 reg166,
                 reg165,
                 reg164,
                 reg162,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg154,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg145,
                 reg143,
                 reg141,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg215,
                 forvar214,
                 forvar211,
                 reg210,
                 reg209,
                 reg207,
                 reg200,
                 forvar199,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 forvar192,
                 reg191,
                 forvar190,
                 reg188,
                 reg187,
                 forvar186,
                 reg185,
                 reg184,
                 forvar181,
                 forvar180,
                 reg175,
                 reg173,
                 reg171,
                 reg170,
                 reg168,
                 reg167,
                 forvar163,
                 reg161,
                 reg160,
                 reg155,
                 reg153,
                 forvar152,
                 forvar151,
                 reg146,
                 reg144,
                 forvar142,
                 reg140,
                 forvar135,
                 forvar134,
                 (1'h0)};
  assign wire133 = (wire128[(2'h3):(1'h1)] ^~ $unsigned(wire129[(3'h5):(3'h4)]));
  always
    @(posedge clk) begin
      for (forvar134 = (1'h0); (forvar134 < (2'h3)); forvar134 = (forvar134 + (1'h1)))
        begin
          for (forvar135 = (1'h0); (forvar135 < (2'h2)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= $unsigned({$signed((wire129 ?
                      $unsigned(wire130) : $unsigned(wire133)))});
              reg137 <= {((7'h40) ?
                      $unsigned(wire129[(3'h6):(1'h1)]) : ((^~$unsigned(wire133)) * (wire131 ?
                          reg136[(2'h3):(1'h1)] : (wire129 ?
                              wire132 : forvar135)))),
                  ($unsigned(wire129[(5'h11):(1'h0)]) >= {({forvar134,
                          forvar134} >>> {forvar134, wire133})})};
              reg138 <= $unsigned($signed(wire129[(4'hb):(2'h2)]));
              reg139 <= ($signed(wire128[(3'h6):(3'h6)]) ? wire129 : (8'hbd));
              reg140 = (+$signed($unsigned((reg139[(5'h11):(3'h7)] + {wire131}))));
            end
          reg141 <= $unsigned($signed((8'hb0)));
          for (forvar142 = (1'h0); (forvar142 < (1'h1)); forvar142 = (forvar142 + (1'h1)))
            begin
              reg143 <= ($signed((((~|(7'h44)) <<< wire131) ?
                  reg140[(1'h0):(1'h0)] : (!(wire129 ?
                      (8'hb6) : reg136)))) - {($signed(wire132[(3'h4):(1'h1)]) ?
                      $unsigned(wire130[(5'h10):(3'h7)]) : ({reg136, reg139} ?
                          wire130[(3'h5):(2'h3)] : (&reg139))),
                  wire131[(5'h11):(2'h2)]});
              reg144 = forvar135[(2'h2):(2'h2)];
            end
        end
      if ($signed((reg140[(2'h2):(1'h0)] ?
          ($signed(reg140) + ((^reg143) ?
              $unsigned((8'hb9)) : $unsigned(reg144))) : (forvar142[(2'h2):(1'h0)] ?
              reg140[(2'h2):(1'h1)] : $signed({reg143, (7'h42)})))))
        begin
          reg145 <= (|(wire128 == $signed(reg144[(5'h12):(3'h7)])));
        end
      else
        begin
          if ({(!(forvar142[(4'ha):(3'h6)] ?
                  reg141[(4'ha):(3'h7)] : (((7'h41) <<< wire130) ^~ (!reg144)))),
              $unsigned({(((8'ha4) ? wire132 : reg137) ?
                      (~^wire131) : $unsigned(forvar134))})})
            begin
              reg146 = (reg141[(3'h7):(1'h0)] ?
                  forvar142[(2'h3):(1'h0)] : reg138);
              reg147 <= {($unsigned((|wire130[(4'hd):(1'h1)])) ?
                      (((!(8'h9c)) ? $unsigned(forvar134) : (8'ha7)) ?
                          $unsigned($unsigned(reg139)) : ($unsigned(reg143) >> (~|reg139))) : reg139[(2'h2):(1'h0)]),
                  (reg141 ?
                      $unsigned($signed(forvar134)) : ({wire129,
                          reg146} <<< reg139))};
              reg148 <= $unsigned(wire129[(4'hc):(3'h6)]);
              reg149 <= (|($unsigned({reg144,
                  (forvar135 ? reg140 : (8'hb9))}) >= wire131));
              reg150 <= {((7'h44) ^~ (~|$signed((^reg141))))};
            end
          else
            begin
              reg146 = $signed({(^((8'ha9) ? $unsigned(reg139) : (+(8'h9f)))),
                  $signed((reg150[(1'h0):(1'h0)] >= reg146))});
            end
        end
      for (forvar151 = (1'h0); (forvar151 < (2'h3)); forvar151 = (forvar151 + (1'h1)))
        begin
          for (forvar152 = (1'h0); (forvar152 < (1'h0)); forvar152 = (forvar152 + (1'h1)))
            begin
              reg153 = (7'h42);
              reg154 <= ($unsigned({{$unsigned(reg141),
                      (~^(8'hb3))}}) - (($unsigned({forvar152,
                      reg147}) > ((^~(8'hbc)) | $unsigned(wire130))) ?
                  {{(reg148 || wire132)}} : forvar135));
              reg155 = (~$signed($unsigned(wire130)));
              reg156 <= reg154;
            end
          if ({wire131[(4'hf):(4'hb)]})
            begin
              reg157 <= $signed({reg155});
              reg158 <= {($signed($unsigned($signed(reg137))) ?
                      ((&forvar135[(3'h4):(2'h2)]) ^ (-$signed((8'ha5)))) : (reg140[(4'ha):(3'h7)] <= ($unsigned(forvar142) << reg154)))};
              reg159 <= $unsigned(($unsigned(((reg147 ?
                      reg154 : forvar142) || forvar152)) ?
                  (&reg149[(4'ha):(3'h4)]) : $unsigned(($unsigned(reg147) ?
                      $signed(reg156) : (reg144 ? (8'ha0) : reg149)))));
              reg160 = (~reg155[(2'h2):(2'h2)]);
            end
          else
            begin
              reg160 = (reg158 ?
                  ($signed($unsigned($signed((7'h41)))) ?
                      $unsigned($unsigned((reg143 ~^ wire131))) : reg146) : reg141[(5'h11):(3'h5)]);
              reg161 = $unsigned((reg150[(1'h0):(1'h0)] ? reg150 : reg136));
              reg162 <= forvar134;
            end
          for (forvar163 = (1'h0); (forvar163 < (2'h2)); forvar163 = (forvar163 + (1'h1)))
            begin
              reg164 <= $signed($signed((8'hb1)));
              reg165 <= ($unsigned(((&(forvar163 >>> reg160)) ?
                      (~$unsigned(reg153)) : (reg137 ?
                          reg156[(5'h11):(4'hc)] : ((7'h42) ?
                              wire128 : (7'h44))))) ?
                  $unsigned(reg138[(3'h6):(2'h3)]) : (^~reg149[(3'h5):(2'h2)]));
              reg166 <= (((8'hb7) == (-$unsigned((wire133 ?
                      wire130 : reg162)))) ?
                  ($signed($unsigned((^~forvar163))) ?
                      $unsigned((!reg141)) : (($unsigned((8'hac)) == ((8'hb1) <<< reg140)) ?
                          (^(-reg156)) : (|$unsigned(wire131)))) : $signed((!$signed($signed(reg156)))));
              reg167 = (+(~&{{reg138[(1'h0):(1'h0)], reg145[(3'h4):(2'h2)]}}));
            end
          if (wire130[(4'h9):(3'h4)])
            begin
              reg168 = reg146;
              reg169 <= (reg143 - $unsigned($signed($signed((-forvar152)))));
              reg170 = $signed($unsigned($signed(($unsigned(reg145) ?
                  $signed(forvar134) : $signed(reg146)))));
              reg171 = (reg167 ?
                  $signed(((reg150[(1'h0):(1'h0)] | (reg169 & reg166)) ?
                      reg141[(3'h4):(2'h3)] : ($signed(reg136) ?
                          $signed(reg146) : reg169[(4'h8):(2'h2)]))) : reg155[(1'h0):(1'h0)]);
            end
          else
            begin
              reg168 = $signed(((+(wire128 ?
                  $unsigned(reg140) : wire129)) > {$unsigned((reg149 ?
                      wire132 : reg166)),
                  (8'hab)}));
              reg169 <= (reg140[(3'h6):(3'h6)] ?
                  $signed((^~reg137[(4'h9):(1'h0)])) : {$signed((~{reg170,
                          reg162}))});
              reg172 <= reg166;
              reg173 = reg149[(4'h8):(1'h1)];
              reg174 <= $signed(reg169[(5'h10):(1'h0)]);
            end
        end
      reg175 = forvar135[(2'h2):(1'h1)];
    end
  assign wire176 = $signed({wire130[(2'h2):(1'h1)]});
  assign wire177 = ((($unsigned((reg159 ?
                       (8'hbc) : wire131)) <<< reg164[(1'h0):(1'h0)]) < ((wire133 ?
                       (~|reg159) : reg157) <<< reg149)) << reg158[(2'h3):(2'h2)]);
  assign wire178 = reg169[(4'h8):(3'h7)];
  assign wire179 = $unsigned((8'hb2));
  always
    @(posedge clk) begin
      for (forvar180 = (1'h0); (forvar180 < (2'h3)); forvar180 = (forvar180 + (1'h1)))
        begin
          for (forvar181 = (1'h0); (forvar181 < (1'h0)); forvar181 = (forvar181 + (1'h1)))
            begin
              reg182 <= $unsigned(($unsigned(reg137) ?
                  (+($signed(reg149) || {reg172,
                      reg158})) : $signed(((reg154 & reg138) ?
                      $unsigned(wire128) : wire177[(2'h3):(2'h2)]))));
              reg183 <= (^~(wire131 | $unsigned({$unsigned(reg150)})));
              reg184 = (|((-reg137[(3'h6):(2'h3)]) ?
                  ($signed($unsigned(wire130)) ?
                      $signed($unsigned(reg183)) : $unsigned((reg147 ?
                          reg143 : reg166))) : wire178));
            end
          reg185 = $signed((reg174 ~^ ((~(|wire130)) ?
              wire177[(2'h2):(2'h2)] : $unsigned(((8'had) ?
                  (8'ha2) : reg138)))));
          for (forvar186 = (1'h0); (forvar186 < (1'h1)); forvar186 = (forvar186 + (1'h1)))
            begin
              reg187 = $unsigned(reg136);
            end
          reg188 = reg183[(4'h8):(1'h0)];
        end
      reg189 <= (reg145[(2'h3):(1'h0)] << $unsigned(reg188[(4'hc):(3'h4)]));
      for (forvar190 = (1'h0); (forvar190 < (1'h0)); forvar190 = (forvar190 + (1'h1)))
        begin
          reg191 = $unsigned(($unsigned($signed($signed((8'hb7)))) ?
              $unsigned(wire176) : ((reg185 ?
                      (~reg158) : (wire131 ? forvar180 : reg137)) ?
                  reg157 : ((~forvar186) ?
                      $signed(forvar186) : (reg147 << reg138)))));
          for (forvar192 = (1'h0); (forvar192 < (3'h4)); forvar192 = (forvar192 + (1'h1)))
            begin
              reg193 <= (~^(reg137 || (wire131[(5'h13):(4'hf)] ^~ forvar181)));
              reg194 = $signed($signed((|($signed(reg156) ?
                  (forvar180 ? (7'h47) : reg193) : $unsigned(reg184)))));
              reg195 = ($unsigned(($unsigned({(7'h40)}) <= ({(8'ha9),
                  reg139} == reg169[(2'h3):(2'h3)]))) < forvar190[(1'h0):(1'h0)]);
              reg196 = $signed($unsigned(({$unsigned(reg149), $signed(reg194)} ?
                  reg162 : (8'ha8))));
              reg197 = $signed($signed((~$unsigned($signed((8'ha9))))));
            end
          reg198 <= ((|({$signed(wire176),
                  $signed(reg137)} && reg143[(1'h0):(1'h0)])) ?
              (wire178 < $unsigned({(reg195 ? reg165 : forvar192),
                  reg138[(3'h6):(3'h6)]})) : $signed((8'ha3)));
          for (forvar199 = (1'h0); (forvar199 < (2'h2)); forvar199 = (forvar199 + (1'h1)))
            begin
              reg200 = ($unsigned(({$unsigned(reg182)} + ((~^wire133) ^ reg196[(3'h5):(2'h2)]))) ?
                  $signed($signed($signed({reg150,
                      reg147}))) : ((reg187[(4'hc):(4'hb)] ?
                          ({forvar190, wire129} ?
                              (reg141 ?
                                  reg183 : reg138) : wire129) : ($unsigned(wire178) ?
                              $signed(reg157) : (reg166 != reg198))) ?
                      (((reg197 <= (7'h41)) - (~&reg184)) & reg157) : ({(forvar199 ?
                                  (8'ha7) : reg188)} ?
                          reg197[(3'h5):(3'h5)] : $unsigned($unsigned((8'h9e))))));
              reg201 <= ($unsigned((~$signed({reg196, reg195}))) ?
                  ($unsigned(reg182[(3'h7):(3'h7)]) ?
                      wire128[(2'h2):(2'h2)] : (7'h40)) : (^$unsigned(reg147)));
              reg202 <= (reg150[(3'h6):(1'h1)] < $unsigned((($unsigned(forvar186) <= wire132[(1'h0):(1'h0)]) ?
                  {(!reg194),
                      (reg165 ^ wire132)} : (~&reg149[(1'h0):(1'h0)]))));
              reg203 <= reg198;
            end
        end
    end
  assign wire204 = $unsigned($signed(wire129));
  always
    @(posedge clk) begin
      reg205 <= $unsigned($signed($signed((reg203[(1'h0):(1'h0)] << wire178[(2'h2):(1'h1)]))));
      reg206 <= {reg158[(2'h3):(1'h1)]};
    end
  always
    @(posedge clk) begin
      if ((7'h47))
        begin
          reg207 = (^~(8'had));
          reg208 <= ({((reg136[(1'h0):(1'h0)] - reg139) ?
                  ((reg162 >>> (8'hbf)) ?
                      $unsigned(reg145) : reg165) : ($unsigned((7'h42)) ?
                      $signed(reg159) : {reg205,
                          reg164}))} << reg154[(3'h4):(1'h1)]);
        end
      else
        begin
          reg207 = $signed($signed((reg158 ?
              (reg208[(2'h2):(1'h0)] ?
                  reg158 : reg158) : (!$unsigned(reg157)))));
          reg209 = (&$unsigned({wire176, $unsigned(reg136[(3'h4):(1'h1)])}));
        end
      reg210 = (!wire177);
      for (forvar211 = (1'h0); (forvar211 < (3'h4)); forvar211 = (forvar211 + (1'h1)))
        begin
          reg212 <= (8'haf);
          reg213 <= (reg136 != reg141);
          for (forvar214 = (1'h0); (forvar214 < (1'h1)); forvar214 = (forvar214 + (1'h1)))
            begin
              reg215 = $signed((forvar211 ?
                  reg183 : $unsigned(($unsigned(reg206) << (reg212 ?
                      reg202 : reg205)))));
            end
        end
    end
endmodule