(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param1907 = {({(~((7'h57) ? (8'hba) : (8'hb5)))} ~^ {({(8'hb3), (7'h4e), (7'h4a)} ? ((8'hb3) >> (8'ha0)) : ((8'h9c) ? (8'hbe) : (7'h49))), (((8'hb9) ? (8'hbe) : (7'h52)) ? ((7'h56) << (8'ha1)) : (-(7'h51)))}), (^~({((8'ha7) ? (8'hb3) : (7'h4c)), (|(8'ha2))} ? (((8'ha5) || (8'hbf)) != ((7'h4a) >= (8'hb6))) : (((8'hb3) ? (7'h55) : (8'ha9)) ? ((8'hb1) ? (8'ha7) : (8'ha4)) : (|(8'ha7))))), (((~&((7'h58) ? (8'hb2) : (7'h40))) + (((8'ha4) >= (7'h41)) << (&(8'hb0)))) ? {(&((7'h54) && (8'ha0))), (~^{(7'h52), (8'hb1)})} : ({(^(7'h4d))} ^~ (^(&(7'h57)))))}, 
parameter param1908 = param1907)
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h15c5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire0;
  input wire signed [(5'h1b):(1'h0)] wire1;
  input wire signed [(4'hd):(1'h0)] wire2;
  input wire [(3'h5):(1'h0)] wire3;
  input wire [(5'h17):(1'h0)] wire4;
  wire [(5'h1a):(1'h0)] wire1906;
  wire signed [(5'h13):(1'h0)] wire5;
  wire signed [(5'h1b):(1'h0)] wire137;
  wire [(3'h5):(1'h0)] wire139;
  wire [(5'h1e):(1'h0)] wire165;
  wire signed [(4'hd):(1'h0)] wire166;
  wire [(5'h12):(1'h0)] wire167;
  wire [(4'h8):(1'h0)] wire169;
  wire signed [(3'h4):(1'h0)] wire1774;
  wire [(5'h15):(1'h0)] wire1776;
  wire signed [(5'h17):(1'h0)] wire1831;
  wire signed [(5'h13):(1'h0)] wire1900;
  wire signed [(4'ha):(1'h0)] wire1902;
  wire [(3'h7):(1'h0)] wire1904;
  reg signed [(5'h12):(1'h0)] reg7 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg12 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg13 = (1'h0);
  reg [(4'h9):(1'h0)] reg14 = (1'h0);
  reg [(3'h6):(1'h0)] reg16 = (1'h0);
  reg [(5'h1f):(1'h0)] reg18 = (1'h0);
  reg [(5'h1c):(1'h0)] reg20 = (1'h0);
  reg [(5'h17):(1'h0)] reg22 = (1'h0);
  reg [(5'h11):(1'h0)] reg23 = (1'h0);
  reg [(5'h1a):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg29 = (1'h0);
  reg [(4'hd):(1'h0)] reg30 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg31 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg32 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg33 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg37 = (1'h0);
  reg signed [(4'he):(1'h0)] reg40 = (1'h0);
  reg [(5'h1e):(1'h0)] reg42 = (1'h0);
  reg [(4'hc):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg49 = (1'h0);
  reg [(5'h14):(1'h0)] reg51 = (1'h0);
  reg [(5'h10):(1'h0)] reg56 = (1'h0);
  reg [(4'hf):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg59 = (1'h0);
  reg [(4'ha):(1'h0)] reg60 = (1'h0);
  reg [(5'h1a):(1'h0)] reg63 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg64 = (1'h0);
  reg [(4'hb):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg68 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg80 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg82 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg85 = (1'h0);
  reg [(5'h15):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg93 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg95 = (1'h0);
  reg [(2'h3):(1'h0)] reg97 = (1'h0);
  reg [(3'h7):(1'h0)] reg98 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg102 = (1'h0);
  reg [(5'h1d):(1'h0)] reg105 = (1'h0);
  reg [(5'h13):(1'h0)] reg108 = (1'h0);
  reg [(5'h1b):(1'h0)] reg109 = (1'h0);
  reg [(4'h8):(1'h0)] reg111 = (1'h0);
  reg [(5'h18):(1'h0)] reg112 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg116 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg118 = (1'h0);
  reg [(5'h1b):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg124 = (1'h0);
  reg [(5'h1d):(1'h0)] reg126 = (1'h0);
  reg [(5'h1c):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg127 = (1'h0);
  reg [(5'h14):(1'h0)] reg129 = (1'h0);
  reg [(4'hb):(1'h0)] reg134 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg135 = (1'h0);
  reg [(3'h7):(1'h0)] reg136 = (1'h0);
  reg [(5'h14):(1'h0)] reg138 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg140 = (1'h0);
  reg [(4'hb):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg144 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg152 = (1'h0);
  reg [(5'h12):(1'h0)] reg154 = (1'h0);
  reg [(4'hf):(1'h0)] reg155 = (1'h0);
  reg [(5'h1b):(1'h0)] reg156 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg157 = (1'h0);
  reg [(5'h16):(1'h0)] reg161 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg170 = (1'h0);
  reg [(5'h1d):(1'h0)] reg171 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg183 = (1'h0);
  reg [(5'h1f):(1'h0)] reg186 = (1'h0);
  reg [(5'h1f):(1'h0)] reg180 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1780 = (1'h0);
  reg [(5'h18):(1'h0)] reg1783 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1784 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1787 = (1'h0);
  reg [(3'h5):(1'h0)] reg1792 = (1'h0);
  reg [(5'h18):(1'h0)] reg1793 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1795 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1796 = (1'h0);
  reg [(5'h13):(1'h0)] reg1798 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1801 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1804 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1806 = (1'h0);
  reg [(4'he):(1'h0)] reg1808 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1810 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1812 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1813 = (1'h0);
  reg [(5'h19):(1'h0)] reg1822 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1825 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1830 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1834 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1838 = (1'h0);
  reg [(4'h8):(1'h0)] reg1844 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1847 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1851 = (1'h0);
  reg [(2'h2):(1'h0)] reg1852 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1856 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1857 = (1'h0);
  reg [(5'h16):(1'h0)] reg1860 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1861 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1863 = (1'h0);
  reg [(4'h9):(1'h0)] reg1864 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1865 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1866 = (1'h0);
  reg [(5'h15):(1'h0)] reg1869 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1872 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1874 = (1'h0);
  reg [(4'hc):(1'h0)] reg1882 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1883 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1884 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1885 = (1'h0);
  reg [(5'h15):(1'h0)] reg1886 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1887 = (1'h0);
  reg [(4'hd):(1'h0)] reg1890 = (1'h0);
  reg [(5'h13):(1'h0)] reg1892 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1894 = (1'h0);
  reg [(3'h5):(1'h0)] reg1899 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1898 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1897 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1896 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1895 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1893 = (1'h0);
  reg [(5'h18):(1'h0)] reg1891 = (1'h0);
  reg [(4'ha):(1'h0)] reg1889 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1888 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1881 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1880 = (1'h0);
  reg [(3'h4):(1'h0)] reg1879 = (1'h0);
  reg [(4'h8):(1'h0)] reg1878 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1877 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1876 = (1'h0);
  reg [(5'h12):(1'h0)] reg1875 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1873 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1871 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1870 = (1'h0);
  reg [(3'h7):(1'h0)] reg1868 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1867 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1862 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1859 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1858 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1855 = (1'h0);
  reg [(3'h4):(1'h0)] reg1854 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1853 = (1'h0);
  reg [(4'hf):(1'h0)] reg1850 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1849 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1848 = (1'h0);
  reg [(3'h6):(1'h0)] reg1846 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1845 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1843 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1842 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1841 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1840 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1839 = (1'h0);
  reg [(5'h10):(1'h0)] reg1837 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1836 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1835 = (1'h0);
  reg [(4'h9):(1'h0)] reg1833 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1832 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1829 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1828 = (1'h0);
  reg [(3'h4):(1'h0)] reg1827 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1826 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1824 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1823 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1821 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1820 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1819 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1818 = (1'h0);
  reg [(4'hb):(1'h0)] reg1817 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1816 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1815 = (1'h0);
  reg [(2'h3):(1'h0)] reg1814 = (1'h0);
  reg [(4'hb):(1'h0)] reg1811 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1809 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1807 = (1'h0);
  reg [(5'h12):(1'h0)] reg1805 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1803 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1799 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1802 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1800 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1799 = (1'h0);
  reg [(5'h10):(1'h0)] reg1797 = (1'h0);
  reg [(4'hd):(1'h0)] reg1794 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1791 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1790 = (1'h0);
  reg [(5'h19):(1'h0)] reg1789 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1788 = (1'h0);
  reg [(4'ha):(1'h0)] reg1786 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1785 = (1'h0);
  reg [(4'he):(1'h0)] reg1782 = (1'h0);
  reg [(2'h3):(1'h0)] reg1781 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1779 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar1778 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1777 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg188 = (1'h0);
  reg [(3'h4):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg185 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg184 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar180 = (1'h0);
  reg [(3'h5):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg178 = (1'h0);
  reg [(5'h13):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg175 = (1'h0);
  reg [(3'h6):(1'h0)] reg172 = (1'h0);
  reg [(4'h9):(1'h0)] reg164 = (1'h0);
  reg [(5'h1b):(1'h0)] reg163 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg162 = (1'h0);
  reg [(5'h1b):(1'h0)] reg160 = (1'h0);
  reg [(4'h8):(1'h0)] reg159 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg158 = (1'h0);
  reg [(3'h4):(1'h0)] reg153 = (1'h0);
  reg [(5'h17):(1'h0)] reg151 = (1'h0);
  reg [(3'h5):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg149 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg146 = (1'h0);
  reg [(5'h16):(1'h0)] forvar144 = (1'h0);
  reg [(5'h18):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg142 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar133 = (1'h0);
  reg [(5'h1d):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar130 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg128 = (1'h0);
  reg [(2'h2):(1'h0)] forvar118 = (1'h0);
  reg [(5'h10):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg123 = (1'h0);
  reg [(4'hd):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar120 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg117 = (1'h0);
  reg [(4'ha):(1'h0)] reg115 = (1'h0);
  reg [(5'h1a):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg107 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg103 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg101 = (1'h0);
  reg [(4'h9):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg96 = (1'h0);
  reg [(4'hf):(1'h0)] forvar94 = (1'h0);
  reg [(5'h10):(1'h0)] reg91 = (1'h0);
  reg [(5'h1f):(1'h0)] reg90 = (1'h0);
  reg [(3'h7):(1'h0)] forvar88 = (1'h0);
  reg [(5'h1a):(1'h0)] reg87 = (1'h0);
  reg [(5'h19):(1'h0)] forvar86 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar75 = (1'h0);
  reg [(4'ha):(1'h0)] forvar84 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg81 = (1'h0);
  reg [(3'h6):(1'h0)] reg76 = (1'h0);
  reg [(5'h1c):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg74 = (1'h0);
  reg [(5'h1a):(1'h0)] reg73 = (1'h0);
  reg [(5'h16):(1'h0)] reg72 = (1'h0);
  reg [(5'h16):(1'h0)] forvar71 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg70 = (1'h0);
  reg [(5'h17):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg66 = (1'h0);
  reg [(5'h13):(1'h0)] reg65 = (1'h0);
  reg [(3'h6):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg61 = (1'h0);
  reg [(5'h17):(1'h0)] forvar54 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg57 = (1'h0);
  reg [(3'h5):(1'h0)] reg55 = (1'h0);
  reg [(4'ha):(1'h0)] reg54 = (1'h0);
  reg [(2'h3):(1'h0)] forvar53 = (1'h0);
  reg [(5'h16):(1'h0)] reg52 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar50 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg48 = (1'h0);
  reg [(5'h19):(1'h0)] reg46 = (1'h0);
  reg signed [(4'he):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg44 = (1'h0);
  reg [(2'h3):(1'h0)] reg43 = (1'h0);
  reg [(5'h17):(1'h0)] reg41 = (1'h0);
  reg [(5'h17):(1'h0)] reg39 = (1'h0);
  reg [(5'h13):(1'h0)] reg38 = (1'h0);
  reg [(2'h3):(1'h0)] reg36 = (1'h0);
  reg [(2'h3):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg34 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg27 = (1'h0);
  reg [(3'h7):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg24 = (1'h0);
  reg [(5'h17):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg19 = (1'h0);
  reg [(5'h17):(1'h0)] reg17 = (1'h0);
  reg [(5'h15):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg10 = (1'h0);
  reg [(3'h5):(1'h0)] reg9 = (1'h0);
  reg [(5'h13):(1'h0)] reg8 = (1'h0);
  reg [(5'h14):(1'h0)] forvar6 = (1'h0);
  assign y = {wire1906,
                 wire5,
                 wire137,
                 wire139,
                 wire165,
                 wire166,
                 wire167,
                 wire169,
                 wire1774,
                 wire1776,
                 wire1831,
                 wire1900,
                 wire1902,
                 wire1904,
                 reg7,
                 reg12,
                 reg13,
                 reg14,
                 reg16,
                 reg18,
                 reg20,
                 reg22,
                 reg23,
                 reg26,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 reg37,
                 reg40,
                 reg42,
                 reg47,
                 reg49,
                 reg51,
                 reg56,
                 reg50,
                 reg58,
                 reg59,
                 reg60,
                 reg63,
                 reg64,
                 reg67,
                 reg68,
                 reg77,
                 reg78,
                 reg79,
                 reg80,
                 reg82,
                 reg85,
                 reg84,
                 reg89,
                 reg92,
                 reg93,
                 reg95,
                 reg97,
                 reg98,
                 reg102,
                 reg105,
                 reg108,
                 reg109,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 reg116,
                 reg118,
                 reg122,
                 reg124,
                 reg126,
                 reg120,
                 reg127,
                 reg129,
                 reg134,
                 reg135,
                 reg136,
                 reg138,
                 reg140,
                 reg145,
                 reg147,
                 reg144,
                 reg152,
                 reg154,
                 reg155,
                 reg156,
                 reg157,
                 reg161,
                 reg168,
                 reg170,
                 reg171,
                 reg173,
                 reg174,
                 reg176,
                 reg182,
                 reg183,
                 reg186,
                 reg180,
                 reg1780,
                 reg1783,
                 reg1784,
                 reg1787,
                 reg1792,
                 reg1793,
                 reg1795,
                 reg1796,
                 reg1798,
                 reg1801,
                 reg1804,
                 reg1806,
                 reg1808,
                 reg1810,
                 reg1812,
                 reg1813,
                 reg1822,
                 reg1825,
                 reg1830,
                 reg1834,
                 reg1838,
                 reg1844,
                 reg1847,
                 reg1851,
                 reg1852,
                 reg1856,
                 reg1857,
                 reg1860,
                 reg1861,
                 reg1863,
                 reg1864,
                 reg1865,
                 reg1866,
                 reg1869,
                 reg1872,
                 reg1874,
                 reg1882,
                 reg1883,
                 reg1884,
                 reg1885,
                 reg1886,
                 reg1887,
                 reg1890,
                 reg1892,
                 reg1894,
                 reg1899,
                 forvar1898,
                 reg1897,
                 reg1896,
                 reg1895,
                 forvar1893,
                 reg1891,
                 reg1889,
                 reg1888,
                 reg1881,
                 reg1880,
                 reg1879,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1875,
                 reg1873,
                 reg1871,
                 reg1870,
                 reg1868,
                 reg1867,
                 reg1862,
                 forvar1859,
                 reg1858,
                 reg1855,
                 reg1854,
                 reg1853,
                 reg1850,
                 reg1849,
                 reg1848,
                 reg1846,
                 reg1845,
                 reg1843,
                 forvar1842,
                 reg1841,
                 reg1840,
                 reg1839,
                 reg1837,
                 reg1836,
                 reg1835,
                 reg1833,
                 forvar1832,
                 reg1829,
                 reg1828,
                 reg1827,
                 reg1826,
                 reg1824,
                 forvar1823,
                 reg1821,
                 reg1820,
                 reg1819,
                 reg1818,
                 reg1817,
                 forvar1816,
                 forvar1815,
                 reg1814,
                 reg1811,
                 forvar1809,
                 reg1807,
                 reg1805,
                 reg1803,
                 reg1799,
                 reg1802,
                 reg1800,
                 forvar1799,
                 reg1797,
                 reg1794,
                 reg1791,
                 reg1790,
                 reg1789,
                 reg1788,
                 reg1786,
                 reg1785,
                 reg1782,
                 reg1781,
                 reg1779,
                 forvar1778,
                 forvar1777,
                 reg188,
                 reg187,
                 reg185,
                 reg184,
                 reg181,
                 forvar180,
                 reg179,
                 reg178,
                 reg177,
                 reg175,
                 reg172,
                 reg164,
                 reg163,
                 reg162,
                 reg160,
                 reg159,
                 reg158,
                 reg153,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg146,
                 forvar144,
                 reg143,
                 reg142,
                 reg141,
                 forvar133,
                 reg132,
                 reg131,
                 forvar130,
                 reg128,
                 forvar118,
                 reg125,
                 reg123,
                 reg121,
                 forvar120,
                 reg119,
                 reg117,
                 reg115,
                 reg110,
                 reg107,
                 reg106,
                 reg104,
                 reg103,
                 reg101,
                 reg100,
                 reg99,
                 reg96,
                 forvar94,
                 reg91,
                 reg90,
                 forvar88,
                 reg87,
                 forvar86,
                 forvar75,
                 forvar84,
                 reg83,
                 reg81,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 forvar71,
                 reg70,
                 reg69,
                 reg66,
                 reg65,
                 reg62,
                 reg61,
                 forvar54,
                 reg53,
                 reg57,
                 reg55,
                 reg54,
                 forvar53,
                 reg52,
                 forvar50,
                 reg48,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg41,
                 reg39,
                 reg38,
                 reg36,
                 reg35,
                 reg34,
                 reg28,
                 reg27,
                 reg25,
                 reg24,
                 reg21,
                 reg19,
                 reg17,
                 reg15,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 forvar6,
                 (1'h0)};
  assign wire5 = wire4[(3'h7):(3'h5)];
  always
    @(posedge clk) begin
      for (forvar6 = (1'h0); (forvar6 < (3'h6)); forvar6 = (forvar6 + (1'h1)))
        begin
          if (($signed(wire0[(2'h2):(1'h0)]) ^~ $unsigned($signed(wire3[(1'h0):(1'h0)]))))
            begin
              reg7 <= (&(wire3[(3'h4):(2'h3)] | $signed(({wire2} && (wire4 ~^ wire4)))));
            end
          else
            begin
              reg7 <= forvar6[(3'h4):(1'h1)];
            end
          if (($unsigned(wire5) > reg7[(3'h4):(1'h0)]))
            begin
              reg8 = wire2;
              reg9 = (~(7'h47));
              reg10 = (wire1 != wire4[(1'h0):(1'h0)]);
              reg11 = (forvar6 ? reg9 : wire5);
              reg12 <= ($signed(wire0) >> wire3);
              reg13 <= (reg9[(3'h5):(3'h5)] ?
                  ($unsigned(($unsigned((8'haf)) + (8'hb1))) ?
                      $unsigned((~reg12)) : (wire4[(5'h11):(3'h7)] + (reg11 ?
                          $signed(reg12) : (wire2 ?
                              reg9 : (8'hbb))))) : $signed((^{(~&(7'h55)),
                      reg8})));
            end
          else
            begin
              reg8 = (reg13[(4'h9):(2'h2)] ?
                  reg8 : ($unsigned(wire4) ?
                      ((^~(wire2 < wire5)) && $unsigned(reg8)) : (~^({reg7} ?
                          (reg10 == wire4) : $unsigned(reg8)))));
              reg9 = $unsigned($unsigned($unsigned($unsigned((wire2 <= reg9)))));
              reg10 = (~$signed(((~&reg12[(1'h1):(1'h0)]) ^~ $unsigned((-reg8)))));
            end
          if ($signed(((^$signed(wire3)) ?
              ($signed(reg8) ?
                  (^(~^(8'ha9))) : reg9[(3'h4):(1'h1)]) : (+$unsigned($signed(reg11))))))
            begin
              reg14 <= reg10[(4'hf):(3'h4)];
              reg15 = $unsigned(($unsigned(($unsigned(wire2) ?
                      (|reg8) : (^~reg8))) ?
                  (&$unsigned($unsigned(wire4))) : reg7[(2'h2):(1'h0)]));
              reg16 <= $signed(reg10[(2'h3):(1'h1)]);
              reg17 = reg12[(1'h1):(1'h1)];
              reg18 <= $signed((-$unsigned((wire5 ?
                  (reg11 <<< wire3) : (+reg9)))));
            end
          else
            begin
              reg15 = (forvar6[(4'h9):(2'h3)] ?
                  wire1 : $unsigned(({$signed(reg12)} ~^ wire4[(4'h8):(3'h7)])));
              reg17 = reg18[(5'h14):(4'hc)];
              reg19 = reg16;
              reg20 <= $signed(reg16[(3'h5):(2'h2)]);
              reg21 = wire4[(4'ha):(1'h0)];
              reg22 <= wire4[(5'h12):(4'hf)];
              reg23 <= (&((-$signed($unsigned(reg19))) < ({(~^reg18),
                  (8'h9c)} < (~^reg14))));
            end
          reg24 = (wire0 || (wire4 ?
              (^{reg11[(2'h2):(2'h2)],
                  (^reg21),
                  {wire2, reg20}}) : ((reg9[(3'h5):(1'h1)] ?
                  reg18[(4'he):(3'h7)] : reg13) - (8'hb8))));
          if ($signed($unsigned((~(7'h46)))))
            begin
              reg25 = $signed({($signed((~reg23)) ^ ((wire3 ?
                      wire2 : reg20) - $unsigned((8'hb7)))),
                  reg9[(2'h3):(1'h1)]});
              reg26 <= (wire2[(4'hb):(4'ha)] == $signed($unsigned({$unsigned(reg12)})));
              reg27 = (reg16[(3'h4):(2'h2)] * $signed((({wire5} ?
                      $unsigned((8'hac)) : (forvar6 ? reg24 : reg19)) ?
                  ($unsigned(wire3) * reg22) : ((wire5 < reg20) ?
                      reg19[(4'ha):(3'h7)] : (reg21 ? reg10 : reg16)))));
              reg28 = reg7[(5'h11):(4'hc)];
            end
          else
            begin
              reg26 <= ((8'hbc) >>> $signed($signed({$unsigned((7'h40)),
                  (~reg27)})));
              reg27 = (8'ha7);
              reg28 = {$signed((($unsigned(wire3) ?
                      (reg25 ?
                          forvar6 : reg27) : $unsigned(wire0)) | $unsigned(reg22[(2'h2):(1'h0)]))),
                  $unsigned((~|(reg14[(2'h3):(1'h0)] < reg15[(5'h13):(5'h10)])))};
            end
        end
    end
  always
    @(posedge clk) begin
      if ((^~(^~($signed($unsigned(wire0)) >= ((reg22 ? wire5 : reg26) ?
          (reg16 ^ reg7) : {reg26})))))
        begin
          reg29 <= $unsigned($unsigned(($unsigned($unsigned(wire2)) | reg16[(1'h0):(1'h0)])));
          reg30 <= wire2[(4'h9):(1'h1)];
          if ((wire3[(2'h3):(1'h0)] ?
              (($unsigned($unsigned((7'h53))) <<< (8'hb4)) ?
                  $unsigned(($signed(reg26) > (wire5 ?
                      reg14 : wire0))) : ({wire4[(5'h12):(4'hc)],
                          ((8'hb7) ? wire5 : reg23)} ?
                      {$signed(reg18),
                          (reg13 ? reg18 : reg7),
                          (reg20 ? reg30 : reg23)} : ($unsigned(reg14) ?
                          (!reg18) : reg20[(3'h5):(2'h3)]))) : ($unsigned((!(~reg7))) && $unsigned(wire1[(4'he):(4'hd)]))))
            begin
              reg31 <= $signed(wire0);
              reg32 <= ($signed(wire3) ?
                  ($unsigned((|(reg12 << wire5))) <<< ($signed((+reg23)) ?
                      $signed(reg23) : reg7)) : reg26[(4'he):(4'hb)]);
              reg33 <= (^(((~(~|wire0)) > wire0[(2'h2):(1'h0)]) ?
                  ((~^{reg14, reg30}) ?
                      $signed(((8'ha1) <= (8'h9e))) : reg7[(5'h12):(4'hb)]) : $unsigned((~&(reg13 ?
                      reg23 : (8'h9f))))));
              reg34 = $signed((((7'h47) * wire3[(1'h0):(1'h0)]) >= wire1[(3'h7):(2'h2)]));
              reg35 = $unsigned($signed(reg33[(1'h1):(1'h0)]));
              reg36 = $signed($unsigned(($signed((wire1 ?
                  reg13 : reg18)) ~^ ((-reg35) >> (~^reg35)))));
            end
          else
            begin
              reg31 <= (reg30[(3'h4):(1'h1)] ^ $signed(reg7));
              reg32 <= ($unsigned({$unsigned((&wire4)),
                  reg30,
                  {reg20,
                      {reg22},
                      reg22[(3'h6):(1'h0)]}}) < wire4[(5'h16):(4'hf)]);
              reg33 <= {reg12[(3'h4):(1'h1)]};
              reg34 = $unsigned(reg13);
              reg37 <= reg18;
            end
        end
      else
        begin
          reg34 = reg37;
          if (((reg32[(1'h0):(1'h0)] ?
              (~(reg23 ?
                  (reg12 <= reg26) : reg36[(2'h3):(1'h1)])) : (reg29[(1'h1):(1'h1)] ?
                  ((-reg12) && reg18) : $signed((&reg14)))) & reg16[(3'h6):(2'h3)]))
            begin
              reg37 <= reg37[(2'h2):(2'h2)];
              reg38 = (&(+$signed((((8'hb7) ?
                  wire5 : reg13) <<< $unsigned(reg37)))));
              reg39 = wire0[(2'h3):(1'h1)];
              reg40 <= reg34;
            end
          else
            begin
              reg35 = ((reg14[(1'h0):(1'h0)] ?
                      {$unsigned($signed(reg40)),
                          ($signed(reg12) ?
                              $signed(wire3) : $unsigned((8'hba)))} : (!$unsigned((^reg36)))) ?
                  reg37[(1'h0):(1'h0)] : wire3[(2'h2):(1'h0)]);
              reg36 = ($unsigned(reg23) ^~ (reg33 ?
                  ((+$unsigned(reg33)) >= reg20[(4'hf):(1'h1)]) : $unsigned({reg20})));
            end
        end
      reg41 = (|{reg7,
          ((^~reg18[(5'h11):(4'he)]) ?
              (7'h4c) : ((wire0 ? reg32 : (8'had)) && (~|wire0)))});
      if (($signed($unsigned($unsigned((reg20 + reg32)))) ?
          (((~&(reg32 ?
              reg41 : reg36)) && (&(wire4 * wire3))) >> (reg12[(3'h4):(1'h1)] >= (&(reg22 ?
              reg20 : reg40)))) : $unsigned((reg40 > {reg33[(3'h7):(2'h3)],
              $unsigned(wire5)}))))
        begin
          if (reg40)
            begin
              reg42 <= (((7'h57) ^~ (((&reg7) | $signed(reg7)) ?
                      ($unsigned(reg31) != (reg12 && reg31)) : {(^~(7'h41)),
                          wire5})) ?
                  $unsigned($signed($unsigned((reg34 ?
                      wire1 : wire0)))) : (~reg14));
            end
          else
            begin
              reg43 = reg35[(2'h2):(2'h2)];
            end
          if ((~($unsigned((^((8'hb8) ? reg39 : reg20))) ?
              wire3 : wire5[(4'hb):(4'h9)])))
            begin
              reg44 = (|reg16);
              reg45 = ($signed(wire3[(2'h2):(1'h1)]) ?
                  {reg33,
                      {(~^(reg43 ? (8'hbf) : reg36))},
                      (~^reg14[(3'h5):(3'h4)])} : reg36);
              reg46 = ($unsigned((^~($unsigned(reg20) && (reg35 <= reg13)))) ?
                  ((reg13[(4'ha):(3'h4)] ?
                      $signed($signed(wire2)) : (~^{reg30,
                          reg45})) != (^$unsigned((reg42 & reg12)))) : {(8'h9d),
                      reg37});
            end
          else
            begin
              reg44 = reg41[(4'hc):(3'h4)];
              reg45 = ((~reg23) ^ $signed(wire0[(3'h5):(2'h3)]));
            end
          if ($unsigned((reg39 <= reg35)))
            begin
              reg47 <= $unsigned({reg34, (-reg33[(2'h2):(1'h0)])});
            end
          else
            begin
              reg48 = ((reg30 << ((~^reg39[(3'h5):(2'h2)]) * (+reg45[(1'h0):(1'h0)]))) ?
                  $signed(reg47[(4'h9):(3'h6)]) : (-reg42[(5'h13):(4'h9)]));
              reg49 <= wire0[(2'h2):(1'h0)];
            end
          for (forvar50 = (1'h0); (forvar50 < (2'h2)); forvar50 = (forvar50 + (1'h1)))
            begin
              reg51 <= reg26[(4'hf):(2'h3)];
              reg52 = $unsigned((&(8'hba)));
            end
          for (forvar53 = (1'h0); (forvar53 < (1'h1)); forvar53 = (forvar53 + (1'h1)))
            begin
              reg54 = reg14[(3'h5):(2'h2)];
              reg55 = reg45;
            end
          reg56 <= wire0;
          reg57 = wire4;
        end
      else
        begin
          reg43 = $unsigned({(((reg44 != reg36) <<< {reg33}) ?
                  reg20[(1'h1):(1'h1)] : $unsigned($signed(reg18))),
              $signed(forvar53[(2'h2):(2'h2)]),
              reg49});
          reg44 = $unsigned((reg56[(1'h1):(1'h0)] ?
              ((7'h4a) <<< ((reg38 ? reg33 : (7'h46)) ?
                  (!reg46) : $unsigned(reg44))) : reg22));
          if ($signed($signed(reg31)))
            begin
              reg47 <= $unsigned($unsigned($signed({{reg57, reg31, wire5},
                  reg37,
                  (reg33 && reg38)})));
              reg48 = reg44;
              reg49 <= $unsigned(reg18);
              reg50 <= $signed(($unsigned($signed(reg39[(1'h0):(1'h0)])) == (8'hb3)));
              reg51 <= reg45;
              reg52 = ($signed($signed(((reg37 ?
                  reg44 : (7'h56)) >>> $signed(wire2)))) < $unsigned({($signed(reg20) > (~^reg56))}));
            end
          else
            begin
              reg47 <= (~^$signed(((!{reg30, reg26}) ?
                  (8'h9c) : $unsigned(wire3))));
              reg49 <= {forvar53[(1'h1):(1'h1)],
                  ((~$unsigned($unsigned((8'hbd)))) ?
                      $unsigned(((reg37 ?
                          reg37 : reg39) <<< reg35[(1'h1):(1'h1)])) : reg44)};
            end
          reg53 = reg32;
          for (forvar54 = (1'h0); (forvar54 < (3'h6)); forvar54 = (forvar54 + (1'h1)))
            begin
              reg55 = $signed(({$signed(((8'hba) > reg26))} ^ reg18[(2'h3):(2'h2)]));
              reg56 <= (8'ha6);
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned(((reg56 ?
          ((~reg47) ?
              $signed(reg32) : reg13[(3'h5):(3'h5)]) : ((reg14 > reg26) ?
              (wire0 || reg20) : reg56)) != reg22)))
        begin
          if ((({reg31[(1'h0):(1'h0)]} | $unsigned(reg37[(2'h2):(1'h0)])) ^~ (8'hac)))
            begin
              reg58 <= ((({reg50, (reg40 >= (7'h48))} >> (+$unsigned(reg56))) ?
                      reg23[(1'h1):(1'h1)] : $unsigned((-(-reg23)))) ?
                  {reg37[(2'h2):(1'h0)],
                      reg23,
                      $unsigned($unsigned($unsigned(reg12)))} : $signed((wire5 ?
                      $signed($unsigned(reg13)) : $signed((-reg20)))));
              reg59 <= (~^($unsigned($signed(reg12)) ?
                  $signed($signed({reg22})) : wire0));
              reg60 <= $unsigned(reg33);
              reg61 = (($signed(reg18) ?
                  $unsigned((reg23 < reg31[(1'h1):(1'h0)])) : $signed((~|$signed(reg32)))) * ((+(reg16 != ((7'h4a) ^ reg58))) || $signed(((reg60 << reg31) != {reg20,
                  wire5}))));
            end
          else
            begin
              reg58 <= (!reg40[(1'h0):(1'h0)]);
              reg61 = reg60[(2'h2):(1'h0)];
              reg62 = ((^~reg16) << (~|((reg20[(4'hf):(1'h0)] ^ (wire1 - (8'hb8))) ?
                  reg42 : reg12)));
              reg63 <= ($signed($unsigned($unsigned($signed(reg16)))) ?
                  (reg18[(3'h7):(1'h1)] ?
                      ({{(8'hbb), wire3}} ?
                          (~^(~reg12)) : $unsigned(reg16[(1'h1):(1'h1)])) : ($unsigned((~&wire1)) ?
                          (reg58 <<< reg13) : $unsigned((reg30 ?
                              wire4 : (8'hb9))))) : (~|$signed(($signed(reg62) ?
                      (~|wire5) : {reg62}))));
              reg64 <= (reg61[(2'h2):(1'h0)] ? reg22[(5'h16):(2'h2)] : reg37);
              reg65 = reg62;
              reg66 = {($unsigned($signed((^reg7))) ~^ (((reg47 ?
                          wire3 : reg29) ?
                      $signed(reg20) : $signed(reg64)) <<< reg64)),
                  {(~|{(wire1 != reg58),
                          (reg31 ? (8'hb4) : reg30),
                          ((7'h4f) ? wire4 : wire2)}),
                      wire5[(5'h10):(4'ha)]},
                  $unsigned(reg20[(5'h1b):(3'h6)])};
            end
          reg67 <= reg66[(4'h8):(2'h3)];
          reg68 <= (-$signed(wire5[(4'h9):(4'h8)]));
          reg69 = reg16;
          reg70 = $unsigned($unsigned(reg42[(5'h1e):(5'h11)]));
          for (forvar71 = (1'h0); (forvar71 < (3'h6)); forvar71 = (forvar71 + (1'h1)))
            begin
              reg72 = ($unsigned(((reg13 ?
                  (^~(8'hb6)) : (reg47 ? (8'hbb) : reg42)) <= (!(wire4 ?
                  reg70 : reg58)))) <<< (|reg12[(3'h6):(3'h6)]));
            end
          reg73 = ((+(reg62 ? wire5 : $signed($unsigned(reg16)))) ?
              $signed({(~^$signed((7'h43)))}) : ((~^(|{reg42,
                      (7'h43),
                      wire3})) ?
                  (+$signed((reg49 ?
                      (7'h40) : reg50))) : (^~reg56[(1'h0):(1'h0)])));
        end
      else
        begin
          reg61 = (($signed($unsigned(reg73[(5'h18):(5'h11)])) ?
                  reg37[(2'h2):(2'h2)] : reg22) ?
              (reg13[(3'h6):(1'h1)] && $unsigned(($signed(reg47) - (reg63 & reg60)))) : $signed(reg56[(2'h2):(1'h1)]));
          reg62 = $signed((($signed((reg51 ?
              wire4 : reg14)) > $unsigned(reg16)) + $unsigned(($signed(reg16) ?
              $signed(reg60) : reg50))));
          reg65 = $signed(((~^(|wire4)) < ((^~(reg70 && reg65)) >> $unsigned((reg14 ^ reg60)))));
        end
      if (wire3[(1'h0):(1'h0)])
        begin
          reg74 = ($signed({(((8'haf) ? reg68 : reg68) && (8'hab))}) ?
              (|forvar71[(3'h5):(1'h0)]) : $signed((^~wire3)));
          reg75 = $unsigned(($signed($unsigned($unsigned(reg66))) <<< ((~$signed(reg56)) ?
              forvar71[(4'hb):(2'h3)] : ((reg60 | forvar71) ?
                  (~&reg66) : (wire1 + reg40)))));
          if ((reg14[(3'h6):(2'h2)] & $signed((reg16 ~^ (8'h9e)))))
            begin
              reg76 = (~|(($unsigned(reg58) ?
                      $signed(reg31) : $unsigned((reg63 > reg32))) ?
                  (^~(+(reg74 | reg62))) : ({reg62,
                          (reg74 ? reg49 : reg18),
                          {(8'hba), (7'h50)}} ?
                      reg63[(5'h10):(4'h8)] : (7'h58))));
              reg77 <= reg75[(4'hf):(3'h5)];
              reg78 <= reg26;
              reg79 <= {reg61[(5'h1a):(3'h6)]};
              reg80 <= reg67;
            end
          else
            begin
              reg76 = ((|(({reg76} ? (-reg75) : ((7'h55) ? wire1 : reg32)) ?
                  reg80 : ((reg26 << reg42) | (reg12 ?
                      reg40 : reg70)))) | ({$signed({reg50})} | $unsigned(($signed(reg33) - (^~reg61)))));
              reg77 <= $signed(reg78[(1'h1):(1'h0)]);
            end
          if ($signed((reg18 + (reg32[(1'h1):(1'h1)] != (~^reg77[(3'h4):(2'h3)])))))
            begin
              reg81 = ($signed(((^reg64[(5'h10):(4'hd)]) ?
                      $unsigned({wire4, (8'haa)}) : (~|$signed(reg77)))) ?
                  $unsigned({reg29,
                      (^~reg65[(1'h0):(1'h0)])}) : reg18[(3'h4):(2'h2)]);
              reg82 <= forvar71[(4'he):(3'h4)];
              reg83 = ($signed(wire3[(3'h4):(2'h2)]) * reg76);
            end
          else
            begin
              reg82 <= {$signed($signed({reg61[(5'h1a):(4'hf)],
                      (reg79 ? reg32 : reg18),
                      (reg72 >>> (7'h40))}))};
            end
          for (forvar84 = (1'h0); (forvar84 < (3'h6)); forvar84 = (forvar84 + (1'h1)))
            begin
              reg85 <= $unsigned(({((reg65 - wire1) ?
                          (reg82 && reg12) : $signed(reg79)),
                      $unsigned(wire5)} ?
                  ((~^(^(7'h47))) ? reg60 : reg82[(2'h2):(2'h2)]) : reg14));
            end
        end
      else
        begin
          reg74 = reg26[(1'h0):(1'h0)];
          for (forvar75 = (1'h0); (forvar75 < (3'h6)); forvar75 = (forvar75 + (1'h1)))
            begin
              reg77 <= {$unsigned($unsigned(reg37))};
              reg78 <= (|(-$signed(reg31[(1'h1):(1'h1)])));
              reg81 = $unsigned($signed(((reg12 ^~ {reg14}) >> ($signed(reg73) ?
                  {reg22, wire1} : $unsigned((8'hb1))))));
              reg82 <= $signed($unsigned($signed(reg7[(1'h1):(1'h0)])));
              reg84 <= {reg70};
            end
        end
      for (forvar86 = (1'h0); (forvar86 < (3'h6)); forvar86 = (forvar86 + (1'h1)))
        begin
          reg87 = ((~reg63[(3'h7):(3'h6)]) ?
              ((&((!reg16) ? reg23[(3'h6):(1'h1)] : (reg16 ^ reg26))) ?
                  ({{(8'ha1), reg68, (8'h9e)}, (^~reg7)} ^~ $signed((reg74 ?
                      reg22 : (8'hb4)))) : $signed(reg80)) : {reg26[(3'h7):(3'h6)],
                  ($signed($signed(wire0)) ?
                      {reg73[(4'he):(4'h9)]} : $unsigned($signed((8'hb4))))});
          for (forvar88 = (1'h0); (forvar88 < (1'h1)); forvar88 = (forvar88 + (1'h1)))
            begin
              reg89 <= $unsigned($signed(((forvar86[(3'h6):(2'h3)] ?
                  {reg85,
                      forvar88,
                      forvar84} : reg31[(1'h1):(1'h0)]) < (reg67[(3'h6):(3'h4)] == (reg20 >> (8'ha7))))));
              reg90 = (7'h46);
              reg91 = {((reg37[(1'h1):(1'h1)] ?
                          (wire3 ?
                              $signed(wire2) : $signed((7'h51))) : $unsigned((reg59 ?
                              (8'hb3) : (7'h4a)))) ?
                      $signed(reg65[(4'h9):(2'h2)]) : reg42),
                  $signed($unsigned(({reg33} ?
                      (reg42 ? reg69 : reg60) : (~reg13))))};
            end
          reg92 <= reg83;
          reg93 <= $unsigned((+$unsigned($signed({reg31}))));
          for (forvar94 = (1'h0); (forvar94 < (2'h2)); forvar94 = (forvar94 + (1'h1)))
            begin
              reg95 <= (^(7'h44));
            end
          if (((&(wire0 < reg95)) ~^ $unsigned((~&$unsigned(reg16)))))
            begin
              reg96 = ({(~|$signed((reg85 <= wire5)))} ?
                  reg65[(5'h12):(3'h6)] : ((reg84 ?
                          ((wire0 ? (7'h49) : wire3) ?
                              reg93 : reg69) : $signed(reg74[(5'h18):(2'h3)])) ?
                      reg22 : ($unsigned($unsigned(reg40)) || (|$unsigned(forvar75)))));
              reg97 <= ((((+((8'ha6) != reg74)) ^ (8'hab)) ^~ $unsigned(((reg75 <= reg92) ?
                  (8'hbb) : $unsigned((7'h4a))))) ~^ (((reg90 ?
                  {reg92} : reg74[(4'hc):(3'h5)]) != $unsigned({reg73,
                  reg13,
                  (8'hb7)})) ^ {(reg20[(5'h14):(5'h14)] ?
                      $signed(wire5) : $signed(wire5))}));
              reg98 <= reg26;
            end
          else
            begin
              reg97 <= ({((forvar75 <<< reg49[(4'hb):(3'h6)]) ?
                          ((~|reg85) ?
                              (reg16 ?
                                  reg76 : reg7) : reg59[(4'ha):(4'ha)]) : ((^~reg49) ?
                              (reg95 ? wire1 : (7'h41)) : $signed(reg18))),
                      (8'had)} ?
                  $signed(forvar71[(1'h0):(1'h0)]) : reg89);
              reg98 <= (({reg18} ~^ $signed($unsigned((forvar84 >> (7'h58))))) ~^ $unsigned($signed(forvar75[(5'h18):(4'ha)])));
              reg99 = $unsigned(($signed((&reg70[(2'h2):(1'h1)])) <= $signed(forvar88[(3'h6):(1'h0)])));
              reg100 = (8'h9d);
              reg101 = $unsigned($unsigned((($unsigned(reg50) ^~ (~reg75)) >= (^(wire3 ?
                  reg23 : reg63)))));
              reg102 <= reg23;
              reg103 = ((reg37 ? reg95 : $unsigned(reg102)) ?
                  reg92[(4'h9):(3'h4)] : $signed($signed($signed({wire0,
                      forvar75,
                      reg83}))));
            end
          if ($unsigned($unsigned(({(wire5 ? reg50 : (8'hb8))} ~^ reg78))))
            begin
              reg104 = $signed($signed($signed(reg102[(2'h3):(1'h0)])));
              reg105 <= $unsigned($signed(wire3[(1'h0):(1'h0)]));
              reg106 = reg97;
              reg107 = reg42;
            end
          else
            begin
              reg105 <= ((~^(reg72[(4'h9):(1'h0)] ^ ($signed((8'hbe)) ?
                      reg62[(2'h2):(1'h0)] : (^reg80)))) ?
                  $unsigned($unsigned(($signed(reg64) >= ((8'ha6) & (7'h46))))) : (^~reg20[(5'h17):(5'h13)]));
              reg108 <= ($signed((((reg18 ^~ reg56) >= (reg84 ?
                          reg64 : reg23)) ?
                      $signed(reg69[(1'h1):(1'h0)]) : $signed((7'h49)))) ?
                  ({{{reg50, forvar88}}, $unsigned((reg68 ? reg73 : reg12))} ?
                      reg97 : reg66) : $signed($unsigned(((reg14 ?
                      (8'hbf) : (8'hbb)) ~^ $signed(reg75)))));
              reg109 <= reg50[(3'h5):(1'h1)];
              reg110 = ((8'ha3) | (reg100 ?
                  ($unsigned((8'hbd)) ?
                      ($unsigned(reg79) ^ (~^reg91)) : {(~&reg92),
                          (+reg29),
                          (reg12 == reg74)}) : (($signed((8'hb8)) || (~^reg102)) ^~ (~$unsigned(reg33)))));
              reg111 <= (reg29[(3'h6):(3'h4)] ?
                  reg107[(1'h1):(1'h1)] : (($signed((~|reg82)) ?
                      forvar86[(5'h12):(1'h1)] : {(~&reg101),
                          (7'h43),
                          (~^(8'hba))}) == reg68));
              reg112 <= (!($unsigned({$signed(reg69), $signed((7'h53))}) ?
                  ($signed(reg87) ~^ $unsigned((reg93 ?
                      reg81 : reg92))) : $signed($signed(reg30))));
              reg113 <= reg87[(2'h2):(2'h2)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg114 <= reg20;
      reg115 = reg114;
      reg116 <= ((8'hba) ?
          (7'h4d) : ({((^~reg77) ?
                      (reg67 ? reg13 : reg95) : $unsigned((8'hbe))),
                  (reg89[(3'h4):(3'h4)] < $unsigned((8'had))),
                  $unsigned((&reg67))} ?
              (((reg51 <= reg112) ? ((7'h45) * reg97) : (~reg84)) ?
                  $unsigned(reg67) : reg108) : wire0[(3'h4):(2'h3)]));
      reg117 = reg77[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      if ({($unsigned(($unsigned(wire5) ~^ wire0[(3'h4):(1'h1)])) ?
              {(wire3 ?
                      $unsigned((7'h4b)) : {reg49, reg63})} : ($signed((reg93 ?
                  reg68 : reg20)) <= (reg97 && (wire5 ^~ reg13)))),
          wire1[(5'h12):(3'h7)],
          (8'hb5)})
        begin
          reg118 <= $signed(reg78);
          reg119 = {reg31[(2'h2):(1'h0)]};
          for (forvar120 = (1'h0); (forvar120 < (3'h5)); forvar120 = (forvar120 + (1'h1)))
            begin
              reg121 = $unsigned(reg116);
              reg122 <= reg108;
              reg123 = (((^(reg64 - reg31[(2'h2):(1'h0)])) ?
                  (-{$unsigned(reg58)}) : (reg33[(1'h0):(1'h0)] ?
                      (^~(reg95 >> reg121)) : $unsigned(reg93))) ^ ({(^((8'hae) && (7'h49))),
                  $unsigned((reg64 > (8'hae))),
                  reg67} >= reg97));
              reg124 <= (7'h51);
              reg125 = reg60;
              reg126 <= (8'hab);
            end
        end
      else
        begin
          for (forvar118 = (1'h0); (forvar118 < (2'h3)); forvar118 = (forvar118 + (1'h1)))
            begin
              reg120 <= reg108[(4'hd):(4'hc)];
              reg122 <= (8'hb3);
              reg124 <= (^~$signed(reg49));
              reg125 = {((7'h4a) << wire0[(1'h0):(1'h0)]),
                  reg97[(1'h0):(1'h0)]};
              reg126 <= $signed(wire3[(3'h4):(2'h2)]);
              reg127 <= $unsigned((^~reg114));
              reg128 = ((8'h9e) ?
                  (|({reg116[(5'h12):(4'hf)],
                      {reg105},
                      reg78[(1'h0):(1'h0)]} ^~ ((reg14 ? forvar118 : reg13) ?
                      reg123[(5'h11):(4'h8)] : $signed(reg78)))) : (7'h47));
            end
          reg129 <= $signed(wire5[(4'ha):(3'h4)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar130 = (1'h0); (forvar130 < (3'h5)); forvar130 = (forvar130 + (1'h1)))
        begin
          reg131 = $signed(((|reg67) ?
              {(~&(~^reg18))} : ($unsigned({reg92,
                  reg112}) ^~ $unsigned((!reg98)))));
          reg132 = ((-(|$unsigned((reg131 != reg29)))) ?
              {reg7[(4'hc):(2'h2)],
                  ((8'hae) ^ $unsigned((|reg109)))} : {((&(reg111 ?
                      reg109 : (8'ha1))) + {reg113[(1'h1):(1'h1)],
                      $signed((7'h4c)),
                      (reg47 ^ (7'h47))}),
                  $signed($signed((~&(8'hac)))),
                  ($signed((reg126 << reg29)) ?
                      reg131[(2'h3):(1'h1)] : (^~reg108[(5'h10):(2'h3)]))});
        end
      for (forvar133 = (1'h0); (forvar133 < (2'h2)); forvar133 = (forvar133 + (1'h1)))
        begin
          reg134 <= reg33[(3'h7):(3'h4)];
          reg135 <= $signed($unsigned($signed($unsigned($unsigned(reg37)))));
          reg136 <= ($unsigned((&reg50[(2'h2):(2'h2)])) ?
              {{((reg82 >> reg37) ? (~|reg105) : {reg37}),
                      ($signed(reg89) != (reg114 >>> reg97))},
                  reg84,
                  $unsigned(((8'hb2) ?
                      {reg113} : (reg30 <<< reg131)))} : reg13);
        end
    end
  assign wire137 = reg23;
  always
    @(posedge clk) begin
      reg138 <= (8'hb6);
    end
  assign wire139 = $signed($signed(reg118));
  always
    @(posedge clk) begin
      reg140 <= reg97[(1'h1):(1'h0)];
      reg141 = {reg112};
      reg142 = $unsigned(reg114[(4'hf):(3'h4)]);
      reg143 = ($unsigned(reg114) >= $signed($signed(($unsigned(reg37) == reg32))));
      if (((+(!$unsigned((!reg82)))) < $signed(reg67)))
        begin
          for (forvar144 = (1'h0); (forvar144 < (3'h5)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 <= $signed((reg127[(2'h3):(1'h0)] >= {(|(~|wire137)),
                  reg31}));
              reg146 = (~|$signed((reg95[(5'h1a):(5'h11)] ~^ $signed((wire4 >>> wire139)))));
              reg147 <= reg105;
            end
        end
      else
        begin
          if (reg141[(5'h17):(4'hb)])
            begin
              reg144 <= $unsigned((reg143[(5'h14):(4'hf)] * ({wire4} ?
                  ($signed(reg49) ? reg59 : $signed(wire137)) : reg47)));
              reg145 <= reg50;
              reg146 = (reg105 || reg14);
              reg148 = $signed((~|((~^(!(8'hb5))) ~^ reg105)));
            end
          else
            begin
              reg144 <= $signed((~($signed((~&reg148)) ~^ $unsigned({reg134}))));
              reg145 <= $unsigned(reg20);
            end
          if ({reg95})
            begin
              reg149 = (~(reg102[(3'h4):(1'h1)] << reg134[(4'h8):(3'h7)]));
              reg150 = {($signed((wire137 ~^ reg124[(4'ha):(3'h7)])) < reg134),
                  $signed($signed(($signed(reg97) ~^ ((7'h48) < reg93))))};
              reg151 = $signed((~$signed((-(wire2 != reg148)))));
              reg152 <= $signed((^(8'hb3)));
              reg153 = $signed(reg63[(5'h10):(4'h9)]);
            end
          else
            begin
              reg152 <= ($signed($unsigned(wire0)) && (reg59 ?
                  {reg79, reg129} : ((~&$unsigned((7'h43))) ?
                      ((reg82 ?
                          reg12 : reg116) ^ (7'h57)) : $signed(((7'h4c) ^ reg92)))));
              reg154 <= reg68[(3'h4):(3'h4)];
              reg155 <= reg26[(3'h7):(1'h1)];
            end
          reg156 <= $unsigned(reg152);
          reg157 <= reg64[(5'h10):(1'h1)];
          if (reg145)
            begin
              reg158 = $unsigned((($unsigned({reg155,
                      reg149}) <= $unsigned((-reg68))) ?
                  ({reg97[(2'h2):(1'h0)]} ?
                      ((!reg111) <<< {(8'hb2),
                          reg156}) : reg63) : ($unsigned((reg82 ?
                      (8'hb6) : reg127)) ^ $unsigned($unsigned(reg141)))));
              reg159 = ($signed({(~&(7'h4a)),
                  $signed((reg56 || reg93))}) | $signed({reg63[(5'h16):(2'h3)]}));
              reg160 = reg47;
            end
          else
            begin
              reg158 = $unsigned(reg63);
              reg161 <= (7'h50);
              reg162 = (((reg12[(3'h5):(3'h4)] & reg155[(4'h8):(3'h5)]) > reg68) - $unsigned($unsigned((^~(wire0 ?
                  reg116 : reg156)))));
              reg163 = ((+(^reg92)) | reg141);
            end
        end
      reg164 = reg102;
    end
  assign wire165 = $unsigned(reg152[(4'hd):(4'hb)]);
  assign wire166 = ($signed(($unsigned($signed(reg29)) ?
                       {(|(8'ha5))} : ($signed(reg47) ?
                           (reg26 && (8'hbb)) : reg105[(2'h3):(1'h0)]))) > ($unsigned(reg33) > reg98));
  assign wire167 = {(reg85[(5'h12):(1'h0)] ?
                           $signed(reg51) : reg30[(3'h6):(1'h0)]),
                       reg13[(4'hd):(1'h0)]};
  always
    @(posedge clk) begin
      reg168 <= wire4[(1'h1):(1'h1)];
    end
  assign wire169 = reg95;
  always
    @(posedge clk) begin
      if ({(((8'hb9) >> reg124) >= $unsigned(reg157[(2'h3):(2'h2)]))})
        begin
          if (($unsigned((((^reg126) | (!wire0)) >= reg49[(4'h9):(2'h3)])) < $signed((($unsigned(reg20) ~^ reg156) <<< reg102))))
            begin
              reg170 <= $unsigned((($unsigned((reg152 ? reg29 : wire1)) ?
                      $unsigned(reg140) : ((reg49 >> reg95) ?
                          (~|reg102) : ((8'h9f) ? wire2 : reg111))) ?
                  {(8'hb9),
                      $signed(reg111),
                      ((!reg136) & reg120[(5'h1b):(5'h12)])} : $signed(((reg7 ?
                          reg7 : reg136) ?
                      (reg112 ? reg77 : reg16) : wire3))));
              reg171 <= (~^((reg49[(4'he):(2'h2)] >= reg58[(5'h17):(2'h3)]) ?
                  (reg18[(5'h12):(4'hc)] ?
                      ($unsigned(reg30) ?
                          $signed(reg37) : (~^reg102)) : ({reg140,
                              reg116,
                              reg127} ?
                          reg152[(4'hb):(4'h9)] : (-reg108))) : $unsigned(reg23[(4'hb):(3'h5)])));
              reg172 = {((((!reg14) | (reg68 << (8'hae))) ?
                          reg129[(2'h3):(2'h2)] : $signed(reg147[(1'h0):(1'h0)])) ?
                      $unsigned((|reg67[(4'h9):(2'h2)])) : {(reg108[(5'h10):(4'he)] <<< (|(7'h56))),
                          $unsigned(reg126[(5'h14):(4'hf)]),
                          (^$unsigned(reg40))}),
                  reg26};
              reg173 <= reg147[(4'hb):(1'h1)];
              reg174 <= $unsigned($unsigned($unsigned((reg13 ?
                  reg170[(5'h1a):(5'h11)] : (-reg135)))));
            end
          else
            begin
              reg172 = $signed($unsigned((((reg173 ?
                  reg63 : (8'haa)) && (!reg168)) >>> wire3[(3'h4):(3'h4)])));
              reg175 = reg93[(2'h2):(1'h0)];
              reg176 <= reg49;
              reg177 = (8'hb5);
              reg178 = (+(~$signed($unsigned(wire4))));
            end
          reg179 = $signed($signed(reg112));
          for (forvar180 = (1'h0); (forvar180 < (3'h4)); forvar180 = (forvar180 + (1'h1)))
            begin
              reg181 = reg63[(4'hb):(3'h6)];
              reg182 <= (8'h9f);
              reg183 <= reg7;
              reg184 = (({$signed((reg22 - reg108)),
                  ({reg140} ?
                      (reg16 + reg181) : reg7[(2'h2):(1'h0)])} <= {{reg56[(2'h2):(1'h1)],
                      $unsigned(reg173),
                      reg47[(2'h3):(2'h3)]},
                  reg30[(4'h8):(3'h7)],
                  $signed(wire5[(3'h7):(3'h7)])}) <<< wire165[(4'hd):(3'h6)]);
            end
          reg185 = $unsigned((forvar180[(4'hb):(4'ha)] >>> reg179[(3'h5):(1'h0)]));
          reg186 <= (!reg56[(2'h2):(1'h0)]);
          reg187 = reg178;
          reg188 = (|{reg183});
        end
      else
        begin
          if (($signed(reg172) && $unsigned(wire4)))
            begin
              reg172 = (~|(reg92[(3'h7):(1'h0)] ?
                  reg184[(4'ha):(3'h6)] : reg188[(5'h10):(1'h0)]));
              reg175 = {(-($signed(reg173) ?
                      reg177[(4'h9):(1'h0)] : {reg155[(1'h1):(1'h1)],
                          {reg188, reg79, reg32}})),
                  ($signed($signed({reg40, reg175})) ?
                      $unsigned(((reg176 ?
                          reg7 : reg147) << reg47[(4'h8):(2'h3)])) : wire165[(1'h1):(1'h1)]),
                  ($unsigned($signed((reg187 == forvar180))) ?
                      (^(!$signed(reg114))) : {({reg59, reg186, reg49} ?
                              (^forvar180) : reg58[(4'hb):(4'h8)]),
                          (reg179[(2'h2):(2'h2)] >= ((7'h48) ?
                              reg126 : (8'haa)))})};
              reg176 <= (+$unsigned((reg156 ?
                  {reg175[(3'h5):(2'h3)],
                      {reg178, (8'h9c), wire0},
                      ((8'hbd) ? (7'h47) : (8'hb0))} : ((7'h47) ?
                      $signed(reg116) : (+reg183)))));
              reg180 <= $unsigned($signed(reg77));
              reg181 = reg173;
              reg182 <= $signed(($signed($unsigned({reg127,
                  reg49,
                  wire3})) + reg89));
            end
          else
            begin
              reg172 = (reg42[(4'hd):(3'h6)] <<< (&reg126));
              reg175 = ($unsigned(((reg120 && $signed(reg67)) != $unsigned(reg173[(1'h1):(1'h0)]))) ?
                  (({{reg134, reg134}} < wire169[(2'h2):(1'h0)]) ?
                      reg89 : (((&reg109) >> (reg67 - reg92)) ?
                          ((reg183 | wire3) ?
                              $signed((8'hae)) : reg177[(3'h7):(3'h7)]) : reg32)) : (reg56 | $unsigned(((~reg23) ?
                      (reg180 <= reg84) : reg31[(1'h0):(1'h0)]))));
            end
        end
    end
  module189 #() modinst1775 (.wire190(reg168), .wire191(reg56), .y(wire1774), .wire195(reg116), .wire193(reg42), .wire194(reg114), .wire192(reg174), .clk(clk));
  assign wire1776 = $signed(($signed(reg182[(3'h4):(1'h0)]) ~^ $unsigned(reg29[(3'h4):(3'h4)])));
  always
    @(posedge clk) begin
      for (forvar1777 = (1'h0); (forvar1777 < (2'h3)); forvar1777 = (forvar1777 + (1'h1)))
        begin
          for (forvar1778 = (1'h0); (forvar1778 < (2'h2)); forvar1778 = (forvar1778 + (1'h1)))
            begin
              reg1779 = $signed((reg180[(4'hc):(2'h3)] >= reg183[(4'hb):(4'ha)]));
              reg1780 <= (-$signed($signed(($signed(forvar1777) | (reg127 ?
                  reg124 : reg60)))));
            end
          reg1781 = ($unsigned({$unsigned($signed(reg47))}) & {$signed((^~$unsigned(wire167)))});
          reg1782 = reg108[(2'h3):(1'h1)];
          reg1783 <= {(reg105 ?
                  ((forvar1777[(5'h13):(3'h6)] ?
                          $unsigned(forvar1778) : (reg67 ? reg37 : reg182)) ?
                      reg170[(4'he):(4'he)] : ((8'ha7) ?
                          $signed((8'hb9)) : (~^reg138))) : reg126),
              wire166};
          reg1784 <= $unsigned($unsigned(wire1[(5'h16):(2'h3)]));
          reg1785 = (^$signed(reg155));
        end
      reg1786 = ((7'h47) ? reg1783[(5'h10):(4'hc)] : reg126);
      reg1787 <= reg7[(1'h0):(1'h0)];
      if ((8'ha1))
        begin
          reg1788 = {$unsigned($signed(reg64)), ((7'h4b) >> reg186)};
          reg1789 = reg157;
          reg1790 = (reg176 * ($unsigned(reg68) >> $unsigned($unsigned($unsigned(reg40)))));
          if ($unsigned(reg180))
            begin
              reg1791 = $unsigned((((|(|reg161)) >>> ($unsigned(reg113) ?
                  $unsigned(reg124) : (reg122 + reg111))) || $signed($unsigned(wire137[(4'ha):(2'h2)]))));
              reg1792 <= $unsigned($signed(reg183[(4'he):(4'he)]));
              reg1793 <= (^reg127);
              reg1794 = (|(!$unsigned(reg26)));
              reg1795 <= ((+(^~$unsigned(reg127))) ?
                  reg49[(5'h12):(4'hb)] : reg1789);
              reg1796 <= $signed((&((8'h9f) ?
                  ({wire166} ? (7'h53) : $unsigned(reg29)) : reg168)));
            end
          else
            begin
              reg1791 = reg14;
              reg1794 = $signed((+reg63));
              reg1795 <= (reg26[(3'h7):(2'h2)] ?
                  {($unsigned((8'ha4)) != (&(8'ha8))),
                      $signed((~(wire167 ?
                          reg134 : reg58)))} : $unsigned($signed(reg122[(5'h17):(3'h6)])));
              reg1797 = (reg116[(5'h16):(3'h6)] ~^ (~({$unsigned(reg122)} ?
                  (-$signed(reg51)) : (~&wire4[(4'h9):(3'h4)]))));
              reg1798 <= $unsigned(reg112);
            end
          for (forvar1799 = (1'h0); (forvar1799 < (2'h3)); forvar1799 = (forvar1799 + (1'h1)))
            begin
              reg1800 = reg33;
              reg1801 <= ($signed(reg59) ?
                  $unsigned($signed(reg42[(3'h6):(1'h0)])) : (reg59[(4'ha):(4'h9)] * reg118));
              reg1802 = (~^((|(^reg1793)) <= (((reg1800 ?
                  (7'h50) : reg135) >> (!reg129)) | ($signed(reg174) <= reg108))));
            end
        end
      else
        begin
          reg1792 <= reg1781;
          if (($unsigned({$unsigned($unsigned(reg97))}) ^ reg32))
            begin
              reg1794 = $signed(wire137[(5'h14):(4'he)]);
              reg1797 = reg1793[(5'h13):(4'h8)];
            end
          else
            begin
              reg1793 <= {{((reg1802[(4'hd):(1'h1)] ?
                              $unsigned(reg129) : (reg118 && reg102)) ?
                          reg140[(1'h1):(1'h0)] : (reg176 - (reg140 != reg1790))),
                      reg109,
                      (reg1789 >>> reg116)}};
              reg1794 = reg1798;
              reg1795 <= $signed((+reg67[(1'h1):(1'h1)]));
              reg1797 = reg63[(4'h9):(1'h0)];
              reg1799 = ((reg95[(4'hf):(4'h8)] >>> reg147[(3'h5):(1'h1)]) & ({($unsigned(reg155) ~^ reg84[(4'hb):(3'h7)]),
                  ((^~reg1780) ? (!reg129) : $unsigned(wire166)),
                  ((reg1788 << (7'h4f)) + $unsigned(reg180))} >= reg84[(4'h9):(3'h7)]));
            end
          if (reg29)
            begin
              reg1800 = $unsigned({$unsigned((reg50[(3'h5):(2'h3)] || (reg113 == reg118)))});
              reg1801 <= $unsigned($unsigned($signed($signed($signed(reg118)))));
              reg1802 = reg84;
              reg1803 = (reg60[(4'h9):(3'h4)] != ((reg1782 >= ((-reg1787) ?
                  $signed(reg18) : ((7'h50) ? reg105 : (7'h4e)))) << reg40));
            end
          else
            begin
              reg1800 = (^(~(8'hb4)));
              reg1802 = reg22;
              reg1803 = ((~&((reg82 - (reg156 > reg113)) <= ((^~reg29) ?
                      $unsigned(reg14) : (reg85 ^~ reg50)))) ?
                  (7'h50) : $unsigned(($signed($unsigned(reg145)) ?
                      reg49 : ($unsigned((8'hb0)) | $unsigned(reg136)))));
              reg1804 <= ($signed({$unsigned(reg1797[(4'hd):(4'hd)])}) ?
                  reg156 : reg1794[(4'hb):(2'h2)]);
              reg1805 = wire167;
              reg1806 <= $unsigned($signed($unsigned((((8'hb9) ?
                      reg1783 : reg59) ?
                  (~&reg12) : $unsigned(reg42)))));
              reg1807 = $unsigned({(reg113[(5'h12):(3'h7)] != {{(8'haf),
                          wire167,
                          reg156},
                      (reg1804 | reg144),
                      {wire167, reg144, reg120}}),
                  (!reg26[(4'h9):(3'h6)]),
                  (7'h45)});
            end
          reg1808 <= reg22;
          for (forvar1809 = (1'h0); (forvar1809 < (3'h4)); forvar1809 = (forvar1809 + (1'h1)))
            begin
              reg1810 <= (^(^(~^((+reg1795) ?
                  (|reg1808) : $unsigned(reg1807)))));
              reg1811 = $signed($signed($unsigned(((reg42 || reg152) - reg49[(2'h2):(1'h1)]))));
              reg1812 <= ((reg1806 >= ($signed((forvar1809 ?
                  (8'hb3) : reg1795)) | reg113[(3'h4):(1'h1)])) ^ (8'ha3));
              reg1813 <= $signed(((~^((reg51 ? reg174 : reg173) ?
                  $unsigned(reg152) : reg85)) * ((!((7'h56) != reg84)) ?
                  reg1799 : (^~reg126))));
              reg1814 = $unsigned((reg1802[(3'h7):(3'h5)] << (|reg129[(3'h5):(1'h0)])));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1815 = (1'h0); (forvar1815 < (2'h3)); forvar1815 = (forvar1815 + (1'h1)))
        begin
          for (forvar1816 = (1'h0); (forvar1816 < (2'h3)); forvar1816 = (forvar1816 + (1'h1)))
            begin
              reg1817 = (8'hb5);
              reg1818 = (-((reg60[(4'h9):(2'h3)] ?
                  (8'hba) : $signed($signed(reg49))) > reg1798[(4'hd):(4'hd)]));
              reg1819 = reg135;
              reg1820 = {(reg136[(1'h0):(1'h0)] ?
                      (reg1783[(4'h9):(2'h2)] ^ (^{(7'h45),
                          reg64})) : {{$signed((8'hb9)),
                              reg136[(3'h4):(2'h3)],
                              $signed(reg1801)},
                          reg120[(5'h19):(3'h4)]})};
              reg1821 = (+$signed((&$signed(wire1774))));
              reg1822 <= (~^(^($signed(reg1801[(4'he):(4'hc)]) || $unsigned((-reg78)))));
            end
          for (forvar1823 = (1'h0); (forvar1823 < (1'h1)); forvar1823 = (forvar1823 + (1'h1)))
            begin
              reg1824 = ((+$unsigned($signed((reg1793 >>> reg173)))) != (reg173 != (~reg140[(2'h2):(1'h0)])));
              reg1825 <= (^((~{$signed(reg95),
                  (&(7'h42)),
                  $unsigned(reg1817)}) < reg56));
              reg1826 = reg31;
              reg1827 = (~&$unsigned(reg16[(3'h4):(1'h0)]));
              reg1828 = ($unsigned((!$unsigned((^reg20)))) ?
                  (((-(reg80 + reg23)) ?
                      (!$signed(reg67)) : $unsigned($unsigned(reg157))) == $unsigned(reg1810[(4'hb):(4'hb)])) : reg64[(4'hc):(2'h3)]);
            end
          reg1829 = reg168[(1'h1):(1'h1)];
          reg1830 <= $unsigned(($signed(wire169[(1'h0):(1'h0)]) ?
              (~&$unsigned((+wire1776))) : (reg89 >> (reg85[(4'hf):(4'h8)] ?
                  (wire139 <<< forvar1815) : (reg92 ^ reg1795)))));
        end
    end
  assign wire1831 = $signed(($unsigned($signed($signed(wire1776))) ?
                        (|wire1[(1'h0):(1'h0)]) : reg1810));
  always
    @(posedge clk) begin
      for (forvar1832 = (1'h0); (forvar1832 < (3'h4)); forvar1832 = (forvar1832 + (1'h1)))
        begin
          reg1833 = reg51;
          if (reg108)
            begin
              reg1834 <= {(((wire1 && reg135) >= (~^$signed(reg1792))) ?
                      reg80[(5'h10):(3'h4)] : {$unsigned($signed(reg182)),
                          {reg112, reg176}})};
              reg1835 = (^~{$unsigned((&(reg145 ? reg1793 : reg47))), reg183});
              reg1836 = {reg161, $unsigned((~{$unsigned((8'ha3)), reg78}))};
              reg1837 = (+reg109);
              reg1838 <= (7'h57);
              reg1839 = $signed({$unsigned((wire0[(1'h1):(1'h0)] ?
                      reg98[(3'h5):(2'h2)] : wire1[(5'h1a):(3'h7)])),
                  $unsigned($unsigned(wire137))});
              reg1840 = reg136;
            end
          else
            begin
              reg1834 <= reg138;
              reg1838 <= ((-$unsigned((+$unsigned(reg50)))) ?
                  reg68[(2'h2):(1'h1)] : $unsigned({$unsigned(reg68)}));
              reg1839 = reg112[(5'h10):(5'h10)];
              reg1840 = reg155;
            end
          reg1841 = ($signed(($unsigned(reg1793) ?
                  (~(reg1801 ? reg98 : reg138)) : reg18[(5'h1d):(4'ha)])) ?
              (((~^reg30[(4'hc):(1'h0)]) ?
                  {{(7'h51)}} : ((!reg145) > reg112)) ~^ (({wire1774} ?
                      $unsigned(reg29) : (~|reg108)) ?
                  ((|reg1784) ?
                      $signed((8'ha1)) : (^(8'hb7))) : ($signed(wire0) == $unsigned((7'h47))))) : ((~$signed((reg84 * (8'hae)))) ?
                  reg144 : reg186[(5'h15):(5'h15)]));
          for (forvar1842 = (1'h0); (forvar1842 < (2'h3)); forvar1842 = (forvar1842 + (1'h1)))
            begin
              reg1843 = ($signed((reg18 ?
                  reg84[(4'hd):(4'hd)] : reg108[(5'h10):(2'h3)])) <<< reg1838);
              reg1844 <= $unsigned($unsigned(($unsigned($unsigned(reg170)) >>> (~|reg92[(4'h8):(3'h4)]))));
              reg1845 = (reg51[(3'h4):(1'h1)] << {reg145});
            end
          reg1846 = ((reg1844 > (($signed(reg183) ?
              $signed(wire137) : reg1841[(1'h0):(1'h0)]) * reg56)) && ((~|({forvar1842} ?
                  reg118[(3'h5):(1'h1)] : (reg1841 && reg84))) ?
              $signed((reg1830[(1'h1):(1'h0)] <= $unsigned(wire4))) : ($signed((^(7'h54))) ?
                  $unsigned((reg51 ^ wire0)) : ((&reg84) == $signed(reg26)))));
          if (reg116)
            begin
              reg1847 <= reg186[(5'h1c):(5'h13)];
            end
          else
            begin
              reg1848 = (~|$unsigned(reg7[(3'h4):(1'h0)]));
              reg1849 = reg68;
              reg1850 = ((-$signed(wire2[(4'h8):(4'h8)])) >> ($signed({reg22[(5'h17):(1'h0)],
                  (reg174 & reg186)}) < $signed(($unsigned(reg1830) > (~reg82)))));
              reg1851 <= reg176[(5'h14):(3'h7)];
              reg1852 <= reg33;
            end
        end
      reg1853 = $signed(wire1774);
      reg1854 = $signed($unsigned(reg82[(2'h3):(2'h3)]));
      if ((^~(~&$signed(((reg135 ? reg56 : reg82) ?
          reg14[(1'h0):(1'h0)] : (+reg145))))))
        begin
          reg1855 = reg176[(5'h12):(5'h12)];
        end
      else
        begin
          reg1855 = (~&($unsigned((^~(~|reg89))) ?
              reg109[(3'h7):(1'h1)] : $signed(reg145[(4'ha):(4'ha)])));
          reg1856 <= reg84;
          reg1857 <= (~|($signed((^~(reg59 ? reg1846 : reg78))) ?
              reg154 : $unsigned((7'h4f))));
        end
      reg1858 = (reg79[(1'h1):(1'h1)] * (reg47 ?
          $unsigned((reg186[(5'h13):(3'h5)] >>> $unsigned((7'h55)))) : ((^~$unsigned(reg20)) && reg1822[(4'he):(3'h4)])));
      for (forvar1859 = (1'h0); (forvar1859 < (2'h2)); forvar1859 = (forvar1859 + (1'h1)))
        begin
          if (reg7[(3'h4):(1'h0)])
            begin
              reg1860 <= ((~&reg180) ?
                  $signed($unsigned((^~$signed(reg118)))) : {($signed(((8'h9f) * reg1855)) ?
                          $unsigned(((7'h4c) ? reg1849 : reg176)) : (+(reg59 ?
                              reg1804 : reg1853))),
                      ($unsigned($signed(reg49)) ?
                          wire3[(3'h5):(2'h3)] : $unsigned((~|reg59)))});
              reg1861 <= $signed(reg155[(2'h3):(2'h2)]);
              reg1862 = $signed($signed(($unsigned($signed(reg1841)) & ($signed(reg51) != {reg155,
                  reg1806,
                  reg124}))));
            end
          else
            begin
              reg1862 = ({{($signed(reg1848) ?
                          $signed(reg1847) : $signed(reg31))},
                  $unsigned((reg42[(5'h1d):(5'h16)] && reg1830))} || reg78);
              reg1863 <= reg1840[(5'h1a):(4'h9)];
              reg1864 <= (reg1852[(1'h1):(1'h0)] ^ (((^~$signed((8'hb4))) ?
                  {(~reg1810),
                      (reg16 ?
                          reg1833 : reg1858)} : (8'ha8)) - (reg1849[(5'h14):(5'h10)] >>> {$unsigned(reg1855),
                  $signed((8'hb8))})));
              reg1865 <= ({$unsigned($unsigned((~&reg1798)))} ?
                  (|($signed(reg105) ^~ ((|reg1850) ?
                      ((7'h48) ? reg14 : reg1808) : reg58))) : reg109);
              reg1866 <= reg111;
              reg1867 = reg124;
              reg1868 = reg145;
            end
          if ((({reg109,
              forvar1832} * $signed((reg67[(3'h4):(2'h3)] && $signed(reg113)))) + reg1783[(1'h0):(1'h0)]))
            begin
              reg1869 <= $signed({(8'hb5),
                  {(^~$signed(reg1846)),
                      $signed((reg168 >>> reg20)),
                      $signed((reg144 ? reg152 : wire0))}});
            end
          else
            begin
              reg1870 = (~&(reg32[(3'h4):(3'h4)] ?
                  (-(reg155 ^ $signed(reg1864))) : $signed(reg1783[(5'h10):(4'hf)])));
              reg1871 = ({(($signed(reg68) ?
                          $unsigned(wire166) : reg111[(3'h7):(3'h4)]) >>> ($signed(reg89) ?
                          $unsigned((8'hb0)) : $unsigned(reg1804))),
                      reg127[(5'h13):(2'h2)]} ?
                  ((|reg1865[(4'h9):(3'h4)]) <= ($unsigned({reg1869,
                          reg168,
                          reg180}) ?
                      reg1813[(4'h9):(3'h6)] : reg1865[(2'h2):(1'h1)])) : (-($signed((^~reg78)) >= (+reg29[(5'h14):(2'h3)]))));
              reg1872 <= reg67[(3'h4):(1'h0)];
              reg1873 = reg1795;
              reg1874 <= ((((+((8'hbd) ? reg120 : (7'h51))) ?
                  $unsigned({(7'h55), reg152, reg108}) : {((8'hb3) ^ reg23),
                      (!reg1857)}) | $signed((~|(wire167 >> wire1)))) & reg1858[(1'h1):(1'h0)]);
              reg1875 = $signed($unsigned({reg174[(4'h9):(1'h1)],
                  reg127[(5'h11):(2'h3)]}));
            end
          reg1876 = $signed(($signed((reg1850[(1'h1):(1'h0)] ^~ (+reg1857))) ?
              ($unsigned((~^reg1796)) - (reg47[(4'ha):(2'h3)] + (reg92 <<< reg37))) : (($unsigned((8'ha1)) ?
                      $signed(reg118) : reg135) ?
                  ((8'ha4) <<< {reg50,
                      reg168,
                      (7'h56)}) : reg1851[(3'h5):(1'h0)])));
          if ($signed((-((wire137[(5'h19):(5'h17)] ? (-reg1810) : (&reg1863)) ?
              (!reg1850[(4'h8):(2'h3)]) : (|forvar1842[(2'h3):(2'h2)])))))
            begin
              reg1877 = $unsigned(($signed(reg79) ?
                  $signed(wire169[(3'h7):(1'h0)]) : reg1796[(3'h5):(3'h5)]));
              reg1878 = $signed((~|$unsigned(($signed(reg129) ?
                  wire0 : $unsigned(reg1876)))));
              reg1879 = ($unsigned(((reg1877 ?
                  $unsigned(reg1796) : reg93[(5'h1a):(3'h7)]) * wire1)) || (reg1837 + ($signed((^reg145)) ?
                  reg1857[(1'h1):(1'h1)] : ((reg171 >>> reg176) * reg127[(3'h6):(3'h6)]))));
              reg1880 = $unsigned(($signed(reg23) ?
                  reg1846[(3'h6):(1'h0)] : (|$unsigned($signed(reg58)))));
              reg1881 = (($unsigned($signed((reg56 ^ reg108))) ^ {(!((8'hb0) ?
                          reg1806 : reg112)),
                      reg1863}) ?
                  reg14 : $unsigned(reg50));
              reg1882 <= wire165[(5'h1d):(5'h14)];
            end
          else
            begin
              reg1882 <= (&{($signed($signed(reg89)) && reg89[(3'h5):(3'h4)]),
                  ((reg1879 || reg1812) ?
                      (reg1801[(5'h17):(5'h14)] ?
                          $signed(reg85) : (reg140 ?
                              (7'h40) : reg1875)) : $signed((~reg51)))});
              reg1883 <= $signed($unsigned(($signed((^reg1874)) ?
                  $unsigned($signed((7'h46))) : (reg1812 ?
                      (|reg155) : (+reg1801)))));
              reg1884 <= reg1796;
              reg1885 <= reg120;
              reg1886 <= $unsigned(({{(~^reg174), {reg1840, reg109}},
                  reg1793[(4'hf):(4'he)],
                  reg113[(3'h4):(2'h3)]} >> (!($unsigned(reg1839) >= reg89))));
              reg1887 <= $unsigned(reg33);
              reg1888 = $unsigned((^~reg40));
            end
          if (reg102[(1'h0):(1'h0)])
            begin
              reg1889 = reg1862;
              reg1890 <= ({((reg1834[(5'h12):(5'h12)] || (^wire4)) ?
                      $unsigned({(8'hb1), reg157, reg1887}) : wire1),
                  $signed({(|reg98),
                      (forvar1832 ? reg155 : reg1810),
                      reg16})} ^ (wire5[(4'hf):(4'h8)] ?
                  reg78[(3'h5):(3'h4)] : {(((8'ha4) ?
                          reg1848 : reg1867) <<< reg26[(4'hc):(4'h9)]),
                      reg1813,
                      $unsigned((&reg182))}));
            end
          else
            begin
              reg1889 = $unsigned($unsigned($unsigned(($signed(reg1848) * (reg1854 ?
                  reg183 : reg171)))));
              reg1891 = $unsigned(($unsigned($signed($unsigned(reg26))) ?
                  $signed({reg136,
                      $unsigned(reg1871),
                      (+reg64)}) : {reg30[(2'h3):(2'h3)],
                      $signed((reg92 ? reg56 : (8'hb3)))}));
              reg1892 <= {(reg1834[(1'h1):(1'h1)] >= reg1796),
                  reg1858,
                  reg168[(1'h0):(1'h0)]};
            end
        end
      for (forvar1893 = (1'h0); (forvar1893 < (2'h2)); forvar1893 = (forvar1893 + (1'h1)))
        begin
          reg1894 <= $unsigned((|(+reg1835[(3'h4):(1'h0)])));
          if (($signed(((7'h54) ?
                  ($signed(reg37) >= forvar1859) : ((~^reg124) ?
                      {(8'ha3), (8'hb9), reg1873} : (reg174 ?
                          (7'h45) : reg1892)))) ?
              wire5 : reg1873[(5'h12):(4'hb)]))
            begin
              reg1895 = (-(~(^$signed($unsigned(reg182)))));
              reg1896 = $signed((reg97 ?
                  ((&$unsigned(reg1845)) <= $signed($unsigned((7'h44)))) : reg64));
            end
          else
            begin
              reg1895 = $unsigned($unsigned($unsigned({$signed((8'hbf)),
                  (wire2 ? reg1808 : reg1849),
                  $signed(reg1836)})));
              reg1896 = $unsigned(reg1896);
            end
          reg1897 = (^$unsigned((reg174 >>> (wire1776 ?
              reg170[(5'h12):(4'hc)] : $unsigned(wire166)))));
          for (forvar1898 = (1'h0); (forvar1898 < (3'h6)); forvar1898 = (forvar1898 + (1'h1)))
            begin
              reg1899 = reg68[(2'h2):(1'h0)];
            end
        end
    end
  module1005 #() modinst1901 (.wire1007(reg1813), .wire1008(reg180), .wire1006(reg1804), .wire1009(reg152), .clk(clk), .y(wire1900), .wire1010(reg1865));
  module1005 #() modinst1903 (wire1902, clk, reg18, reg1890, reg1795, reg102, reg26);
  module189 #() modinst1905 (wire1904, clk, reg1834, reg29, reg64, reg1796, reg114, wire166);
  assign wire1906 = $unsigned(($unsigned((!(~|(8'hb6)))) ?
                        $signed(((wire2 != reg114) && $signed(reg98))) : reg1780[(4'ha):(4'ha)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module189
#(parameter param1773 = ((|{{(&(7'h58)), (&(8'hbd)), ((8'h9f) && (8'hba))}}) > (((~|(8'hae)) + ((^(7'h51)) ? ((8'hbb) ? (7'h52) : (8'ha4)) : ((8'hbb) ? (8'h9f) : (7'h4f)))) || ((((8'hbc) ? (8'hbd) : (7'h4e)) ? ((7'h4c) != (7'h51)) : (7'h40)) ? (((8'ha7) * (7'h55)) ? (!(7'h4c)) : ((8'h9f) ~^ (8'hb2))) : (((8'ha6) != (8'ha5)) ? (~(7'h54)) : ((8'hbd) ? (8'hbb) : (8'ha2)))))))
(y, clk, wire195, wire194, wire193, wire192, wire191, wire190);
  output wire [(32'h3be2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire195;
  input wire [(5'h17):(1'h0)] wire194;
  input wire signed [(5'h17):(1'h0)] wire193;
  input wire signed [(2'h3):(1'h0)] wire192;
  input wire [(5'h10):(1'h0)] wire191;
  input wire signed [(4'hb):(1'h0)] wire190;
  wire signed [(4'h9):(1'h0)] wire1772;
  wire signed [(5'h15):(1'h0)] wire1739;
  wire signed [(4'h9):(1'h0)] wire1697;
  wire [(5'h19):(1'h0)] wire1613;
  wire signed [(5'h19):(1'h0)] wire1494;
  wire signed [(4'hb):(1'h0)] wire754;
  wire [(5'h14):(1'h0)] wire718;
  wire [(5'h17):(1'h0)] wire717;
  wire [(4'hc):(1'h0)] wire584;
  wire [(5'h17):(1'h0)] wire516;
  wire signed [(5'h18):(1'h0)] wire351;
  wire [(5'h10):(1'h0)] wire350;
  reg [(4'he):(1'h0)] reg1770 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1762 = (1'h0);
  reg [(5'h13):(1'h0)] reg1761 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1757 = (1'h0);
  reg [(3'h5):(1'h0)] reg1755 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1753 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1752 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1747 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1744 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1742 = (1'h0);
  reg [(4'h8):(1'h0)] reg1741 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1740 = (1'h0);
  reg [(5'h14):(1'h0)] reg1738 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1728 = (1'h0);
  reg [(5'h17):(1'h0)] reg1734 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1733 = (1'h0);
  reg [(4'hf):(1'h0)] reg1732 = (1'h0);
  reg [(4'hb):(1'h0)] reg1731 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1726 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1725 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1724 = (1'h0);
  reg [(2'h2):(1'h0)] reg1722 = (1'h0);
  reg [(5'h13):(1'h0)] reg1721 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1719 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1717 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1714 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1712 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1708 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1705 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1700 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1696 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1695 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1694 = (1'h0);
  reg [(4'h9):(1'h0)] reg1690 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1688 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1686 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1683 = (1'h0);
  reg [(3'h6):(1'h0)] reg1680 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1679 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1677 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1675 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1673 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1671 = (1'h0);
  reg [(3'h7):(1'h0)] reg1670 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1668 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1665 = (1'h0);
  reg [(4'hf):(1'h0)] reg1664 = (1'h0);
  reg [(5'h17):(1'h0)] reg1658 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1657 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1655 = (1'h0);
  reg [(4'hf):(1'h0)] reg1654 = (1'h0);
  reg [(4'he):(1'h0)] reg1651 = (1'h0);
  reg [(3'h5):(1'h0)] reg1649 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1647 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1646 = (1'h0);
  reg [(3'h4):(1'h0)] reg1644 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1643 = (1'h0);
  reg [(5'h10):(1'h0)] reg1637 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1636 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1632 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1627 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1621 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1620 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1618 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1617 = (1'h0);
  reg [(4'hc):(1'h0)] reg1615 = (1'h0);
  reg [(5'h17):(1'h0)] reg1614 = (1'h0);
  reg [(4'he):(1'h0)] reg1612 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1610 = (1'h0);
  reg [(3'h5):(1'h0)] reg1609 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1607 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1606 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1605 = (1'h0);
  reg [(5'h13):(1'h0)] reg1604 = (1'h0);
  reg [(2'h3):(1'h0)] reg1603 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1600 = (1'h0);
  reg [(5'h13):(1'h0)] reg1599 = (1'h0);
  reg [(3'h6):(1'h0)] reg1598 = (1'h0);
  reg [(2'h2):(1'h0)] reg1596 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1594 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1591 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1589 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1587 = (1'h0);
  reg [(5'h18):(1'h0)] reg1586 = (1'h0);
  reg [(5'h17):(1'h0)] reg1584 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1583 = (1'h0);
  reg [(4'hb):(1'h0)] reg1580 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1578 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1577 = (1'h0);
  reg [(5'h13):(1'h0)] reg1576 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1575 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1572 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1571 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1566 = (1'h0);
  reg [(5'h18):(1'h0)] reg1563 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1562 = (1'h0);
  reg [(3'h4):(1'h0)] reg1560 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1559 = (1'h0);
  reg [(4'hd):(1'h0)] reg1558 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1555 = (1'h0);
  reg [(5'h11):(1'h0)] reg1554 = (1'h0);
  reg [(3'h5):(1'h0)] reg1552 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1551 = (1'h0);
  reg [(3'h6):(1'h0)] reg1550 = (1'h0);
  reg [(3'h6):(1'h0)] reg1549 = (1'h0);
  reg [(5'h18):(1'h0)] reg1548 = (1'h0);
  reg [(4'hc):(1'h0)] reg1544 = (1'h0);
  reg [(4'h8):(1'h0)] reg1539 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1537 = (1'h0);
  reg [(4'ha):(1'h0)] reg1534 = (1'h0);
  reg [(5'h12):(1'h0)] reg1533 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1532 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1529 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1528 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1527 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1525 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1524 = (1'h0);
  reg [(3'h6):(1'h0)] reg1523 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1514 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1517 = (1'h0);
  reg [(4'hf):(1'h0)] reg1516 = (1'h0);
  reg [(5'h16):(1'h0)] reg1508 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1507 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1501 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1500 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1497 = (1'h0);
  reg [(4'he):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg892 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg891 = (1'h0);
  reg [(5'h1e):(1'h0)] reg889 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg884 = (1'h0);
  reg [(4'he):(1'h0)] reg881 = (1'h0);
  reg [(2'h3):(1'h0)] reg880 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg879 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg878 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg874 = (1'h0);
  reg [(3'h4):(1'h0)] reg872 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg871 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg870 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg866 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg863 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg859 = (1'h0);
  reg [(5'h11):(1'h0)] reg858 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg856 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg847 = (1'h0);
  reg signed [(4'he):(1'h0)] reg853 = (1'h0);
  reg [(3'h7):(1'h0)] reg850 = (1'h0);
  reg [(5'h12):(1'h0)] reg849 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg844 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg842 = (1'h0);
  reg [(4'he):(1'h0)] reg841 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg839 = (1'h0);
  reg [(5'h10):(1'h0)] reg837 = (1'h0);
  reg [(5'h1f):(1'h0)] reg818 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg834 = (1'h0);
  reg [(5'h16):(1'h0)] reg833 = (1'h0);
  reg [(5'h1f):(1'h0)] reg832 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg828 = (1'h0);
  reg [(4'hb):(1'h0)] reg827 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg815 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg813 = (1'h0);
  reg [(5'h1b):(1'h0)] reg811 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg810 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg809 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg808 = (1'h0);
  reg [(4'hc):(1'h0)] reg805 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg803 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg801 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg798 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg796 = (1'h0);
  reg [(5'h1c):(1'h0)] reg795 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg793 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg790 = (1'h0);
  reg [(5'h1d):(1'h0)] reg789 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg787 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg785 = (1'h0);
  reg [(5'h14):(1'h0)] reg783 = (1'h0);
  reg [(5'h1a):(1'h0)] reg782 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg779 = (1'h0);
  reg [(5'h11):(1'h0)] reg778 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg776 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg775 = (1'h0);
  reg [(5'h13):(1'h0)] reg774 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg773 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg769 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg767 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg763 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg762 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg760 = (1'h0);
  reg signed [(4'he):(1'h0)] reg757 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg750 = (1'h0);
  reg [(4'h8):(1'h0)] reg747 = (1'h0);
  reg [(4'h8):(1'h0)] reg745 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg744 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg742 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg741 = (1'h0);
  reg [(4'ha):(1'h0)] reg736 = (1'h0);
  reg [(5'h1a):(1'h0)] reg734 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg731 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg730 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg728 = (1'h0);
  reg [(4'h9):(1'h0)] reg727 = (1'h0);
  reg [(5'h1c):(1'h0)] reg726 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg713 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg709 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg708 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg707 = (1'h0);
  reg signed [(4'he):(1'h0)] reg705 = (1'h0);
  reg [(5'h16):(1'h0)] reg704 = (1'h0);
  reg [(3'h5):(1'h0)] reg703 = (1'h0);
  reg [(4'h8):(1'h0)] reg702 = (1'h0);
  reg [(3'h7):(1'h0)] reg700 = (1'h0);
  reg [(5'h13):(1'h0)] reg699 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg698 = (1'h0);
  reg [(4'hc):(1'h0)] reg696 = (1'h0);
  reg [(5'h11):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg689 = (1'h0);
  reg [(5'h10):(1'h0)] reg688 = (1'h0);
  reg [(5'h13):(1'h0)] reg683 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg678 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg675 = (1'h0);
  reg signed [(4'he):(1'h0)] reg674 = (1'h0);
  reg [(4'hd):(1'h0)] reg673 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg672 = (1'h0);
  reg [(4'hd):(1'h0)] reg671 = (1'h0);
  reg [(5'h16):(1'h0)] reg669 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg664 = (1'h0);
  reg [(4'h8):(1'h0)] reg663 = (1'h0);
  reg [(5'h11):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg657 = (1'h0);
  reg [(2'h2):(1'h0)] reg655 = (1'h0);
  reg [(3'h4):(1'h0)] reg654 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg653 = (1'h0);
  reg [(5'h13):(1'h0)] reg652 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg650 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg649 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg648 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg646 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg645 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg643 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg641 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg639 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg636 = (1'h0);
  reg [(4'h8):(1'h0)] reg635 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg634 = (1'h0);
  reg [(3'h7):(1'h0)] reg627 = (1'h0);
  reg [(5'h15):(1'h0)] reg624 = (1'h0);
  reg [(4'h8):(1'h0)] reg620 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg619 = (1'h0);
  reg [(4'he):(1'h0)] reg618 = (1'h0);
  reg [(4'h9):(1'h0)] reg617 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg616 = (1'h0);
  reg [(5'h12):(1'h0)] reg613 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg610 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg607 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg606 = (1'h0);
  reg [(5'h13):(1'h0)] reg604 = (1'h0);
  reg [(4'hb):(1'h0)] reg602 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg600 = (1'h0);
  reg [(2'h2):(1'h0)] reg597 = (1'h0);
  reg [(5'h13):(1'h0)] reg593 = (1'h0);
  reg [(4'h8):(1'h0)] reg592 = (1'h0);
  reg [(5'h11):(1'h0)] reg591 = (1'h0);
  reg [(5'h13):(1'h0)] reg589 = (1'h0);
  reg [(5'h1b):(1'h0)] reg587 = (1'h0);
  reg [(4'h8):(1'h0)] reg515 = (1'h0);
  reg [(5'h1c):(1'h0)] reg514 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg512 = (1'h0);
  reg [(5'h17):(1'h0)] reg511 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg509 = (1'h0);
  reg [(5'h1a):(1'h0)] reg507 = (1'h0);
  reg [(3'h5):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg503 = (1'h0);
  reg [(5'h18):(1'h0)] reg502 = (1'h0);
  reg [(5'h18):(1'h0)] reg501 = (1'h0);
  reg [(5'h19):(1'h0)] reg496 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg494 = (1'h0);
  reg [(5'h17):(1'h0)] reg493 = (1'h0);
  reg [(2'h2):(1'h0)] reg492 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg491 = (1'h0);
  reg [(3'h4):(1'h0)] reg490 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg484 = (1'h0);
  reg [(5'h14):(1'h0)] reg483 = (1'h0);
  reg [(5'h1a):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg475 = (1'h0);
  reg [(5'h1b):(1'h0)] reg474 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg472 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg471 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg470 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg468 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg462 = (1'h0);
  reg [(4'hd):(1'h0)] reg460 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg453 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg447 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg446 = (1'h0);
  reg [(5'h11):(1'h0)] reg445 = (1'h0);
  reg [(5'h1f):(1'h0)] reg444 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg440 = (1'h0);
  reg [(5'h16):(1'h0)] reg438 = (1'h0);
  reg signed [(4'he):(1'h0)] reg436 = (1'h0);
  reg [(3'h7):(1'h0)] reg435 = (1'h0);
  reg [(5'h1a):(1'h0)] reg434 = (1'h0);
  reg [(5'h19):(1'h0)] reg430 = (1'h0);
  reg [(3'h6):(1'h0)] reg429 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg424 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg421 = (1'h0);
  reg [(5'h10):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg415 = (1'h0);
  reg [(2'h2):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg402 = (1'h0);
  reg [(5'h17):(1'h0)] reg399 = (1'h0);
  reg [(4'h9):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg396 = (1'h0);
  reg [(5'h14):(1'h0)] reg393 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg389 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg386 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg383 = (1'h0);
  reg [(4'hc):(1'h0)] reg376 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg373 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg370 = (1'h0);
  reg [(5'h1a):(1'h0)] reg366 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg365 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg364 = (1'h0);
  reg [(5'h16):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg360 = (1'h0);
  reg [(3'h4):(1'h0)] reg359 = (1'h0);
  reg [(3'h4):(1'h0)] reg346 = (1'h0);
  reg [(5'h10):(1'h0)] reg345 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg343 = (1'h0);
  reg [(4'ha):(1'h0)] reg341 = (1'h0);
  reg [(5'h10):(1'h0)] reg339 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg338 = (1'h0);
  reg [(2'h2):(1'h0)] reg335 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg331 = (1'h0);
  reg [(5'h11):(1'h0)] reg330 = (1'h0);
  reg [(3'h6):(1'h0)] reg327 = (1'h0);
  reg [(3'h7):(1'h0)] reg316 = (1'h0);
  reg [(5'h14):(1'h0)] reg324 = (1'h0);
  reg [(5'h11):(1'h0)] reg321 = (1'h0);
  reg [(5'h1f):(1'h0)] reg320 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg319 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg318 = (1'h0);
  reg [(2'h2):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg313 = (1'h0);
  reg [(3'h7):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg307 = (1'h0);
  reg [(4'hb):(1'h0)] reg302 = (1'h0);
  reg [(2'h3):(1'h0)] reg300 = (1'h0);
  reg [(5'h11):(1'h0)] reg299 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg293 = (1'h0);
  reg [(5'h1c):(1'h0)] reg287 = (1'h0);
  reg [(3'h4):(1'h0)] reg284 = (1'h0);
  reg [(5'h17):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg280 = (1'h0);
  reg [(5'h1f):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg269 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg268 = (1'h0);
  reg [(5'h15):(1'h0)] reg265 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg263 = (1'h0);
  reg [(5'h1b):(1'h0)] reg259 = (1'h0);
  reg [(2'h2):(1'h0)] reg258 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg256 = (1'h0);
  reg [(3'h7):(1'h0)] reg255 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg252 = (1'h0);
  reg [(5'h1a):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg248 = (1'h0);
  reg [(5'h18):(1'h0)] reg245 = (1'h0);
  reg [(5'h1f):(1'h0)] reg244 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg243 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg238 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg237 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg236 = (1'h0);
  reg [(3'h6):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg231 = (1'h0);
  reg [(5'h1d):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg227 = (1'h0);
  reg [(5'h1f):(1'h0)] reg225 = (1'h0);
  reg [(5'h14):(1'h0)] reg218 = (1'h0);
  reg [(5'h16):(1'h0)] reg216 = (1'h0);
  reg [(3'h6):(1'h0)] reg215 = (1'h0);
  reg [(4'h9):(1'h0)] reg210 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg208 = (1'h0);
  reg [(5'h1f):(1'h0)] reg206 = (1'h0);
  reg [(5'h13):(1'h0)] reg205 = (1'h0);
  reg [(5'h14):(1'h0)] reg203 = (1'h0);
  reg [(4'hf):(1'h0)] reg201 = (1'h0);
  reg [(5'h1b):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1771 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1769 = (1'h0);
  reg [(2'h3):(1'h0)] reg1768 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar1767 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1766 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1765 = (1'h0);
  reg [(4'hf):(1'h0)] reg1764 = (1'h0);
  reg [(5'h12):(1'h0)] reg1763 = (1'h0);
  reg [(3'h7):(1'h0)] reg1760 = (1'h0);
  reg [(4'ha):(1'h0)] reg1759 = (1'h0);
  reg [(4'hb):(1'h0)] reg1758 = (1'h0);
  reg [(5'h18):(1'h0)] reg1756 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1754 = (1'h0);
  reg [(4'hf):(1'h0)] reg1751 = (1'h0);
  reg [(5'h15):(1'h0)] reg1750 = (1'h0);
  reg [(5'h16):(1'h0)] reg1749 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1740 = (1'h0);
  reg [(5'h19):(1'h0)] reg1748 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1747 = (1'h0);
  reg [(3'h7):(1'h0)] reg1746 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1745 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1743 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1737 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1736 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1735 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1719 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1730 = (1'h0);
  reg [(2'h3):(1'h0)] reg1729 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1728 = (1'h0);
  reg [(4'h9):(1'h0)] reg1727 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1723 = (1'h0);
  reg [(4'hc):(1'h0)] reg1720 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1718 = (1'h0);
  reg [(5'h12):(1'h0)] reg1716 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1715 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1713 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1711 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1710 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1709 = (1'h0);
  reg [(4'hb):(1'h0)] reg1707 = (1'h0);
  reg [(3'h7):(1'h0)] reg1706 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1704 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1703 = (1'h0);
  reg [(2'h3):(1'h0)] reg1702 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1701 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1699 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar1698 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1693 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1692 = (1'h0);
  reg [(4'ha):(1'h0)] reg1691 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1689 = (1'h0);
  reg [(5'h14):(1'h0)] reg1687 = (1'h0);
  reg [(2'h3):(1'h0)] reg1685 = (1'h0);
  reg [(2'h3):(1'h0)] reg1684 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar1682 = (1'h0);
  reg [(5'h16):(1'h0)] reg1681 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1676 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1674 = (1'h0);
  reg [(5'h18):(1'h0)] reg1678 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1676 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1674 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1672 = (1'h0);
  reg [(5'h17):(1'h0)] reg1669 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1667 = (1'h0);
  reg [(4'he):(1'h0)] reg1666 = (1'h0);
  reg [(4'he):(1'h0)] reg1663 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1662 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1661 = (1'h0);
  reg [(5'h10):(1'h0)] reg1660 = (1'h0);
  reg [(5'h15):(1'h0)] reg1659 = (1'h0);
  reg [(4'hd):(1'h0)] reg1656 = (1'h0);
  reg [(2'h2):(1'h0)] reg1653 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1652 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1650 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1614 = (1'h0);
  reg [(2'h2):(1'h0)] reg1648 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1645 = (1'h0);
  reg [(5'h18):(1'h0)] reg1642 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1641 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1640 = (1'h0);
  reg [(5'h17):(1'h0)] reg1639 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1638 = (1'h0);
  reg [(5'h11):(1'h0)] reg1635 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1634 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1633 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1631 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1630 = (1'h0);
  reg [(3'h6):(1'h0)] reg1629 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1628 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1626 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1625 = (1'h0);
  reg [(5'h19):(1'h0)] reg1624 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1623 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1622 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1619 = (1'h0);
  reg [(5'h16):(1'h0)] reg1616 = (1'h0);
  reg [(5'h14):(1'h0)] reg1611 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1608 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1602 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1601 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1597 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1595 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1593 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1592 = (1'h0);
  reg [(4'hf):(1'h0)] reg1590 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1588 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1585 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1582 = (1'h0);
  reg [(5'h16):(1'h0)] reg1581 = (1'h0);
  reg [(4'ha):(1'h0)] reg1579 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1574 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1573 = (1'h0);
  reg [(5'h18):(1'h0)] reg1570 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1569 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1568 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1567 = (1'h0);
  reg [(4'ha):(1'h0)] reg1565 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1564 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1561 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1557 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1556 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1553 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1547 = (1'h0);
  reg [(5'h18):(1'h0)] reg1546 = (1'h0);
  reg [(5'h19):(1'h0)] reg1545 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1543 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1542 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1541 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1540 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1538 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1536 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1535 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1531 = (1'h0);
  reg [(5'h19):(1'h0)] reg1530 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1526 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1522 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1521 = (1'h0);
  reg [(4'h9):(1'h0)] reg1520 = (1'h0);
  reg [(2'h3):(1'h0)] reg1519 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1518 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1515 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1514 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1513 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1512 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1511 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1510 = (1'h0);
  reg [(3'h5):(1'h0)] reg1509 = (1'h0);
  reg [(5'h14):(1'h0)] reg1506 = (1'h0);
  reg [(2'h2):(1'h0)] reg1505 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar1504 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1503 = (1'h0);
  reg [(5'h16):(1'h0)] reg1502 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1499 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1498 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1496 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg894 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg893 = (1'h0);
  reg [(4'hb):(1'h0)] reg890 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar888 = (1'h0);
  reg [(3'h6):(1'h0)] forvar887 = (1'h0);
  reg [(4'ha):(1'h0)] reg886 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg885 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg883 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg882 = (1'h0);
  reg [(5'h12):(1'h0)] reg877 = (1'h0);
  reg [(3'h5):(1'h0)] forvar876 = (1'h0);
  reg [(4'h8):(1'h0)] reg875 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg873 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar869 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg867 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg865 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg862 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg861 = (1'h0);
  reg [(5'h10):(1'h0)] reg860 = (1'h0);
  reg [(5'h1e):(1'h0)] reg857 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar855 = (1'h0);
  reg [(5'h10):(1'h0)] reg854 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar842 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg852 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg848 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar847 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg845 = (1'h0);
  reg [(5'h13):(1'h0)] reg843 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg838 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg836 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg835 = (1'h0);
  reg [(2'h2):(1'h0)] forvar829 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg814 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar811 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg831 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg830 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg829 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg826 = (1'h0);
  reg [(3'h6):(1'h0)] reg825 = (1'h0);
  reg [(5'h1b):(1'h0)] reg824 = (1'h0);
  reg [(5'h17):(1'h0)] reg823 = (1'h0);
  reg [(5'h17):(1'h0)] reg822 = (1'h0);
  reg [(5'h19):(1'h0)] reg821 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg820 = (1'h0);
  reg [(2'h3):(1'h0)] reg819 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar818 = (1'h0);
  reg [(5'h1c):(1'h0)] reg817 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg816 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar814 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg812 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg807 = (1'h0);
  reg [(5'h1a):(1'h0)] reg806 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg804 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg802 = (1'h0);
  reg [(3'h4):(1'h0)] forvar778 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar772 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg800 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg799 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg797 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg794 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg792 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg791 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg788 = (1'h0);
  reg [(4'h8):(1'h0)] reg786 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg784 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg780 = (1'h0);
  reg [(5'h19):(1'h0)] reg777 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg772 = (1'h0);
  reg [(5'h1f):(1'h0)] reg771 = (1'h0);
  reg [(3'h5):(1'h0)] reg770 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar768 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar766 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg765 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar764 = (1'h0);
  reg [(3'h7):(1'h0)] forvar761 = (1'h0);
  reg [(3'h5):(1'h0)] forvar759 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg758 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar756 = (1'h0);
  reg [(5'h14):(1'h0)] reg755 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg753 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg752 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg751 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg749 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg748 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar746 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar743 = (1'h0);
  reg [(4'he):(1'h0)] forvar740 = (1'h0);
  reg [(2'h2):(1'h0)] reg739 = (1'h0);
  reg [(5'h14):(1'h0)] reg738 = (1'h0);
  reg [(5'h1e):(1'h0)] reg737 = (1'h0);
  reg [(2'h2):(1'h0)] reg735 = (1'h0);
  reg [(3'h7):(1'h0)] reg733 = (1'h0);
  reg [(4'he):(1'h0)] forvar732 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg729 = (1'h0);
  reg [(2'h3):(1'h0)] reg725 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg723 = (1'h0);
  reg [(4'hc):(1'h0)] forvar722 = (1'h0);
  reg [(5'h1d):(1'h0)] reg721 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg720 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg719 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg715 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg714 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg712 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg711 = (1'h0);
  reg [(5'h1d):(1'h0)] reg710 = (1'h0);
  reg [(5'h15):(1'h0)] reg706 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg701 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg697 = (1'h0);
  reg signed [(4'he):(1'h0)] reg695 = (1'h0);
  reg [(4'ha):(1'h0)] reg694 = (1'h0);
  reg [(4'he):(1'h0)] reg692 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg691 = (1'h0);
  reg [(5'h1e):(1'h0)] reg690 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg687 = (1'h0);
  reg [(4'ha):(1'h0)] reg686 = (1'h0);
  reg [(5'h1f):(1'h0)] reg685 = (1'h0);
  reg [(4'hb):(1'h0)] reg684 = (1'h0);
  reg [(5'h1b):(1'h0)] reg682 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg681 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg680 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar679 = (1'h0);
  reg [(5'h15):(1'h0)] reg677 = (1'h0);
  reg signed [(4'he):(1'h0)] reg676 = (1'h0);
  reg [(4'hb):(1'h0)] forvar670 = (1'h0);
  reg [(5'h19):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg666 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg665 = (1'h0);
  reg [(4'hd):(1'h0)] reg662 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar661 = (1'h0);
  reg [(4'he):(1'h0)] forvar660 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg658 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg656 = (1'h0);
  reg [(4'hd):(1'h0)] forvar650 = (1'h0);
  reg [(4'hd):(1'h0)] reg622 = (1'h0);
  reg [(5'h1f):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg647 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg644 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg640 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg637 = (1'h0);
  reg [(4'hf):(1'h0)] reg633 = (1'h0);
  reg [(5'h1d):(1'h0)] reg632 = (1'h0);
  reg [(5'h1e):(1'h0)] reg631 = (1'h0);
  reg [(3'h7):(1'h0)] reg630 = (1'h0);
  reg [(5'h1b):(1'h0)] reg629 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg628 = (1'h0);
  reg [(5'h1d):(1'h0)] reg626 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg625 = (1'h0);
  reg [(3'h6):(1'h0)] reg623 = (1'h0);
  reg [(4'hc):(1'h0)] forvar622 = (1'h0);
  reg [(5'h15):(1'h0)] reg621 = (1'h0);
  reg [(5'h19):(1'h0)] reg615 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg614 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg611 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg609 = (1'h0);
  reg [(4'ha):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg605 = (1'h0);
  reg [(5'h13):(1'h0)] forvar603 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg601 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg599 = (1'h0);
  reg [(5'h15):(1'h0)] forvar598 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg595 = (1'h0);
  reg [(5'h15):(1'h0)] reg594 = (1'h0);
  reg [(5'h17):(1'h0)] reg590 = (1'h0);
  reg [(3'h6):(1'h0)] reg588 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg508 = (1'h0);
  reg [(4'hf):(1'h0)] forvar506 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar504 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg500 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg498 = (1'h0);
  reg [(5'h15):(1'h0)] reg497 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg495 = (1'h0);
  reg [(4'hf):(1'h0)] reg489 = (1'h0);
  reg [(5'h1a):(1'h0)] reg488 = (1'h0);
  reg [(5'h18):(1'h0)] reg487 = (1'h0);
  reg [(4'hc):(1'h0)] reg486 = (1'h0);
  reg signed [(4'he):(1'h0)] reg485 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg481 = (1'h0);
  reg [(5'h1e):(1'h0)] reg479 = (1'h0);
  reg [(5'h15):(1'h0)] reg478 = (1'h0);
  reg [(4'hd):(1'h0)] reg477 = (1'h0);
  reg [(2'h2):(1'h0)] reg476 = (1'h0);
  reg [(5'h15):(1'h0)] forvar473 = (1'h0);
  reg [(5'h11):(1'h0)] reg469 = (1'h0);
  reg [(3'h5):(1'h0)] reg467 = (1'h0);
  reg [(4'h9):(1'h0)] reg466 = (1'h0);
  reg [(5'h16):(1'h0)] reg465 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar464 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg463 = (1'h0);
  reg [(5'h12):(1'h0)] forvar461 = (1'h0);
  reg [(5'h18):(1'h0)] forvar449 = (1'h0);
  reg [(2'h2):(1'h0)] reg459 = (1'h0);
  reg [(3'h7):(1'h0)] reg458 = (1'h0);
  reg [(5'h1d):(1'h0)] reg457 = (1'h0);
  reg [(5'h15):(1'h0)] reg455 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg454 = (1'h0);
  reg [(5'h11):(1'h0)] reg452 = (1'h0);
  reg [(5'h16):(1'h0)] reg451 = (1'h0);
  reg [(5'h12):(1'h0)] reg450 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg449 = (1'h0);
  reg [(5'h19):(1'h0)] reg448 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg443 = (1'h0);
  reg [(4'hc):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg439 = (1'h0);
  reg signed [(4'he):(1'h0)] reg437 = (1'h0);
  reg [(5'h14):(1'h0)] reg433 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg432 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg431 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg428 = (1'h0);
  reg [(5'h14):(1'h0)] forvar427 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg426 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg425 = (1'h0);
  reg [(5'h1a):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg422 = (1'h0);
  reg [(5'h11):(1'h0)] reg420 = (1'h0);
  reg [(5'h15):(1'h0)] forvar419 = (1'h0);
  reg [(4'hb):(1'h0)] forvar418 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg417 = (1'h0);
  reg [(5'h1d):(1'h0)] reg413 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg412 = (1'h0);
  reg [(5'h1b):(1'h0)] reg411 = (1'h0);
  reg [(4'he):(1'h0)] reg410 = (1'h0);
  reg [(2'h2):(1'h0)] reg409 = (1'h0);
  reg [(3'h7):(1'h0)] reg408 = (1'h0);
  reg [(4'hd):(1'h0)] reg407 = (1'h0);
  reg [(4'ha):(1'h0)] forvar406 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg400 = (1'h0);
  reg [(4'hf):(1'h0)] reg397 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg395 = (1'h0);
  reg [(4'hd):(1'h0)] reg394 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg392 = (1'h0);
  reg [(5'h14):(1'h0)] forvar391 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar390 = (1'h0);
  reg [(4'he):(1'h0)] reg387 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg385 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg384 = (1'h0);
  reg signed [(4'he):(1'h0)] reg382 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg381 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg380 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg379 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg378 = (1'h0);
  reg [(4'h8):(1'h0)] reg377 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg375 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg374 = (1'h0);
  reg signed [(4'he):(1'h0)] reg372 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar369 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar367 = (1'h0);
  reg [(5'h12):(1'h0)] forvar363 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg361 = (1'h0);
  reg [(5'h1a):(1'h0)] reg358 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg357 = (1'h0);
  reg [(5'h1b):(1'h0)] reg356 = (1'h0);
  reg [(5'h1f):(1'h0)] reg355 = (1'h0);
  reg [(4'hf):(1'h0)] reg354 = (1'h0);
  reg [(5'h17):(1'h0)] forvar353 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg352 = (1'h0);
  reg [(3'h4):(1'h0)] reg349 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg348 = (1'h0);
  reg [(4'h9):(1'h0)] reg347 = (1'h0);
  reg [(4'hf):(1'h0)] reg344 = (1'h0);
  reg [(3'h6):(1'h0)] reg342 = (1'h0);
  reg [(4'h8):(1'h0)] reg340 = (1'h0);
  reg [(3'h6):(1'h0)] reg337 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg336 = (1'h0);
  reg [(3'h4):(1'h0)] reg334 = (1'h0);
  reg [(4'hf):(1'h0)] reg333 = (1'h0);
  reg [(5'h18):(1'h0)] reg332 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg329 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar328 = (1'h0);
  reg [(4'hc):(1'h0)] reg326 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg325 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg323 = (1'h0);
  reg [(2'h3):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar316 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg308 = (1'h0);
  reg [(4'h9):(1'h0)] reg306 = (1'h0);
  reg [(5'h10):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg304 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg303 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg301 = (1'h0);
  reg [(5'h10):(1'h0)] reg298 = (1'h0);
  reg [(5'h10):(1'h0)] reg297 = (1'h0);
  reg [(5'h1a):(1'h0)] reg296 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg295 = (1'h0);
  reg [(5'h1c):(1'h0)] reg294 = (1'h0);
  reg [(5'h12):(1'h0)] forvar292 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg291 = (1'h0);
  reg signed [(4'he):(1'h0)] reg290 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar289 = (1'h0);
  reg [(3'h4):(1'h0)] reg288 = (1'h0);
  reg [(5'h10):(1'h0)] reg286 = (1'h0);
  reg [(3'h4):(1'h0)] reg285 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar282 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg281 = (1'h0);
  reg [(4'hb):(1'h0)] reg279 = (1'h0);
  reg [(4'h8):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg275 = (1'h0);
  reg [(4'hc):(1'h0)] reg274 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar272 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg271 = (1'h0);
  reg [(3'h7):(1'h0)] reg267 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg266 = (1'h0);
  reg [(5'h1a):(1'h0)] reg264 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg262 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg261 = (1'h0);
  reg signed [(4'he):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg257 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg254 = (1'h0);
  reg [(5'h14):(1'h0)] reg253 = (1'h0);
  reg [(5'h18):(1'h0)] reg251 = (1'h0);
  reg [(5'h11):(1'h0)] reg250 = (1'h0);
  reg [(5'h17):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg246 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg242 = (1'h0);
  reg [(5'h12):(1'h0)] forvar241 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg240 = (1'h0);
  reg [(5'h11):(1'h0)] reg239 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg235 = (1'h0);
  reg [(4'hb):(1'h0)] forvar234 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar233 = (1'h0);
  reg [(5'h10):(1'h0)] reg229 = (1'h0);
  reg [(4'h9):(1'h0)] reg226 = (1'h0);
  reg [(4'h9):(1'h0)] reg224 = (1'h0);
  reg [(5'h1b):(1'h0)] reg223 = (1'h0);
  reg signed [(4'he):(1'h0)] reg222 = (1'h0);
  reg [(5'h14):(1'h0)] reg221 = (1'h0);
  reg [(5'h18):(1'h0)] reg220 = (1'h0);
  reg [(3'h5):(1'h0)] forvar219 = (1'h0);
  reg signed [(4'he):(1'h0)] reg217 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar214 = (1'h0);
  reg [(3'h7):(1'h0)] reg213 = (1'h0);
  reg [(5'h14):(1'h0)] forvar212 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg211 = (1'h0);
  reg [(5'h1b):(1'h0)] reg209 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg207 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg204 = (1'h0);
  reg [(5'h14):(1'h0)] reg202 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar200 = (1'h0);
  reg [(3'h5):(1'h0)] reg198 = (1'h0);
  reg [(5'h14):(1'h0)] reg197 = (1'h0);
  reg [(2'h3):(1'h0)] forvar196 = (1'h0);
  assign y = {wire1772,
                 wire1739,
                 wire1697,
                 wire1613,
                 wire1494,
                 wire754,
                 wire718,
                 wire717,
                 wire584,
                 wire516,
                 wire351,
                 wire350,
                 reg1770,
                 reg1762,
                 reg1761,
                 reg1757,
                 reg1755,
                 reg1753,
                 reg1752,
                 reg1747,
                 reg1744,
                 reg1742,
                 reg1741,
                 reg1740,
                 reg1738,
                 reg1728,
                 reg1734,
                 reg1733,
                 reg1732,
                 reg1731,
                 reg1726,
                 reg1725,
                 reg1724,
                 reg1722,
                 reg1721,
                 reg1719,
                 reg1717,
                 reg1714,
                 reg1712,
                 reg1708,
                 reg1705,
                 reg1700,
                 reg1696,
                 reg1695,
                 reg1694,
                 reg1690,
                 reg1688,
                 reg1686,
                 reg1683,
                 reg1680,
                 reg1679,
                 reg1677,
                 reg1675,
                 reg1673,
                 reg1671,
                 reg1670,
                 reg1668,
                 reg1665,
                 reg1664,
                 reg1658,
                 reg1657,
                 reg1655,
                 reg1654,
                 reg1651,
                 reg1649,
                 reg1647,
                 reg1646,
                 reg1644,
                 reg1643,
                 reg1637,
                 reg1636,
                 reg1632,
                 reg1627,
                 reg1621,
                 reg1620,
                 reg1618,
                 reg1617,
                 reg1615,
                 reg1614,
                 reg1612,
                 reg1610,
                 reg1609,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 reg1603,
                 reg1600,
                 reg1599,
                 reg1598,
                 reg1596,
                 reg1594,
                 reg1591,
                 reg1589,
                 reg1587,
                 reg1586,
                 reg1584,
                 reg1583,
                 reg1580,
                 reg1578,
                 reg1577,
                 reg1576,
                 reg1575,
                 reg1572,
                 reg1571,
                 reg1566,
                 reg1563,
                 reg1562,
                 reg1560,
                 reg1559,
                 reg1558,
                 reg1555,
                 reg1554,
                 reg1552,
                 reg1551,
                 reg1550,
                 reg1549,
                 reg1548,
                 reg1544,
                 reg1539,
                 reg1537,
                 reg1534,
                 reg1533,
                 reg1532,
                 reg1529,
                 reg1528,
                 reg1527,
                 reg1525,
                 reg1524,
                 reg1523,
                 reg1514,
                 reg1517,
                 reg1516,
                 reg1508,
                 reg1507,
                 reg1501,
                 reg1500,
                 reg1497,
                 reg895,
                 reg892,
                 reg891,
                 reg889,
                 reg884,
                 reg881,
                 reg880,
                 reg879,
                 reg878,
                 reg874,
                 reg872,
                 reg871,
                 reg870,
                 reg866,
                 reg864,
                 reg863,
                 reg859,
                 reg858,
                 reg856,
                 reg847,
                 reg853,
                 reg850,
                 reg849,
                 reg846,
                 reg844,
                 reg842,
                 reg841,
                 reg839,
                 reg837,
                 reg818,
                 reg834,
                 reg833,
                 reg832,
                 reg828,
                 reg827,
                 reg815,
                 reg813,
                 reg811,
                 reg810,
                 reg809,
                 reg808,
                 reg805,
                 reg803,
                 reg801,
                 reg798,
                 reg796,
                 reg795,
                 reg793,
                 reg790,
                 reg789,
                 reg787,
                 reg785,
                 reg783,
                 reg782,
                 reg781,
                 reg779,
                 reg778,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 reg769,
                 reg767,
                 reg763,
                 reg762,
                 reg760,
                 reg757,
                 reg750,
                 reg747,
                 reg745,
                 reg744,
                 reg742,
                 reg741,
                 reg736,
                 reg734,
                 reg731,
                 reg730,
                 reg728,
                 reg727,
                 reg726,
                 reg724,
                 reg713,
                 reg709,
                 reg708,
                 reg707,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 reg700,
                 reg699,
                 reg698,
                 reg696,
                 reg693,
                 reg689,
                 reg688,
                 reg683,
                 reg678,
                 reg675,
                 reg674,
                 reg673,
                 reg672,
                 reg671,
                 reg669,
                 reg667,
                 reg664,
                 reg663,
                 reg659,
                 reg657,
                 reg655,
                 reg654,
                 reg653,
                 reg652,
                 reg650,
                 reg649,
                 reg648,
                 reg646,
                 reg645,
                 reg643,
                 reg641,
                 reg639,
                 reg638,
                 reg636,
                 reg635,
                 reg634,
                 reg627,
                 reg624,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg613,
                 reg612,
                 reg610,
                 reg607,
                 reg606,
                 reg604,
                 reg602,
                 reg600,
                 reg597,
                 reg593,
                 reg592,
                 reg591,
                 reg589,
                 reg587,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 reg509,
                 reg507,
                 reg505,
                 reg503,
                 reg502,
                 reg501,
                 reg496,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 reg484,
                 reg483,
                 reg480,
                 reg475,
                 reg474,
                 reg472,
                 reg471,
                 reg470,
                 reg468,
                 reg462,
                 reg460,
                 reg456,
                 reg453,
                 reg447,
                 reg446,
                 reg445,
                 reg444,
                 reg440,
                 reg438,
                 reg436,
                 reg435,
                 reg434,
                 reg430,
                 reg429,
                 reg424,
                 reg421,
                 reg416,
                 reg415,
                 reg414,
                 reg403,
                 reg402,
                 reg399,
                 reg398,
                 reg396,
                 reg393,
                 reg389,
                 reg388,
                 reg386,
                 reg383,
                 reg376,
                 reg373,
                 reg371,
                 reg370,
                 reg366,
                 reg365,
                 reg364,
                 reg362,
                 reg360,
                 reg359,
                 reg346,
                 reg345,
                 reg343,
                 reg341,
                 reg339,
                 reg338,
                 reg335,
                 reg331,
                 reg330,
                 reg327,
                 reg316,
                 reg324,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg313,
                 reg312,
                 reg311,
                 reg307,
                 reg302,
                 reg300,
                 reg299,
                 reg293,
                 reg287,
                 reg284,
                 reg283,
                 reg280,
                 reg278,
                 reg276,
                 reg273,
                 reg270,
                 reg269,
                 reg268,
                 reg265,
                 reg263,
                 reg259,
                 reg258,
                 reg256,
                 reg255,
                 reg252,
                 reg249,
                 reg248,
                 reg245,
                 reg244,
                 reg243,
                 reg238,
                 reg237,
                 reg236,
                 reg232,
                 reg231,
                 reg230,
                 reg228,
                 reg227,
                 reg225,
                 reg218,
                 reg216,
                 reg215,
                 reg210,
                 reg208,
                 reg206,
                 reg205,
                 reg203,
                 reg201,
                 reg199,
                 reg1771,
                 reg1769,
                 reg1768,
                 forvar1767,
                 forvar1766,
                 reg1765,
                 reg1764,
                 reg1763,
                 reg1760,
                 reg1759,
                 reg1758,
                 reg1756,
                 reg1754,
                 reg1751,
                 reg1750,
                 reg1749,
                 forvar1740,
                 reg1748,
                 forvar1747,
                 reg1746,
                 reg1745,
                 reg1743,
                 reg1737,
                 reg1736,
                 forvar1735,
                 forvar1719,
                 reg1730,
                 reg1729,
                 forvar1728,
                 reg1727,
                 reg1723,
                 reg1720,
                 reg1718,
                 reg1716,
                 reg1715,
                 reg1713,
                 forvar1711,
                 reg1710,
                 forvar1709,
                 reg1707,
                 reg1706,
                 reg1704,
                 forvar1703,
                 reg1702,
                 reg1701,
                 reg1699,
                 forvar1698,
                 forvar1693,
                 reg1692,
                 reg1691,
                 reg1689,
                 reg1687,
                 reg1685,
                 reg1684,
                 forvar1682,
                 reg1681,
                 reg1676,
                 forvar1674,
                 reg1678,
                 forvar1676,
                 reg1674,
                 reg1672,
                 reg1669,
                 reg1667,
                 reg1666,
                 reg1663,
                 reg1662,
                 forvar1661,
                 reg1660,
                 reg1659,
                 reg1656,
                 reg1653,
                 reg1652,
                 forvar1650,
                 forvar1614,
                 reg1648,
                 reg1645,
                 reg1642,
                 forvar1641,
                 reg1640,
                 reg1639,
                 reg1638,
                 reg1635,
                 forvar1634,
                 reg1633,
                 forvar1631,
                 reg1630,
                 reg1629,
                 reg1628,
                 reg1626,
                 reg1625,
                 reg1624,
                 forvar1623,
                 reg1622,
                 reg1619,
                 reg1616,
                 reg1611,
                 reg1608,
                 forvar1602,
                 reg1601,
                 reg1597,
                 forvar1595,
                 reg1593,
                 reg1592,
                 reg1590,
                 reg1588,
                 forvar1585,
                 reg1582,
                 reg1581,
                 reg1579,
                 reg1574,
                 reg1573,
                 reg1570,
                 forvar1569,
                 reg1568,
                 reg1567,
                 reg1565,
                 forvar1564,
                 reg1561,
                 reg1557,
                 reg1556,
                 reg1553,
                 reg1547,
                 reg1546,
                 reg1545,
                 reg1543,
                 forvar1542,
                 reg1541,
                 reg1540,
                 reg1538,
                 forvar1536,
                 reg1535,
                 reg1531,
                 reg1530,
                 forvar1526,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1519,
                 reg1518,
                 reg1515,
                 forvar1514,
                 reg1513,
                 reg1512,
                 reg1511,
                 reg1510,
                 reg1509,
                 reg1506,
                 reg1505,
                 forvar1504,
                 reg1503,
                 reg1502,
                 reg1499,
                 forvar1498,
                 forvar1496,
                 reg894,
                 reg893,
                 reg890,
                 forvar888,
                 forvar887,
                 reg886,
                 reg885,
                 reg883,
                 reg882,
                 reg877,
                 forvar876,
                 reg875,
                 reg873,
                 forvar869,
                 reg868,
                 reg867,
                 reg865,
                 reg862,
                 reg861,
                 reg860,
                 reg857,
                 forvar855,
                 reg854,
                 forvar842,
                 reg852,
                 reg851,
                 reg848,
                 forvar847,
                 reg845,
                 reg843,
                 reg840,
                 reg838,
                 reg836,
                 reg835,
                 forvar829,
                 reg814,
                 forvar811,
                 reg831,
                 reg830,
                 reg829,
                 reg826,
                 reg825,
                 reg824,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 forvar818,
                 reg817,
                 reg816,
                 forvar814,
                 reg812,
                 reg807,
                 reg806,
                 reg804,
                 reg802,
                 forvar778,
                 forvar772,
                 reg800,
                 reg799,
                 reg797,
                 reg794,
                 reg792,
                 reg791,
                 reg788,
                 reg786,
                 reg784,
                 reg780,
                 reg777,
                 reg772,
                 reg771,
                 reg770,
                 forvar768,
                 forvar766,
                 reg765,
                 forvar764,
                 forvar761,
                 forvar759,
                 reg758,
                 forvar756,
                 reg755,
                 reg753,
                 reg752,
                 reg751,
                 reg749,
                 reg748,
                 forvar746,
                 forvar743,
                 forvar740,
                 reg739,
                 reg738,
                 reg737,
                 reg735,
                 reg733,
                 forvar732,
                 reg729,
                 reg725,
                 reg723,
                 forvar722,
                 reg721,
                 reg720,
                 reg719,
                 reg716,
                 reg715,
                 reg714,
                 reg712,
                 reg711,
                 reg710,
                 reg706,
                 reg701,
                 reg697,
                 reg695,
                 reg694,
                 reg692,
                 reg691,
                 reg690,
                 reg687,
                 reg686,
                 reg685,
                 reg684,
                 reg682,
                 reg681,
                 reg680,
                 forvar679,
                 reg677,
                 reg676,
                 forvar670,
                 reg668,
                 reg666,
                 reg665,
                 reg662,
                 forvar661,
                 forvar660,
                 reg658,
                 reg656,
                 forvar650,
                 reg622,
                 reg651,
                 reg647,
                 reg644,
                 reg642,
                 reg640,
                 reg637,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg626,
                 reg625,
                 reg623,
                 forvar622,
                 reg621,
                 reg615,
                 reg614,
                 reg611,
                 reg609,
                 reg608,
                 reg605,
                 forvar603,
                 reg601,
                 reg599,
                 forvar598,
                 reg596,
                 reg595,
                 reg594,
                 reg590,
                 reg588,
                 reg586,
                 reg510,
                 reg508,
                 forvar506,
                 forvar504,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg495,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg482,
                 reg481,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 forvar473,
                 reg469,
                 reg467,
                 reg466,
                 reg465,
                 forvar464,
                 reg463,
                 forvar461,
                 forvar449,
                 reg459,
                 reg458,
                 reg457,
                 reg455,
                 reg454,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg443,
                 reg442,
                 reg441,
                 reg439,
                 reg437,
                 reg433,
                 reg432,
                 reg431,
                 reg428,
                 forvar427,
                 reg426,
                 reg425,
                 reg423,
                 reg422,
                 reg420,
                 forvar419,
                 forvar418,
                 reg417,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 forvar406,
                 reg405,
                 reg404,
                 reg401,
                 reg400,
                 reg397,
                 reg395,
                 reg394,
                 reg392,
                 forvar391,
                 forvar390,
                 reg387,
                 reg385,
                 reg384,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg375,
                 reg374,
                 reg372,
                 forvar369,
                 reg368,
                 forvar367,
                 forvar363,
                 reg361,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 forvar353,
                 reg352,
                 reg349,
                 reg348,
                 reg347,
                 reg344,
                 reg342,
                 reg340,
                 reg337,
                 reg336,
                 reg334,
                 reg333,
                 reg332,
                 reg329,
                 forvar328,
                 reg326,
                 reg325,
                 reg323,
                 reg322,
                 forvar316,
                 reg315,
                 reg314,
                 reg310,
                 reg309,
                 reg308,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg301,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 forvar292,
                 reg291,
                 reg290,
                 forvar289,
                 reg288,
                 reg286,
                 reg285,
                 forvar282,
                 reg281,
                 reg279,
                 reg277,
                 reg275,
                 reg274,
                 forvar272,
                 reg271,
                 reg267,
                 reg266,
                 reg264,
                 reg262,
                 reg261,
                 reg260,
                 reg257,
                 reg254,
                 reg253,
                 reg251,
                 reg250,
                 reg241,
                 reg247,
                 reg246,
                 reg242,
                 forvar241,
                 reg240,
                 reg239,
                 reg235,
                 forvar234,
                 forvar233,
                 reg229,
                 reg226,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 reg217,
                 forvar214,
                 reg213,
                 forvar212,
                 reg211,
                 reg209,
                 reg207,
                 reg204,
                 reg202,
                 forvar200,
                 reg198,
                 reg197,
                 forvar196,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar196 = (1'h0); (forvar196 < (2'h2)); forvar196 = (forvar196 + (1'h1)))
        begin
          if ($signed((wire194[(3'h7):(3'h7)] != {((wire194 ?
                  wire194 : wire194) >> $signed(wire191)),
              (~(~|(7'h53)))})))
            begin
              reg197 = ((wire190[(1'h0):(1'h0)] ?
                      $signed((~&$unsigned(wire191))) : ((&$unsigned(forvar196)) != wire194)) ?
                  $unsigned((+$unsigned((wire195 & wire191)))) : $signed(forvar196));
            end
          else
            begin
              reg197 = $signed(wire194);
            end
          reg198 = forvar196[(2'h3):(2'h3)];
          reg199 <= (7'h4c);
        end
      for (forvar200 = (1'h0); (forvar200 < (1'h0)); forvar200 = (forvar200 + (1'h1)))
        begin
          if (($unsigned($signed(({wire190} >= reg198))) ?
              $unsigned(wire193) : (&{$signed((wire193 ? wire193 : wire195)),
                  ($unsigned(reg198) && reg197),
                  ((wire190 ^ (8'ha1)) <= $unsigned(wire194))})))
            begin
              reg201 <= (~$signed((forvar200 ?
                  forvar196[(2'h2):(2'h2)] : reg197[(4'hf):(3'h4)])));
              reg202 = $signed($signed({wire195[(5'h12):(2'h3)]}));
              reg203 <= $signed(reg198);
              reg204 = $signed(((^$signed(reg197)) ^ $signed((&(reg199 ?
                  (8'hb3) : (8'hbd))))));
              reg205 <= (!($signed(((wire194 ? wire194 : reg203) ?
                      $signed(reg203) : (wire190 >> wire190))) ?
                  $unsigned(wire194[(5'h10):(4'h9)]) : forvar200[(3'h4):(1'h1)]));
            end
          else
            begin
              reg202 = wire190;
              reg203 <= $unsigned($signed((-(^(~(7'h46))))));
              reg204 = (reg197 ?
                  ($signed((reg205[(4'hc):(1'h1)] ?
                      ((8'h9c) <<< reg204) : (+wire194))) > reg197[(4'he):(4'hb)]) : (!{(^~(wire192 ~^ (7'h4f))),
                      $unsigned(wire191),
                      (^(wire195 ? wire195 : reg205))}));
              reg205 <= {($signed(reg201) >> $unsigned($signed($signed(wire190))))};
              reg206 <= $unsigned($unsigned(((7'h46) ?
                  $unsigned(reg199) : (reg198[(2'h3):(1'h0)] >>> (wire193 ?
                      reg198 : (7'h4d))))));
              reg207 = $unsigned(reg205[(5'h10):(4'h9)]);
              reg208 <= ((~|(|wire191)) >= wire194[(1'h1):(1'h0)]);
            end
          reg209 = $unsigned($unsigned((~&(-reg203))));
          reg210 <= $signed((&wire194));
        end
      if ({reg209[(5'h1b):(4'h8)],
          (^($unsigned($signed((7'h55))) || reg199)),
          forvar196})
        begin
          reg211 = $signed(((^(~&$signed((8'ha9)))) - (|reg206)));
        end
      else
        begin
          reg211 = {wire194[(3'h7):(3'h5)]};
        end
    end
  always
    @(posedge clk) begin
      for (forvar212 = (1'h0); (forvar212 < (1'h1)); forvar212 = (forvar212 + (1'h1)))
        begin
          reg213 = $unsigned(reg208[(1'h0):(1'h0)]);
          for (forvar214 = (1'h0); (forvar214 < (3'h6)); forvar214 = (forvar214 + (1'h1)))
            begin
              reg215 <= reg210;
              reg216 <= (reg206[(5'h19):(5'h17)] ?
                  $signed((forvar214 ^~ (-(reg215 ?
                      reg203 : reg215)))) : (!(forvar212[(1'h0):(1'h0)] ?
                      (!$signed(reg206)) : {$signed((7'h4b)),
                          (reg208 ? wire190 : wire195)})));
              reg217 = (&reg215);
              reg218 <= ($signed(reg206) ?
                  $signed(((~|$unsigned((7'h43))) ?
                      (!reg208[(2'h2):(1'h0)]) : (|(reg215 ?
                          wire195 : wire192)))) : reg201);
            end
          for (forvar219 = (1'h0); (forvar219 < (2'h2)); forvar219 = (forvar219 + (1'h1)))
            begin
              reg220 = (!reg210[(3'h4):(2'h2)]);
              reg221 = reg203;
              reg222 = ((^~{($signed((8'ha8)) ?
                          wire195 : wire194[(4'hf):(4'ha)]),
                      $unsigned((reg221 ? reg215 : wire193)),
                      ((8'ha7) * forvar214)}) ?
                  (8'hb8) : wire191);
              reg223 = reg201[(1'h0):(1'h0)];
              reg224 = {$signed(reg215),
                  forvar214[(1'h0):(1'h0)],
                  reg216[(5'h13):(3'h6)]};
            end
          if (reg210[(4'h8):(3'h5)])
            begin
              reg225 <= {reg217, reg217[(3'h6):(3'h6)]};
              reg226 = reg203[(5'h14):(4'h9)];
              reg227 <= (~$signed((|forvar219[(2'h3):(2'h3)])));
              reg228 <= (!(&$signed((forvar212 << {(7'h4e), reg227}))));
              reg229 = $unsigned($signed($unsigned(($unsigned(wire193) - $unsigned(reg223)))));
              reg230 <= ($unsigned((((reg222 ? reg225 : reg206) ?
                      (wire193 ?
                          forvar212 : reg215) : $signed((8'hae))) ~^ reg224)) ?
                  wire191 : $signed((~|reg229)));
              reg231 <= reg205[(3'h7):(2'h3)];
            end
          else
            begin
              reg226 = ($unsigned($signed($signed(reg224))) >>> ($signed(reg218[(4'he):(1'h0)]) ?
                  (^~$unsigned($unsigned(reg215))) : ($unsigned(reg216) ?
                      $unsigned($unsigned(reg224)) : reg231)));
              reg227 <= (+$unsigned(reg208));
              reg228 <= reg216;
              reg230 <= $signed(wire194);
              reg231 <= wire194;
              reg232 <= ((~|$signed(reg226[(1'h0):(1'h0)])) & reg228);
            end
        end
      for (forvar233 = (1'h0); (forvar233 < (2'h2)); forvar233 = (forvar233 + (1'h1)))
        begin
          for (forvar234 = (1'h0); (forvar234 < (3'h6)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 = (((((7'h54) <= $signed(reg210)) ^ (-reg205)) || (((wire192 ?
                  reg206 : forvar214) << (reg203 == reg205)) >>> $unsigned(((7'h43) ~^ wire194)))) >= ($signed($unsigned($unsigned((7'h53)))) ?
                  $signed(reg226) : reg231));
              reg236 <= $unsigned({$signed($signed(reg206[(5'h1d):(5'h11)]))});
              reg237 <= {(~^(~|{$unsigned((8'hac))}))};
              reg238 <= (-$signed($signed(reg203[(4'he):(1'h0)])));
              reg239 = reg218[(3'h6):(1'h1)];
            end
        end
      reg240 = {$unsigned($signed(forvar212)), reg221};
      if ($signed({(+$unsigned(((8'h9d) ? wire194 : (8'hb3)))), (8'hae)}))
        begin
          for (forvar241 = (1'h0); (forvar241 < (3'h4)); forvar241 = (forvar241 + (1'h1)))
            begin
              reg242 = $signed((~|((-wire192) <= $signed($unsigned(reg235)))));
              reg243 <= reg205[(2'h3):(2'h3)];
              reg244 <= $signed((^~(8'haa)));
              reg245 <= forvar212[(4'h8):(1'h0)];
              reg246 = $signed(reg213);
            end
          reg247 = (^(~&wire194));
        end
      else
        begin
          reg241 = wire191[(3'h7):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      if ({wire190[(2'h2):(2'h2)],
          $unsigned((reg228 ?
              $unsigned({reg230}) : ({reg218} ?
                  $unsigned(wire190) : (8'hb7))))})
        begin
          reg248 <= (!reg227[(4'hd):(4'hb)]);
          reg249 <= $signed((+reg245[(2'h2):(1'h0)]));
          reg250 = reg205;
          reg251 = reg249;
        end
      else
        begin
          reg248 <= (reg206 <= wire191);
          if (wire194)
            begin
              reg249 <= reg227[(5'h15):(4'h9)];
              reg252 <= {(&reg228), (&(^reg244)), reg206[(4'hc):(3'h7)]};
              reg253 = (reg248[(3'h4):(1'h0)] ?
                  ($unsigned($signed((wire192 ?
                      reg228 : wire194))) && (|(~reg205[(4'he):(4'hb)]))) : reg206);
              reg254 = $unsigned(reg249[(5'h18):(4'hc)]);
              reg255 <= reg228[(4'hb):(4'h8)];
              reg256 <= $signed($unsigned((|reg208)));
            end
          else
            begin
              reg249 <= $unsigned((&$unsigned({reg236})));
              reg252 <= $signed(reg206);
              reg255 <= {(~|$signed(((reg253 >= reg255) ?
                      wire195 : {reg232, reg250}))),
                  $signed(reg238[(1'h1):(1'h1)])};
              reg257 = reg208[(2'h2):(2'h2)];
              reg258 <= (reg215[(1'h1):(1'h1)] && wire194[(3'h4):(1'h1)]);
              reg259 <= wire195[(2'h3):(1'h1)];
              reg260 = (($unsigned(($signed((7'h41)) ~^ (reg232 ?
                          reg250 : reg225))) ?
                      $unsigned($signed((+reg238))) : reg257[(4'hd):(4'ha)]) ?
                  ((reg231 < ($signed(reg205) >>> $unsigned(wire190))) ?
                      $signed(reg228) : (!(!(reg201 ?
                          wire194 : reg228)))) : $unsigned((~^reg208[(1'h0):(1'h0)])));
            end
        end
    end
  always
    @(posedge clk) begin
      reg261 = $unsigned((~($signed(reg255[(3'h6):(1'h0)]) ?
          $signed($unsigned(reg203)) : ((!reg245) ?
              $unsigned(reg238) : reg201[(4'hc):(4'hb)]))));
    end
  always
    @(posedge clk) begin
      if ((reg225 >> ($unsigned(((&reg228) ?
              (reg243 << reg243) : (reg244 + (7'h4f)))) ?
          $unsigned($signed($unsigned(wire195))) : (~|(~^reg206)))))
        begin
          reg262 = (reg249[(4'hb):(2'h2)] ?
              $signed((({reg255, wire195} ?
                      (reg252 ? reg244 : reg215) : reg236[(1'h1):(1'h1)]) ?
                  {(reg232 ? (8'ha8) : wire194), reg259} : ({reg255,
                      reg245,
                      reg231} <= $unsigned(reg216)))) : reg225);
        end
      else
        begin
          if (reg216)
            begin
              reg263 <= ($signed(reg262[(3'h4):(2'h3)]) + (~|((reg216[(4'h8):(2'h3)] ?
                      reg225[(4'hc):(1'h1)] : {wire192, reg215, reg248}) ?
                  $signed(reg210) : $unsigned((~&(8'ha6))))));
              reg264 = (7'h4e);
              reg265 <= (8'hae);
              reg266 = $signed($unsigned($unsigned(wire194[(4'he):(1'h0)])));
              reg267 = reg244[(2'h2):(2'h2)];
            end
          else
            begin
              reg263 <= $signed((8'ha9));
              reg265 <= ((+reg208) ? (~&(wire190 - (8'ha4))) : reg259);
              reg268 <= (|$signed(reg245));
              reg269 <= reg205[(4'hc):(4'h8)];
              reg270 <= $signed($signed(reg245));
            end
          reg271 = (-$unsigned($signed({$signed(reg210),
              reg264,
              (reg268 ? reg259 : reg244)})));
          for (forvar272 = (1'h0); (forvar272 < (2'h3)); forvar272 = (forvar272 + (1'h1)))
            begin
              reg273 <= (reg262[(3'h5):(2'h3)] == ({(|reg206[(4'h8):(3'h5)])} ?
                  (reg237 ?
                      $unsigned($signed(reg230)) : ((forvar272 ?
                          reg208 : reg231) && $unsigned(reg216))) : $signed((|reg244))));
            end
          if ((reg269[(5'h18):(3'h5)] <= (reg270[(4'hd):(1'h1)] ?
              (reg243 <<< ((reg236 > reg228) ?
                  $signed(reg205) : (reg269 ? reg236 : reg201))) : forvar272)))
            begin
              reg274 = $unsigned(($unsigned($unsigned((reg216 ?
                  reg266 : (8'ha4)))) >> $signed(($signed(reg255) != $unsigned(reg232)))));
              reg275 = reg271[(4'h9):(4'h9)];
              reg276 <= wire193[(4'hf):(4'hf)];
              reg277 = (8'hbf);
              reg278 <= ({{((!reg245) ?
                          $signed(reg244) : reg273[(4'hf):(3'h6)]),
                      $signed($unsigned(wire193)),
                      ({reg273} ? (forvar272 < (8'hb4)) : $signed(reg245))},
                  $unsigned($signed($signed(reg256)))} * reg274[(3'h4):(3'h4)]);
              reg279 = ({$signed((wire195[(1'h0):(1'h0)] | reg276[(3'h5):(3'h4)]))} ?
                  ({$signed(reg267)} ?
                      reg255[(1'h0):(1'h0)] : $signed($unsigned((reg231 + (8'hb5))))) : $unsigned({(~&reg269)}));
            end
          else
            begin
              reg274 = reg227;
              reg275 = {reg256, ($unsigned(wire191) ^~ reg215[(2'h2):(1'h1)])};
              reg276 <= $signed($unsigned((((7'h54) & reg275[(4'h9):(3'h7)]) >> reg206[(3'h5):(3'h5)])));
              reg277 = reg225;
              reg278 <= (reg274[(3'h7):(1'h0)] + (-reg279[(3'h5):(3'h5)]));
              reg280 <= reg278;
              reg281 = $unsigned((reg258 ?
                  $signed(($unsigned(wire191) * (reg269 == reg255))) : $signed(reg265[(4'ha):(3'h4)])));
            end
          for (forvar282 = (1'h0); (forvar282 < (1'h0)); forvar282 = (forvar282 + (1'h1)))
            begin
              reg283 <= (~|((reg203[(4'h8):(4'h8)] * reg270) ~^ $signed((~$signed(reg203)))));
              reg284 <= ({reg231[(4'hf):(4'h8)],
                      $signed(reg269[(2'h2):(1'h1)]),
                      (8'had)} ?
                  reg243[(3'h6):(1'h0)] : (($unsigned(((8'hb4) ?
                          reg231 : reg280)) < $signed($signed(reg283))) ?
                      {$unsigned(wire190),
                          (~$unsigned((7'h44)))} : (^~{reg199[(5'h12):(3'h7)],
                          (reg280 << (8'ha5))})));
              reg285 = ($signed(((reg264 ? (|reg243) : (reg269 >>> reg243)) ?
                      (((7'h4d) && reg236) ?
                          (reg262 ? (8'ha5) : reg203) : (reg237 ?
                              reg238 : (7'h54))) : {reg248[(1'h1):(1'h1)],
                          $unsigned(reg238),
                          (-reg265)})) ?
                  $signed(({(reg273 ? reg264 : reg231),
                      $unsigned(reg281),
                      {reg270}} > $signed($unsigned(reg259)))) : $signed($signed((reg256[(5'h11):(5'h10)] ?
                      (~^reg258) : $signed(reg236)))));
              reg286 = reg210[(4'h8):(3'h7)];
              reg287 <= ({$signed(($signed((7'h4c)) & $signed(wire191)))} ?
                  ((reg199[(5'h13):(4'hf)] ?
                      {$signed(reg227)} : ((reg218 ?
                          reg256 : reg216) ^~ reg255)) || ({(reg248 ?
                          (7'h58) : reg278)} >= $unsigned({reg208}))) : (reg237[(3'h6):(2'h2)] ^~ reg205[(3'h4):(1'h1)]));
            end
          reg288 = reg228[(5'h13):(5'h13)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar289 = (1'h0); (forvar289 < (1'h1)); forvar289 = (forvar289 + (1'h1)))
        begin
          reg290 = reg245[(2'h2):(2'h2)];
          reg291 = (reg237[(2'h2):(1'h1)] ?
              (+{$unsigned($unsigned(reg225))}) : (~&reg231));
          for (forvar292 = (1'h0); (forvar292 < (2'h2)); forvar292 = (forvar292 + (1'h1)))
            begin
              reg293 <= (reg278 ?
                  (~|(|(wire191 ~^ $signed(reg291)))) : $unsigned($signed(reg263)));
              reg294 = reg203[(4'h9):(4'h8)];
              reg295 = {reg258[(1'h1):(1'h0)],
                  reg259,
                  {(^$unsigned(reg248[(1'h1):(1'h1)])),
                      (~$signed((7'h53))),
                      (8'hbc)}};
              reg296 = reg295[(1'h0):(1'h0)];
              reg297 = (|reg230);
              reg298 = reg268;
              reg299 <= ($signed({$signed(wire190),
                      (-(~^reg227)),
                      (!(reg249 ? reg280 : reg278))}) ?
                  (|reg265) : $unsigned((~^({reg263,
                      reg210} == reg291[(2'h3):(2'h3)]))));
            end
          if ($unsigned(reg199))
            begin
              reg300 <= (-$signed((((7'h50) && (|reg210)) <<< {(^reg245)})));
              reg301 = reg270;
              reg302 <= (reg284 | $unsigned(($signed($signed(reg259)) > reg263)));
            end
          else
            begin
              reg300 <= $signed($unsigned($unsigned({((7'h4b) >> wire194)})));
              reg301 = reg218[(4'hd):(4'h8)];
              reg303 = reg269;
              reg304 = (+$signed(reg232[(1'h0):(1'h0)]));
              reg305 = reg228[(2'h2):(1'h0)];
              reg306 = reg296;
            end
          reg307 <= (reg215[(1'h1):(1'h0)] ~^ $signed(reg306[(2'h2):(1'h0)]));
          reg308 = ($unsigned((reg236 - wire195)) ?
              ((reg236[(1'h1):(1'h0)] || reg278) ~^ reg227) : {$signed(wire195[(2'h2):(2'h2)]),
                  (~(-(wire194 ? reg201 : (8'ha7)))),
                  (~|reg258)});
        end
      if ($signed(((^{$unsigned(reg230), (-reg210), reg300}) ?
          $signed($unsigned($unsigned(reg215))) : (-(&(forvar292 ?
              reg237 : reg252))))))
        begin
          if (((^($signed((reg199 ? reg255 : reg205)) ?
              (reg300 < (wire190 <<< reg299)) : reg218)) || ({$signed($signed(reg300)),
                  reg216[(5'h15):(4'hd)],
                  {(reg299 ? reg258 : (8'hb5)),
                      $signed(reg232),
                      $signed(reg295)}} ?
              {(~|(7'h54)), $unsigned(((7'h55) ^ reg256))} : (reg290 ?
                  $unsigned($signed(reg230)) : reg218[(4'he):(4'h8)]))))
            begin
              reg309 = (^~(wire190 >> $unsigned(reg249)));
              reg310 = (($signed(((~|reg208) ?
                  reg265 : (reg227 ?
                      (7'h42) : reg276))) * $signed(reg231)) * ((~|reg280[(3'h6):(3'h5)]) ?
                  $signed({(reg206 & (8'hbf))}) : (&(+((8'hb4) ~^ reg228)))));
              reg311 <= $unsigned((^~$unsigned(forvar289[(1'h1):(1'h1)])));
              reg312 <= reg205[(4'hc):(3'h4)];
            end
          else
            begin
              reg311 <= (((^~(^~$signed(wire192))) ?
                      reg296[(2'h3):(2'h3)] : (($signed(reg208) <<< reg236[(3'h5):(2'h2)]) ?
                          reg276[(2'h3):(1'h0)] : reg283)) ?
                  $signed(reg298) : (8'ha0));
              reg312 <= ($signed((+reg283[(3'h5):(2'h2)])) ?
                  $unsigned(reg269[(3'h6):(1'h0)]) : (forvar289[(3'h7):(3'h6)] >= reg215[(1'h1):(1'h0)]));
              reg313 <= $signed(((reg290 < reg228) << (~|reg216)));
              reg314 = (~^($signed({reg201[(4'hf):(4'hb)]}) & ($signed({reg258,
                  reg291,
                  reg308}) != reg206[(4'hc):(3'h7)])));
              reg315 = ($signed(($unsigned($unsigned(wire193)) ^ $signed((reg301 > reg296)))) ?
                  $signed($unsigned({reg230, (reg215 > reg269)})) : wire190);
            end
          for (forvar316 = (1'h0); (forvar316 < (2'h3)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg317 <= forvar316;
              reg318 <= ($unsigned($signed($signed($unsigned(reg298)))) ?
                  (reg205 != (reg225[(3'h6):(1'h0)] || (|$signed(reg301)))) : ($unsigned(reg268[(3'h6):(1'h0)]) >>> $unsigned(reg265[(4'hb):(3'h6)])));
              reg319 <= $signed((&$unsigned($signed(forvar292[(1'h0):(1'h0)]))));
              reg320 <= {$signed(reg248),
                  (~|$unsigned((&(~&reg294)))),
                  $unsigned($signed($signed((reg312 <<< reg301))))};
              reg321 <= reg295[(3'h6):(1'h1)];
              reg322 = reg205;
              reg323 = reg284;
            end
          reg324 <= reg323;
        end
      else
        begin
          reg309 = (^~(~^reg270));
          reg311 <= reg306[(1'h0):(1'h0)];
          if ((8'hb5))
            begin
              reg314 = (~^reg232);
              reg315 = reg199;
              reg316 <= (reg298 ?
                  $signed($unsigned(($unsigned((7'h4e)) != (reg273 ?
                      (8'hb7) : reg297)))) : reg323[(5'h1f):(5'h10)]);
              reg317 <= $unsigned((-{((reg319 <<< reg216) ?
                      $signed(reg205) : {reg317})}));
              reg318 <= reg228[(5'h18):(5'h17)];
              reg319 <= reg249;
              reg320 <= (8'hac);
            end
          else
            begin
              reg314 = reg301[(1'h1):(1'h0)];
              reg316 <= $signed($unsigned(($signed(reg263[(3'h6):(1'h0)]) ?
                  (!reg228) : (8'hb8))));
              reg322 = ((~^reg215) << {($signed(reg318[(3'h4):(1'h0)]) ?
                      (^$signed(reg228)) : reg276[(3'h6):(2'h3)]),
                  reg293});
              reg324 <= $unsigned({$unsigned({{reg307, reg230, reg228}}),
                  reg310,
                  (reg291 ? reg206 : reg230[(1'h0):(1'h0)])});
              reg325 = $signed((reg243[(3'h6):(1'h1)] ?
                  (&({reg280, (8'hb2)} ?
                      (-reg270) : (reg256 - reg300))) : $signed(reg309[(4'h9):(3'h6)])));
              reg326 = ($signed({(~|reg206[(2'h3):(2'h3)]),
                  ($signed(reg227) ?
                      (reg276 ?
                          reg244 : reg297) : (reg227 >> reg296))}) & reg228[(5'h10):(4'hd)]);
            end
        end
      reg327 <= reg215[(2'h3):(2'h2)];
      for (forvar328 = (1'h0); (forvar328 < (2'h3)); forvar328 = (forvar328 + (1'h1)))
        begin
          reg329 = forvar316[(2'h3):(1'h0)];
          reg330 <= (reg312[(1'h1):(1'h1)] ?
              (~|(($unsigned(reg273) ^ (~reg201)) < (|$unsigned((8'hb9))))) : reg252[(3'h5):(1'h0)]);
          reg331 <= (+forvar328[(5'h15):(4'hc)]);
          reg332 = {{reg210}};
        end
      reg333 = $unsigned($unsigned((~^reg327)));
    end
  always
    @(posedge clk) begin
      if (((|(({reg228} == $signed((8'ha5))) < $signed(wire190[(4'h9):(2'h3)]))) ?
          $signed((~^reg293[(3'h4):(3'h4)])) : (reg299[(4'ha):(1'h1)] ?
              {({reg258} ? (reg269 ? reg230 : (7'h49)) : (-wire194)),
                  ((reg249 ? reg225 : wire190) ?
                      reg331 : {reg327,
                          (8'h9d),
                          reg330})} : {(!$unsigned((8'hbe))),
                  {(reg284 ? reg263 : wire190), (~|reg331)}})))
        begin
          if ((8'hba))
            begin
              reg334 = (reg327 >= reg313);
              reg335 <= ($unsigned($unsigned($unsigned({reg316}))) ?
                  reg312[(2'h2):(1'h0)] : {(|$unsigned($unsigned(reg265))),
                      (~&((reg316 ^ reg280) ?
                          (~&wire192) : $unsigned(reg210)))});
              reg336 = (($unsigned($signed((^~reg284))) & reg205[(3'h4):(2'h3)]) < $signed((-((-reg259) && $signed(reg268)))));
              reg337 = reg265;
            end
          else
            begin
              reg334 = (reg293 == reg232);
              reg336 = reg316[(1'h1):(1'h0)];
              reg338 <= reg278[(3'h6):(1'h0)];
              reg339 <= reg320[(3'h7):(3'h4)];
              reg340 = $signed($unsigned(reg320[(4'h8):(3'h7)]));
              reg341 <= {reg336};
              reg342 = ((reg208[(2'h2):(1'h1)] > (~&reg218)) ?
                  ($unsigned($signed((reg206 ^~ (8'hac)))) << $unsigned(reg243)) : reg258);
            end
          if (reg245)
            begin
              reg343 <= reg225;
            end
          else
            begin
              reg343 <= $unsigned(((reg334[(1'h1):(1'h1)] ?
                  (reg319[(2'h3):(1'h1)] != (reg256 < wire192)) : reg330[(4'h8):(4'h8)]) && {(^~reg248),
                  reg206[(5'h1c):(2'h2)]}));
              reg344 = ((&reg248[(1'h0):(1'h0)]) | ((~&(~&(|reg284))) ^~ $signed({reg249[(4'hf):(1'h0)],
                  $unsigned(reg228)})));
              reg345 <= reg208[(1'h0):(1'h0)];
              reg346 <= (reg256 << reg237[(2'h2):(2'h2)]);
            end
          reg347 = $unsigned(((~|$signed((7'h4c))) ?
              $signed($signed($signed(reg311))) : reg256[(5'h16):(4'hb)]));
          reg348 = (reg199[(3'h6):(3'h4)] | $signed((reg337 ?
              ((reg205 ? (7'h49) : wire193) + $unsigned(reg265)) : reg330)));
          reg349 = {(^((^{reg206}) ? ($signed(wire192) | (~reg231)) : reg302))};
        end
      else
        begin
          reg334 = reg265[(3'h4):(1'h0)];
          if ((^~({(reg252[(3'h4):(1'h0)] ?
                  reg287[(4'hb):(2'h2)] : (reg302 >>> (8'hb9))),
              reg225[(5'h1f):(5'h10)]} >>> $unsigned(reg324))))
            begin
              reg335 <= $signed($unsigned((~^(reg269[(5'h15):(3'h6)] ?
                  (reg252 & reg346) : {reg313}))));
              reg336 = reg346[(2'h3):(2'h3)];
              reg337 = ((|$unsigned(((-reg244) ?
                  reg216[(5'h16):(5'h15)] : reg259))) * $unsigned($signed((((8'h9c) ?
                      reg348 : (8'hb7)) ?
                  $signed((7'h52)) : (7'h57)))));
              reg340 = reg225[(4'hb):(2'h3)];
              reg342 = (reg340[(3'h5):(3'h4)] ?
                  $unsigned($unsigned(reg230[(3'h7):(2'h3)])) : $unsigned($unsigned(reg201)));
              reg344 = reg249;
            end
          else
            begin
              reg336 = {reg293, wire195[(4'h9):(1'h1)], {(7'h48)}};
              reg338 <= (reg334 >>> reg206);
              reg339 <= (&($signed(reg206[(3'h6):(3'h6)]) ? reg319 : reg243));
            end
        end
    end
  assign wire350 = (8'hb9);
  assign wire351 = reg327;
  always
    @(posedge clk) begin
      reg352 = reg345;
      for (forvar353 = (1'h0); (forvar353 < (3'h4)); forvar353 = (forvar353 + (1'h1)))
        begin
          if ((-{(+$unsigned($unsigned(reg339))),
              (!(!wire350[(4'h8):(1'h0)])),
              $unsigned((reg215 <<< $unsigned(reg338)))}))
            begin
              reg354 = {reg231[(1'h0):(1'h0)], wire195};
              reg355 = ($unsigned($unsigned(($unsigned(reg341) ^~ reg354))) > reg269);
              reg356 = (wire193[(5'h12):(4'h9)] < $unsigned(($signed(reg237) > ({forvar353,
                  reg287} <<< forvar353[(5'h15):(5'h10)]))));
              reg357 = reg228[(4'hf):(4'hc)];
              reg358 = ($unsigned($signed(($unsigned(reg216) || $signed(reg338)))) >> reg263);
            end
          else
            begin
              reg359 <= (-reg203);
              reg360 <= (+(reg249[(2'h3):(2'h3)] & $signed({reg354[(4'he):(3'h5)],
                  $unsigned((8'ha7)),
                  (8'hbf)})));
              reg361 = (8'hbe);
              reg362 <= reg215[(3'h5):(2'h3)];
            end
          for (forvar363 = (1'h0); (forvar363 < (2'h3)); forvar363 = (forvar363 + (1'h1)))
            begin
              reg364 <= reg248;
              reg365 <= $unsigned({reg199[(5'h13):(4'hd)],
                  ({{wire193, reg244, reg338},
                          (reg319 ? reg249 : reg263),
                          reg280[(4'h8):(3'h7)]} ?
                      ($signed(reg331) ?
                          $unsigned(reg293) : $unsigned(reg230)) : ((reg330 ?
                          wire190 : wire194) | reg268[(4'h8):(3'h7)]))});
              reg366 <= ($unsigned(reg280[(1'h0):(1'h0)]) >>> $unsigned((^reg228)));
            end
        end
      for (forvar367 = (1'h0); (forvar367 < (3'h4)); forvar367 = (forvar367 + (1'h1)))
        begin
          reg368 = ((((~{reg269}) ?
                  (!$unsigned(reg248)) : ((&(7'h4f)) ?
                      wire195 : reg331[(3'h5):(2'h2)])) ?
              reg318[(3'h4):(3'h4)] : reg236[(1'h0):(1'h0)]) || reg228[(5'h12):(1'h0)]);
          for (forvar369 = (1'h0); (forvar369 < (2'h2)); forvar369 = (forvar369 + (1'h1)))
            begin
              reg370 <= (!((^reg236[(3'h4):(1'h0)]) ?
                  $signed($unsigned(forvar367[(5'h11):(4'hd)])) : {(~^(reg338 != reg269)),
                      $signed(reg248[(1'h0):(1'h0)])}));
              reg371 <= reg230[(4'he):(2'h3)];
              reg372 = $unsigned(reg245[(2'h3):(1'h0)]);
              reg373 <= ($unsigned({((7'h52) ?
                      (reg338 >> reg372) : (reg335 != (8'hb8))),
                  forvar369[(4'hc):(4'ha)]}) == (reg346 ?
                  $signed((~wire194)) : (|(reg216[(4'hd):(4'hc)] ?
                      reg352 : forvar367[(4'hd):(1'h1)]))));
              reg374 = ($signed((forvar367 ?
                      (reg225[(5'h1d):(5'h1c)] || {reg210}) : wire193)) ?
                  (7'h58) : (&(((reg269 ? wire191 : reg355) || {reg317,
                      reg338}) ^~ reg360[(5'h17):(4'ha)])));
              reg375 = $signed(($signed((~^(^reg284))) ?
                  reg366[(1'h0):(1'h0)] : $signed($unsigned(reg299))));
              reg376 <= reg293;
            end
          reg377 = forvar353[(4'hb):(4'h8)];
          reg378 = $signed({reg358[(4'hc):(4'hb)],
              {(reg228[(5'h1a):(2'h2)] ? $signed(reg354) : $signed(wire350)),
                  ($unsigned(reg331) ? (~^reg249) : {reg373})}});
          reg379 = $unsigned(reg273);
          if ({reg376,
              {$unsigned(reg265[(5'h10):(4'hc)]),
                  {$signed(reg321[(4'hf):(4'h9)]),
                      reg359[(1'h1):(1'h1)],
                      (~(reg227 ? reg377 : wire193))},
                  $signed({reg263[(2'h3):(1'h1)]})}})
            begin
              reg380 = ($signed({($unsigned(reg278) ?
                      (reg287 ?
                          reg365 : (8'ha5)) : (wire350 || reg320))}) > $signed($signed(reg366)));
              reg381 = $unsigned(reg358);
              reg382 = $unsigned($unsigned(reg265));
              reg383 <= {(^(reg343 + reg374))};
              reg384 = ({(((reg238 | reg320) <<< reg366[(5'h10):(4'hd)]) ~^ {$unsigned(reg248)}),
                  $unsigned((!reg299))} & reg238[(3'h4):(3'h4)]);
              reg385 = $unsigned(reg338);
              reg386 <= {(~|((reg276[(3'h6):(3'h4)] < $unsigned(reg225)) > reg361[(3'h7):(2'h2)])),
                  forvar367[(5'h16):(4'hf)]};
            end
          else
            begin
              reg380 = {reg345[(3'h7):(1'h0)]};
              reg383 <= ($signed({reg360}) ^~ $signed(reg370[(3'h5):(1'h0)]));
              reg384 = (&({reg243[(3'h7):(1'h1)],
                  {{reg365, reg380}},
                  ($unsigned(reg232) >= {(7'h47)})} < ((reg338 ?
                      $signed(reg358) : (8'ha2)) ?
                  reg227[(4'ha):(3'h5)] : reg216[(1'h0):(1'h0)])));
            end
          reg387 = {reg255[(1'h1):(1'h1)],
              $unsigned({(!(~&reg273)), (!{reg354, (7'h51)})}),
              $signed($signed(((^~reg299) ?
                  {reg379, reg243, reg384} : (&reg273))))};
        end
      reg388 <= ($signed(reg311[(3'h6):(3'h5)]) ?
          $unsigned(reg205) : (+$unsigned(forvar369)));
      reg389 <= reg358;
      for (forvar390 = (1'h0); (forvar390 < (1'h0)); forvar390 = (forvar390 + (1'h1)))
        begin
          for (forvar391 = (1'h0); (forvar391 < (3'h6)); forvar391 = (forvar391 + (1'h1)))
            begin
              reg392 = ((({(!reg299)} ?
                          ((wire194 ?
                              reg379 : reg268) ^ (8'haf)) : ($signed(reg230) ?
                              $signed(reg228) : reg278)) ?
                      $unsigned($unsigned($unsigned(wire192))) : (~^$unsigned((reg341 <= reg389)))) ?
                  ((-$signed((reg378 ?
                      (7'h45) : reg379))) >= reg354) : (|$signed(reg236)));
              reg393 <= reg352;
              reg394 = ({(reg364 <<< ($signed(reg392) ?
                          ((8'h9e) ^ wire193) : (reg346 ~^ reg360)))} ?
                  reg381 : reg387[(1'h0):(1'h0)]);
              reg395 = (&((8'hae) ?
                  ((reg319[(2'h2):(1'h1)] | (&(8'hb1))) * $signed($signed((8'had)))) : reg299));
              reg396 <= (-$signed((((reg230 * reg249) ?
                  (|reg205) : $signed(reg307)) != $signed(reg199[(4'he):(4'h9)]))));
            end
          reg397 = $signed($signed($signed($signed(reg311))));
          if (reg227)
            begin
              reg398 <= reg385;
              reg399 <= {$signed(reg379),
                  (reg376 ?
                      $unsigned((reg324 ?
                          wire193[(5'h12):(3'h5)] : (reg300 ^~ reg268))) : reg299[(4'hc):(4'hb)])};
              reg400 = (8'h9e);
              reg401 = ((8'hb5) < wire194);
              reg402 <= $unsigned($signed((reg265 || (7'h47))));
            end
          else
            begin
              reg400 = ((~&($signed((reg276 >= reg394)) ?
                      $signed($unsigned(reg238)) : {(wire190 ^ (8'h9f))})) ?
                  (reg218 ^ $unsigned($signed((7'h49)))) : $signed($unsigned({(wire351 >= reg287),
                      (wire193 ? reg287 : (8'hb0))})));
              reg401 = reg230;
              reg402 <= ((8'ha4) ^~ reg386);
              reg403 <= reg283[(2'h2):(1'h1)];
              reg404 = $unsigned(reg366);
              reg405 = $unsigned(((~|($unsigned(reg388) + (8'ha9))) < $signed((|{wire190,
                  (8'ha6)}))));
            end
          for (forvar406 = (1'h0); (forvar406 < (2'h3)); forvar406 = (forvar406 + (1'h1)))
            begin
              reg407 = {$unsigned((7'h4b)),
                  (reg320 ?
                      ((8'hb5) && ($signed((8'had)) >>> (reg379 & reg276))) : $unsigned((((8'ha7) <= reg318) ?
                          $unsigned((7'h4d)) : reg356[(4'he):(4'ha)])))};
              reg408 = reg396;
              reg409 = reg252;
              reg410 = $signed(reg377);
              reg411 = reg356[(3'h7):(3'h6)];
            end
          if (reg389[(2'h2):(2'h2)])
            begin
              reg412 = ((reg243 ?
                      ((^$signed(wire351)) ?
                          $signed($signed(reg409)) : reg380) : (7'h45)) ?
                  reg236[(3'h5):(2'h2)] : (~^$signed({$unsigned(reg302),
                      {reg411, reg402}})));
              reg413 = $unsigned((^~forvar391[(4'hd):(4'hd)]));
              reg414 <= (reg388[(4'hf):(3'h7)] ?
                  wire350[(2'h3):(1'h1)] : (($signed((-reg379)) >= $unsigned((reg355 ?
                      reg374 : reg244))) ^ $signed({$unsigned((7'h56))})));
            end
          else
            begin
              reg414 <= reg284[(1'h1):(1'h0)];
              reg415 <= (reg382[(4'hc):(4'hc)] ?
                  reg327 : ({reg372[(4'ha):(1'h0)], reg370[(3'h6):(1'h1)]} ?
                      ((((8'hae) < reg218) ?
                              (^~reg365) : reg381[(3'h4):(1'h1)]) ?
                          ((-reg377) >> $unsigned((8'ha3))) : {wire351[(2'h3):(1'h1)]}) : ((reg366[(5'h18):(4'h9)] >> $unsigned(reg381)) ?
                          reg368 : (reg380[(2'h2):(1'h1)] != {reg387,
                              (8'hbc),
                              reg225}))));
              reg416 <= reg313;
              reg417 = reg216;
            end
        end
      for (forvar418 = (1'h0); (forvar418 < (2'h2)); forvar418 = (forvar418 + (1'h1)))
        begin
          for (forvar419 = (1'h0); (forvar419 < (3'h6)); forvar419 = (forvar419 + (1'h1)))
            begin
              reg420 = wire351[(4'hf):(4'hb)];
              reg421 <= reg216;
              reg422 = forvar390;
              reg423 = (|wire350[(4'h8):(3'h4)]);
              reg424 <= ($signed(($unsigned(reg387) ?
                  {(^~forvar406),
                      (reg393 ? reg368 : reg355),
                      forvar391[(4'hf):(3'h7)]} : {reg408,
                      $signed(reg318),
                      ((8'hb7) != reg358)})) <<< reg284);
              reg425 = (&reg377[(4'h8):(3'h5)]);
            end
          reg426 = (~^(wire192 == (($signed(reg302) <<< $signed(reg364)) ?
              $unsigned(reg358) : $unsigned($unsigned(reg409)))));
          for (forvar427 = (1'h0); (forvar427 < (2'h3)); forvar427 = (forvar427 + (1'h1)))
            begin
              reg428 = {($unsigned($unsigned(reg320[(5'h1e):(4'h8)])) ?
                      (~|$signed(reg265[(4'h9):(3'h4)])) : (reg393[(4'hc):(3'h5)] > $unsigned($unsigned((7'h56))))),
                  $unsigned(reg252[(2'h2):(1'h0)]),
                  ((reg299 + reg330) ?
                      reg330[(3'h5):(2'h3)] : ((-(^~reg316)) + $signed(reg317[(2'h2):(1'h0)])))};
              reg429 <= reg230;
              reg430 <= (8'ha6);
              reg431 = (reg414[(1'h0):(1'h0)] >> (({(reg386 ~^ reg206),
                          (&reg370)} ?
                      reg287[(4'hc):(1'h0)] : reg416[(2'h3):(1'h1)]) ?
                  reg389 : {((~^reg249) ?
                          $signed(reg359) : wire350[(3'h6):(2'h2)]),
                      $unsigned(reg413)}));
              reg432 = (($signed((reg365 * (reg248 ? reg312 : reg400))) ?
                      reg245 : ($unsigned((reg428 ? reg199 : reg324)) ?
                          ($unsigned(reg232) & (wire195 && forvar363)) : (!reg313))) ?
                  $unsigned(reg355) : (^~forvar391));
            end
          reg433 = $signed((~$unsigned((reg413 ?
              (reg269 ? reg203 : reg392) : forvar419[(5'h15):(1'h1)]))));
          reg434 <= (~({{(reg385 >= (8'ha3)), (7'h41)}} <= {($unsigned(reg421) ?
                  (^~(8'ha8)) : reg346[(3'h4):(2'h3)])}));
          reg435 <= (|$unsigned(reg397[(2'h2):(1'h1)]));
        end
    end
  always
    @(posedge clk) begin
      if ({$signed(reg201[(4'ha):(3'h4)]),
          (((~reg293) << $unsigned($signed(reg313))) ?
              reg218[(5'h12):(4'hf)] : $unsigned((((8'ha2) || reg320) ?
                  reg341[(2'h2):(2'h2)] : {reg399, reg263, reg331})))})
        begin
          reg436 <= (reg258 ^ {$signed((reg365[(3'h5):(2'h3)] > (~|reg317)))});
          reg437 = $signed(((^reg362[(1'h1):(1'h0)]) ?
              $unsigned((&(7'h4d))) : {(reg312[(3'h7):(1'h0)] ?
                      (reg393 - reg280) : reg225[(5'h10):(4'hb)])}));
          if (((^~(reg243 ?
                  ((reg345 | reg215) ~^ (8'hb4)) : ((~&reg399) >= reg278))) ?
              (!($signed(reg429) > (+(reg424 | reg243)))) : reg245[(4'h9):(3'h4)]))
            begin
              reg438 <= {reg230, reg359[(1'h1):(1'h0)], $signed(reg416)};
            end
          else
            begin
              reg439 = reg402[(2'h3):(1'h0)];
              reg440 <= (!(~|reg256));
              reg441 = reg232;
              reg442 = $unsigned(reg439[(3'h7):(1'h0)]);
              reg443 = {($signed(reg441[(4'h9):(4'h8)]) ?
                      reg302[(4'hb):(4'h9)] : {$signed(((8'ha0) ?
                              reg341 : reg324))})};
              reg444 <= reg256;
              reg445 <= $signed((8'hbd));
            end
          reg446 <= reg439[(4'hf):(4'ha)];
          reg447 <= reg319[(1'h1):(1'h1)];
          if ((((~^$signed(reg283)) ?
                  ($unsigned($signed((8'hb5))) < (~reg236[(2'h3):(2'h2)])) : reg388) ?
              ((|(!(reg263 ^~ (8'hb4)))) ?
                  (($unsigned((8'h9d)) ?
                          $signed(reg441) : (reg389 <<< reg316)) ?
                      $unsigned($signed(reg441)) : $unsigned((|reg206))) : ((^(reg435 < reg273)) ~^ (+(|reg362)))) : reg201))
            begin
              reg448 = (reg243[(4'ha):(2'h3)] ?
                  reg399 : {$unsigned(reg263),
                      (-{{reg313}, (7'h4e)}),
                      ($signed(reg320) >= reg373[(2'h2):(1'h0)])});
              reg449 = reg313;
              reg450 = $signed(($unsigned($unsigned((reg258 ?
                  (8'hbe) : reg293))) <<< wire350));
              reg451 = $signed(reg324);
              reg452 = $signed($unsigned($unsigned((+(~^reg441)))));
              reg453 <= {$unsigned($signed((^~(reg416 <= reg265)))),
                  ($signed($signed($unsigned(reg208))) != ((&(reg403 + reg218)) ?
                      reg436[(4'h8):(3'h4)] : reg330[(3'h4):(2'h3)])),
                  $signed(reg430)};
              reg454 = reg312[(3'h5):(1'h0)];
            end
          else
            begin
              reg453 <= ((^$unsigned(($unsigned(reg359) || (reg278 ?
                  reg341 : reg444)))) == ({(!reg436)} * (7'h46)));
              reg454 = wire350[(4'he):(3'h5)];
              reg455 = (~^({reg206[(5'h10):(3'h4)], (|reg414)} | (^~(reg389 ?
                  (^~reg436) : (reg249 << reg313)))));
              reg456 <= (reg445[(4'hc):(4'ha)] || (!((&reg270[(1'h1):(1'h0)]) <= wire192)));
              reg457 = (((~^(reg376 <<< (8'ha4))) & reg280) >= (wire191 ?
                  {((+(7'h4f)) ?
                          $unsigned(reg283) : wire192)} : $unsigned(reg269[(4'he):(4'hc)])));
              reg458 = reg268;
              reg459 = $unsigned($signed((~^$signed((reg203 ?
                  reg442 : reg371)))));
            end
        end
      else
        begin
          if ($unsigned(reg210[(1'h1):(1'h1)]))
            begin
              reg437 = (($unsigned(((~^reg276) && (reg287 ?
                      (7'h4d) : reg343))) <<< reg370[(4'hd):(4'h9)]) ?
                  reg365[(1'h0):(1'h0)] : reg230[(5'h1a):(4'hc)]);
              reg438 <= (&reg216);
              reg439 = $unsigned(reg366[(3'h6):(2'h3)]);
              reg440 <= reg434[(5'h14):(4'hd)];
            end
          else
            begin
              reg437 = $unsigned($unsigned((reg371[(4'hb):(4'h9)] & ({(7'h58),
                  reg454} + reg370[(4'hc):(4'ha)]))));
              reg438 <= $signed($unsigned(wire193[(4'h8):(3'h7)]));
              reg440 <= $unsigned(((reg320 ?
                  $signed((reg268 || reg364)) : $unsigned($unsigned((7'h4b)))) && ({reg302[(3'h4):(2'h2)],
                      (reg319 ? reg383 : reg307),
                      ((8'ha3) ? reg434 : reg362)} ?
                  reg441 : ($unsigned((7'h4a)) ?
                      $signed(reg245) : reg284[(2'h2):(1'h0)]))));
              reg441 = {(reg386[(4'h9):(3'h6)] ?
                      $signed($unsigned((reg273 <<< reg424))) : ((~|(reg280 & reg245)) ?
                          $unsigned((+reg448)) : $unsigned(reg450[(4'hd):(3'h5)])))};
              reg442 = (~&((^($unsigned(reg402) >> reg331[(3'h4):(3'h4)])) == (($unsigned(reg284) ?
                      (reg450 | reg446) : $unsigned(reg278)) ?
                  ($signed(reg399) ? reg438 : (8'hac)) : reg424)));
              reg444 <= (((reg386 ^~ (reg230 ?
                      reg446[(3'h7):(1'h1)] : (reg429 | (8'ha6)))) >= (($signed((8'had)) ?
                          $unsigned(wire195) : (+reg341)) ?
                      (~|$unsigned(reg339)) : $signed($signed(reg442)))) ?
                  (reg245[(3'h6):(1'h0)] << reg237[(1'h0):(1'h0)]) : $unsigned(reg237));
              reg445 <= reg386[(1'h1):(1'h0)];
            end
          reg448 = reg321[(4'hc):(4'h9)];
          for (forvar449 = (1'h0); (forvar449 < (2'h3)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg450 = $signed((((^~{reg231}) & reg276[(2'h3):(1'h1)]) >> reg435));
              reg451 = (((~&reg270[(4'hc):(4'hc)]) || reg451[(4'hd):(1'h1)]) ?
                  reg245[(2'h2):(1'h1)] : (7'h54));
              reg452 = $signed(reg287[(5'h18):(4'ha)]);
              reg453 <= {(&$unsigned((+(~(7'h40))))),
                  ($signed(((~(8'hb6)) ^ ((8'hb4) << reg436))) ?
                      reg444[(5'h18):(4'ha)] : (((!reg244) ?
                          reg360[(4'h9):(4'h9)] : $unsigned((8'hbc))) >= (((7'h43) ?
                              (8'ha7) : reg259) ?
                          reg389[(1'h0):(1'h0)] : (!reg439))))};
              reg454 = (reg346 ~^ $signed(reg245[(4'ha):(3'h7)]));
              reg456 <= (reg398 ?
                  $unsigned((((reg284 >= reg249) << (reg447 ?
                      wire192 : reg278)) > $signed((reg366 ?
                      reg440 : reg205)))) : $signed($signed((+reg456[(5'h11):(1'h0)]))));
            end
          reg460 <= (+(wire192[(2'h3):(1'h0)] < ($unsigned(reg331[(3'h6):(3'h5)]) ?
              $unsigned((reg447 ? (7'h54) : reg237)) : $signed((-reg316)))));
        end
      for (forvar461 = (1'h0); (forvar461 < (3'h6)); forvar461 = (forvar461 + (1'h1)))
        begin
          reg462 <= (~($unsigned($signed((reg335 ? reg457 : (8'hbb)))) ?
              $signed($unsigned(reg430)) : ((~|reg225) || $signed(reg256[(5'h1b):(5'h12)]))));
          reg463 = $signed((+(forvar449 || reg302[(3'h5):(1'h1)])));
        end
      for (forvar464 = (1'h0); (forvar464 < (1'h1)); forvar464 = (forvar464 + (1'h1)))
        begin
          if ((((~$unsigned($unsigned(reg393))) ?
                  reg362[(3'h5):(1'h0)] : $signed((~|((7'h4c) >= wire191)))) ?
              (^~(7'h49)) : reg434[(5'h18):(4'h9)]))
            begin
              reg465 = {(8'ha8), reg331[(1'h0):(1'h0)]};
              reg466 = reg324[(5'h10):(3'h5)];
              reg467 = $signed({reg376,
                  reg203,
                  (((reg278 ? reg396 : reg441) ?
                          {reg269, reg465} : reg451[(4'hc):(4'hb)]) ?
                      reg321 : $signed($unsigned(reg335)))});
            end
          else
            begin
              reg465 = ((~&(8'ha4)) <<< $signed($unsigned($unsigned((wire191 ?
                  reg402 : reg434)))));
              reg468 <= {reg416};
              reg469 = ((-$signed({$unsigned(reg388)})) ?
                  (reg450 == reg312) : $signed(({(~|reg263),
                      (reg276 ?
                          (8'ha1) : reg300)} >>> $signed($unsigned((7'h4b))))));
              reg470 <= {$signed(reg366[(4'h8):(3'h5)]),
                  (^(({reg312, reg452, reg312} && reg259) * (~(~reg434))))};
              reg471 <= (~^(7'h46));
            end
          reg472 <= reg245[(5'h10):(4'hf)];
          for (forvar473 = (1'h0); (forvar473 < (3'h6)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 <= (~^$unsigned((reg227[(5'h17):(1'h0)] - reg302)));
            end
        end
      reg475 <= wire193[(5'h17):(2'h3)];
      if (wire191[(3'h5):(2'h3)])
        begin
          reg476 = reg339;
          if (({$unsigned($unsigned($signed(reg472)))} ?
              ($unsigned(wire193) ?
                  $signed($unsigned(((8'hba) ?
                      reg320 : reg345))) : (reg370[(4'hd):(3'h5)] < reg370[(4'he):(3'h5)])) : forvar473[(5'h11):(5'h10)]))
            begin
              reg477 = $signed(((+{$unsigned(reg316)}) ?
                  (($signed((7'h4e)) | $unsigned(reg459)) && (8'haa)) : (reg231 >> $unsigned(reg474))));
              reg478 = reg360[(5'h12):(4'hf)];
              reg479 = $unsigned({reg205[(4'hf):(1'h0)],
                  (reg445[(3'h5):(1'h0)] <= (!$unsigned(reg448))),
                  reg364});
              reg480 <= (7'h52);
              reg481 = (!$signed(($unsigned($signed(reg449)) >>> {((8'hb9) != (7'h56))})));
            end
          else
            begin
              reg477 = (~&$unsigned((8'hb8)));
              reg478 = (reg283 ?
                  (!$unsigned((~$unsigned(reg335)))) : reg402[(5'h12):(4'h8)]);
              reg480 <= $signed($signed(forvar473[(4'hc):(3'h7)]));
              reg481 = reg338;
              reg482 = $signed((~^reg435[(1'h1):(1'h0)]));
            end
          if (($unsigned((|{(~|reg338),
              $unsigned(reg312)})) || ((~^$unsigned(reg403)) | reg317[(2'h2):(2'h2)])))
            begin
              reg483 <= (&reg243);
              reg484 <= $unsigned(($unsigned(reg287) ?
                  (&$unsigned((|(8'hbd)))) : $signed($unsigned($unsigned(reg300)))));
              reg485 = (8'hab);
            end
          else
            begin
              reg485 = (+wire351);
              reg486 = (8'hae);
              reg487 = $unsigned((($signed(((7'h4e) ?
                  reg452 : reg466)) * ($unsigned(reg362) <<< reg284[(2'h2):(1'h0)])) > $signed({(reg479 ~^ reg388)})));
              reg488 = ({$signed(reg244),
                  $unsigned($unsigned(((8'ha1) <= reg421)))} + $signed((!({reg415,
                      (7'h4e)} ?
                  $signed(reg338) : (~|reg236)))));
              reg489 = {$signed($unsigned(((+(8'ha3)) ?
                      $signed(reg402) : (8'hbd)))),
                  ({wire192} <<< ($signed((reg360 ?
                      reg389 : reg479)) && ((reg472 & reg199) ?
                      reg218[(1'h1):(1'h1)] : (reg365 && reg478)))),
                  ((reg245 ~^ reg270) <<< reg360[(5'h18):(4'hf)])};
              reg490 <= $unsigned($unsigned((7'h40)));
              reg491 <= ({(~^(8'ha4))} || ($signed(reg446[(4'h8):(3'h5)]) ?
                  reg389 : (8'h9c)));
            end
          if ((|$unsigned($signed(((wire195 | (7'h53)) ?
              $unsigned(reg321) : (reg437 ? (7'h55) : wire190))))))
            begin
              reg492 <= $signed((reg403 <= reg205));
              reg493 <= $unsigned($signed((^~(reg280 ?
                  $signed(reg438) : $signed(reg231)))));
              reg494 <= $unsigned({($signed(reg421) * $unsigned($signed(wire195))),
                  $unsigned(reg481[(3'h7):(3'h4)])});
              reg495 = $signed($signed(((reg227 >>> reg482) ?
                  reg468 : $signed((^reg383)))));
              reg496 <= $signed($signed($signed($signed(reg398))));
              reg497 = {(reg455[(3'h5):(1'h0)] <<< reg434)};
            end
          else
            begin
              reg495 = {reg236[(4'h8):(2'h3)],
                  reg273[(4'he):(3'h6)],
                  (reg216[(5'h12):(4'he)] ?
                      wire195 : ($unsigned(reg339) ?
                          {((8'hb7) ? reg457 : reg376),
                              (reg256 ? wire350 : reg370)} : $signed((reg307 ?
                              reg414 : reg486))))};
              reg497 = $unsigned($unsigned((|reg389[(3'h6):(1'h0)])));
              reg498 = (8'had);
              reg499 = ({(+reg230[(1'h1):(1'h0)])} < (!$unsigned($signed($signed(reg386)))));
              reg500 = ({((7'h4b) ? reg388 : (^~{reg255, reg424, reg487})),
                      ((~&((8'hb2) ?
                          reg449 : reg438)) != (~^((8'had) ^~ reg475)))} ?
                  ({{$signed(reg287), reg416}} ?
                      $unsigned(reg402) : $signed(($unsigned(reg273) <<< $unsigned((8'haa))))) : (($signed({reg450,
                          reg276}) <<< reg489) ?
                      (^~((reg338 != reg252) ?
                          (reg458 ?
                              (8'haf) : reg345) : reg302)) : $signed(reg481[(1'h1):(1'h1)])));
              reg501 <= {reg477};
              reg502 <= reg300[(1'h0):(1'h0)];
            end
          reg503 <= forvar449;
        end
      else
        begin
          reg480 <= $signed($unsigned($signed(reg440[(1'h0):(1'h0)])));
        end
      for (forvar504 = (1'h0); (forvar504 < (1'h1)); forvar504 = (forvar504 + (1'h1)))
        begin
          reg505 <= reg280;
          for (forvar506 = (1'h0); (forvar506 < (2'h2)); forvar506 = (forvar506 + (1'h1)))
            begin
              reg507 <= reg463[(4'hd):(3'h7)];
              reg508 = (reg218[(2'h3):(1'h0)] ?
                  $unsigned((reg269[(3'h6):(3'h6)] ?
                      reg312 : ($signed(wire190) ?
                          reg311[(5'h15):(4'h9)] : (reg206 <= (8'hbd))))) : ($signed(($unsigned(reg284) ?
                      $unsigned(reg507) : {(8'hb6),
                          (7'h4b),
                          reg445})) ^ $signed($signed((~wire192)))));
              reg509 <= (8'ha0);
              reg510 = reg269[(4'h8):(3'h6)];
              reg511 <= reg430[(3'h4):(2'h2)];
            end
          if ((|({($unsigned(reg458) >>> (reg339 & reg495))} ?
              reg475 : reg489[(3'h6):(1'h0)])))
            begin
              reg512 <= $signed({(reg393 & forvar464[(5'h19):(2'h3)]),
                  $unsigned((~^reg206[(3'h5):(3'h4)]))});
              reg513 <= $signed($signed($unsigned(($signed(reg203) ~^ reg434))));
              reg514 <= (&($signed($signed(reg398[(3'h5):(1'h0)])) ^ (~^reg415[(3'h5):(2'h3)])));
              reg515 <= (reg480[(5'h19):(5'h18)] > $unsigned(((~|$unsigned((8'hbf))) && {reg365[(2'h3):(1'h1)]})));
            end
          else
            begin
              reg512 <= ($unsigned(reg480[(4'hb):(4'h8)]) ?
                  ($signed(($signed(reg483) == reg467)) ?
                      $signed(($unsigned(reg203) ~^ reg440)) : ($unsigned($signed(reg421)) ?
                          $unsigned($unsigned(reg366)) : reg439[(4'he):(4'hd)])) : (^$unsigned(reg270)));
              reg513 <= (~^({((reg216 + reg259) <= reg307),
                      reg269[(5'h16):(3'h6)],
                      $unsigned($signed(reg244))} ?
                  (^~reg416) : $unsigned(reg399[(3'h5):(3'h4)])));
            end
        end
    end
  assign wire516 = $signed($signed(reg244));
  module517 #() modinst585 (.wire518(reg460), .wire521(reg483), .wire519(reg311), .wire520(reg440), .clk(clk), .y(wire584));
  always
    @(posedge clk) begin
      if ({reg370})
        begin
          if (reg503)
            begin
              reg586 = $signed(((8'hbb) | (reg208[(1'h0):(1'h0)] <<< (^reg366))));
            end
          else
            begin
              reg587 <= {(8'ha9)};
            end
          if ({{(reg258 ^ ({reg216, reg321} || (wire195 ? (7'h4a) : (8'had)))),
                  ((-(reg365 * (8'ha7))) ?
                      (-{reg256, (8'hb7), reg393}) : (reg371[(4'hf):(4'hf)] ?
                          reg335 : reg270)),
                  $unsigned({(8'hab), reg514, reg284[(2'h2):(2'h2)]})},
              $unsigned(reg248[(3'h5):(2'h2)])})
            begin
              reg588 = reg228;
              reg589 <= $signed(($signed((~&reg255)) <<< ($signed((reg493 << reg339)) >> $unsigned($unsigned((8'ha9))))));
              reg590 = wire351[(4'hf):(4'hc)];
              reg591 <= ({reg365[(4'ha):(3'h5)],
                  (^(~|(reg370 ? reg513 : reg227))),
                  reg480[(5'h15):(5'h12)]} <= (^$signed((reg430[(5'h15):(3'h7)] != (~&reg396)))));
            end
          else
            begin
              reg589 <= reg273;
              reg590 = {(reg438[(4'hc):(3'h6)] == $unsigned($unsigned(reg396[(3'h5):(1'h1)])))};
              reg591 <= $unsigned($unsigned(reg324[(4'hf):(2'h3)]));
              reg592 <= {$unsigned(wire194[(5'h15):(4'h8)]),
                  wire191[(3'h7):(3'h6)],
                  (wire195 ?
                      ({$signed(reg331), (+reg270), reg216[(3'h4):(2'h2)]} ?
                          (8'hac) : (|$unsigned(reg460))) : $unsigned($signed({(7'h40),
                          (8'hb5)})))};
            end
          reg593 <= (($signed(reg592) & (^~(reg300 ?
              $unsigned(reg429) : $unsigned(reg210)))) * $signed({{(!reg249),
                  $unsigned(reg312),
                  wire351[(3'h6):(2'h3)]},
              $signed({reg587}),
              $signed(((8'haa) ? reg591 : reg259))}));
        end
      else
        begin
          if ($signed((8'h9c)))
            begin
              reg587 <= reg366[(4'hd):(4'h8)];
              reg589 <= {{(($signed(reg225) ^ (^reg265)) > reg429)},
                  $unsigned((reg590 == ($signed(wire190) ?
                      reg276[(1'h0):(1'h0)] : (~|(7'h54))))),
                  $signed((reg331[(4'he):(1'h0)] ?
                      {(+reg471),
                          (^~(8'h9f)),
                          $unsigned(reg273)} : $unsigned(wire192[(1'h0):(1'h0)])))};
              reg590 = ((~|reg588) ?
                  ((^~reg446[(2'h3):(2'h3)]) ?
                      $unsigned((!reg321)) : reg592) : ((~|(((8'hb2) ?
                              reg346 : reg511) ?
                          $unsigned(reg238) : (~reg232))) ?
                      (|reg507[(4'hf):(1'h1)]) : reg206));
              reg591 <= reg393;
              reg594 = ((reg311 ?
                      (~&reg424) : ($signed(reg389) <<< (reg218 ?
                          (^~reg335) : $unsigned(reg256)))) ?
                  (+({(reg444 & reg456)} ?
                      (!$signed(reg480)) : $signed((wire584 >= reg399)))) : $unsigned(((((8'hbc) ?
                          reg276 : (8'ha6)) ?
                      (+reg502) : reg216) != ((reg302 ?
                      reg456 : reg339) <= $unsigned(reg388)))));
              reg595 = reg201;
              reg596 = (reg398[(2'h2):(2'h2)] && (reg456[(1'h0):(1'h0)] < (7'h4e)));
            end
          else
            begin
              reg586 = (~reg462[(1'h0):(1'h0)]);
              reg588 = (reg284 > reg276);
              reg590 = (reg216[(3'h5):(2'h2)] ?
                  ($unsigned((~&reg383[(5'h15):(5'h11)])) ^ $signed($unsigned((reg263 < reg512)))) : $signed((reg589 ?
                      (reg370 < reg396[(3'h6):(3'h4)]) : reg238[(2'h3):(1'h0)])));
              reg594 = $unsigned(reg293);
            end
          reg597 <= ((|$unsigned(reg208[(1'h1):(1'h0)])) ^~ reg278);
          for (forvar598 = (1'h0); (forvar598 < (3'h6)); forvar598 = (forvar598 + (1'h1)))
            begin
              reg599 = $signed(reg330);
            end
        end
      if ($signed($unsigned(((~(7'h51)) ^~ ((reg586 - reg490) ?
          $signed(wire350) : $unsigned(reg588))))))
        begin
          reg600 <= (7'h47);
          reg601 = reg270;
        end
      else
        begin
          reg600 <= $signed((&($unsigned($signed(reg472)) ?
              ((~^reg414) ?
                  {reg215, reg248} : (reg346 == reg490)) : $signed(reg501))));
          reg602 <= (($unsigned((~|(~^reg248))) ~^ (($unsigned((8'hb0)) ^ reg396) <<< reg453[(3'h6):(2'h2)])) ?
              reg215[(3'h6):(1'h1)] : (reg507 >>> (((reg491 ?
                          (7'h47) : reg312) ?
                      reg588[(3'h4):(2'h2)] : $signed((8'haf))) ?
                  $unsigned((reg445 ? reg283 : reg313)) : {reg493,
                      reg330,
                      {reg460}})));
          for (forvar603 = (1'h0); (forvar603 < (2'h3)); forvar603 = (forvar603 + (1'h1)))
            begin
              reg604 <= $signed({(reg493 ?
                      ({reg471, (8'haa), wire516} ?
                          ((8'h9c) ? reg586 : (8'hbc)) : (reg492 ?
                              reg376 : reg430)) : $unsigned($signed(reg218))),
                  reg484[(2'h2):(1'h1)]});
              reg605 = $signed((((8'h9f) ?
                  (^(reg593 ^ reg475)) : (-reg393)) > reg263[(1'h0):(1'h0)]));
              reg606 <= ((^~((~&reg324) ?
                      {{reg365, (8'hb7), reg203}, reg330} : {(wire191 ?
                              reg386 : reg208)})) ?
                  reg263 : {$signed(reg511[(2'h3):(1'h0)]), reg231});
              reg607 <= (8'hb1);
              reg608 = $signed((((|(reg602 | reg216)) ~^ reg444[(4'ha):(4'ha)]) - (~|reg311[(4'hc):(3'h5)])));
            end
          if (reg230)
            begin
              reg609 = $signed(($signed($signed($signed(reg396))) ?
                  {reg438[(3'h7):(1'h1)],
                      ($unsigned(reg216) ?
                          ((8'h9e) >= reg210) : reg255[(1'h0):(1'h0)])} : (reg474 ?
                      ((reg608 ? reg513 : reg330) ?
                          $signed(reg283) : (reg218 >= reg238)) : (((7'h45) || reg453) <= (reg430 * reg511)))));
              reg610 <= reg609[(1'h0):(1'h0)];
              reg611 = wire191[(4'hc):(1'h1)];
              reg612 <= (reg376 ^~ (($unsigned({reg330}) >>> reg339[(4'hf):(4'hc)]) <= reg503[(4'h8):(1'h0)]));
              reg613 <= (!{({((8'hae) ? reg215 : reg243),
                      (8'hb4)} == $unsigned($unsigned((8'hab))))});
            end
          else
            begin
              reg610 <= $signed($signed($unsigned((^(-reg270)))));
              reg611 = reg256;
              reg612 <= $signed(((~(+(reg468 ?
                  reg252 : reg371))) * (~(7'h44))));
              reg614 = reg227;
              reg615 = (^~{{reg447,
                      reg319[(2'h3):(1'h0)],
                      $signed($signed(reg607))},
                  (+((8'hb7) && reg236[(3'h5):(3'h5)]))});
            end
          if (reg512[(5'h11):(5'h11)])
            begin
              reg616 <= (({(((8'haf) ?
                          (8'hab) : reg480) - $signed(reg474))} & $unsigned(reg365)) ?
                  $signed(((~^reg359) + reg597)) : $unsigned(($signed((wire584 ?
                          reg269 : reg210)) ?
                      $signed((^~reg610)) : ((reg614 ? reg460 : reg225) ?
                          {reg613} : reg606[(2'h2):(1'h0)]))));
              reg617 <= $signed(reg273);
              reg618 <= reg610[(5'h14):(5'h10)];
              reg619 <= {reg396[(4'hc):(1'h1)]};
            end
          else
            begin
              reg616 <= (^(|((~^(|reg589)) && ((~^reg365) ?
                  (reg321 ? wire350 : reg607) : {reg258, reg445}))));
            end
        end
      reg620 <= ($signed(($unsigned((wire195 - reg269)) ?
              reg599[(5'h16):(4'he)] : (reg424 <= $unsigned(reg311)))) ?
          $unsigned((((!reg587) ?
              reg430[(4'he):(4'he)] : {reg490}) & $unsigned((|reg330)))) : reg456[(3'h4):(1'h0)]);
      reg621 = reg591;
      if (((&$unsigned(reg259[(3'h4):(1'h0)])) ?
          (7'h41) : $signed($signed($unsigned((^reg270))))))
        begin
          for (forvar622 = (1'h0); (forvar622 < (2'h3)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 = (-((reg492 << reg307) ?
                  $unsigned((~&$unsigned((8'ha6)))) : ((~^reg468) ?
                      (~^$signed(reg263)) : (-(reg203 ? reg594 : reg605)))));
              reg624 <= $signed($signed(reg612[(4'he):(3'h4)]));
              reg625 = reg359[(1'h1):(1'h0)];
              reg626 = ({reg416[(2'h3):(1'h1)],
                      $signed((reg341[(2'h3):(1'h0)] ? reg283 : (~forvar603))),
                      ($signed((!reg280)) < ((~&wire516) && (~^forvar598)))} ?
                  $unsigned(reg502) : reg496);
              reg627 <= reg609[(4'h9):(3'h7)];
              reg628 = (reg611[(4'he):(3'h5)] ?
                  $signed($signed(reg206)) : (~^$signed(($unsigned((8'hb7)) ?
                      reg364[(1'h1):(1'h0)] : $signed((7'h4c))))));
            end
          if (reg245)
            begin
              reg629 = $signed((&(~&reg424[(4'he):(3'h6)])));
              reg630 = reg243[(2'h3):(1'h1)];
              reg631 = $signed(reg429[(3'h4):(1'h1)]);
              reg632 = $unsigned({reg494[(5'h16):(4'hb)]});
              reg633 = (&(reg225[(5'h10):(3'h6)] ?
                  reg447 : {((~^(8'hbf)) >= (-reg364))}));
            end
          else
            begin
              reg629 = $unsigned($unsigned(reg317[(2'h2):(1'h0)]));
              reg634 <= (~|($unsigned((~^(reg238 ? (7'h4c) : reg293))) ?
                  reg480 : $signed($unsigned((reg588 >= reg515)))));
            end
          reg635 <= reg446[(3'h7):(1'h0)];
          if (reg255)
            begin
              reg636 <= $unsigned(((((|reg307) ?
                  ((8'ha7) != reg388) : reg238[(2'h2):(2'h2)]) - (wire350[(4'ha):(2'h2)] ?
                  $signed(forvar622) : (reg618 ^~ reg218))) >= reg300[(1'h0):(1'h0)]));
              reg637 = (reg362 >= ($signed($signed((reg324 ?
                  reg623 : reg362))) | $unsigned($signed({reg636,
                  reg252,
                  reg608}))));
              reg638 <= (!(!{$unsigned((&reg225))}));
              reg639 <= $unsigned((7'h42));
            end
          else
            begin
              reg637 = {reg208[(1'h1):(1'h0)],
                  (reg383 | (((~^(8'hb8)) ? (&(7'h48)) : (!reg201)) ?
                      ((8'hb0) ?
                          (~^(8'hb7)) : reg493[(4'h8):(1'h0)]) : {(reg609 - reg258)})),
                  {$signed((reg276[(3'h4):(2'h2)] ?
                          (~&reg383) : (wire584 ^~ reg619)))}};
              reg638 <= reg496;
              reg640 = reg225;
              reg641 <= $signed($unsigned(reg509[(5'h1a):(4'he)]));
              reg642 = ($unsigned({($unsigned(reg592) ?
                          $unsigned(reg496) : {reg615, reg383, reg244}),
                      (~(wire190 ? reg609 : reg610))}) ?
                  reg364[(2'h2):(1'h1)] : $unsigned(reg507[(4'ha):(1'h0)]));
              reg643 <= reg634;
              reg644 = $signed($signed($signed((~|reg396))));
            end
          reg645 <= (8'hae);
          reg646 <= $unsigned({$unsigned(($unsigned(reg231) ?
                  (^(7'h44)) : $unsigned(reg604))),
              reg293});
          if (reg203)
            begin
              reg647 = reg602;
              reg648 <= ((reg589[(5'h12):(5'h12)] ?
                      $signed(reg237) : {(~$signed(reg604))}) ?
                  (&{$signed((~|(7'h48)))}) : (((reg346 ~^ reg587[(4'h8):(1'h1)]) ?
                      ($signed(reg316) << (~&wire351)) : {(^reg227),
                          (!reg470),
                          (wire351 && reg635)}) ~^ {$signed(reg273[(4'hd):(2'h3)]),
                      (&$unsigned(reg480))}));
              reg649 <= {$signed(reg421),
                  $signed(((^$unsigned(reg312)) ?
                      ((reg601 ? reg496 : reg252) ?
                          $signed(reg393) : {reg238}) : reg609)),
                  $signed(reg370)};
              reg650 <= reg599;
              reg651 = (-$unsigned($unsigned(reg616[(1'h0):(1'h0)])));
            end
          else
            begin
              reg648 <= (7'h43);
            end
        end
      else
        begin
          reg622 = forvar622;
          if ($signed((~{$unsigned((reg456 ? (7'h42) : reg638))})))
            begin
              reg624 <= (^(((^~$signed(reg647)) && (~&(wire516 ?
                  reg633 : reg421))) || reg512));
              reg627 <= (~$signed(reg249));
              reg634 <= $unsigned($unsigned({reg320,
                  $unsigned($unsigned(reg421))}));
              reg637 = (7'h41);
              reg638 <= (^{reg480[(4'hd):(4'ha)], reg626[(5'h15):(5'h14)]});
              reg640 = ((reg276[(1'h1):(1'h1)] ?
                  {$signed((-(7'h4b))),
                      ((reg248 ~^ (7'h4b)) ? (reg307 << reg453) : reg468),
                      (^(reg331 ?
                          reg492 : reg436))} : ($unsigned($signed(reg474)) >>> reg421[(1'h0):(1'h0)])) ^~ {(&wire584),
                  $unsigned(((reg629 ? reg636 : reg398) ?
                      (!reg444) : $signed(reg208))),
                  (|{$signed(reg632)})});
              reg641 <= ($unsigned((($signed(reg593) >>> $unsigned(reg265)) - (~&(+(7'h51))))) & (~|$signed((8'haf))));
            end
          else
            begin
              reg623 = $signed(reg496);
              reg624 <= (reg646 >>> {$signed(((~&reg216) ?
                      $unsigned(reg456) : reg327)),
                  wire191});
              reg627 <= $signed({reg490});
              reg628 = $signed($signed((~^(8'ha3))));
              reg629 = $unsigned(($signed(((7'h52) + reg493[(4'hc):(3'h6)])) ?
                  $unsigned((~|reg650)) : reg429[(2'h2):(2'h2)]));
            end
          reg643 <= $unsigned($unsigned(((-reg230[(4'he):(3'h6)]) || ($unsigned(reg642) ^~ reg243[(2'h2):(2'h2)]))));
          reg645 <= (reg287[(5'h11):(4'hf)] ?
              $unsigned(((!(^~reg263)) <<< ((reg644 || reg601) ^~ (|reg494)))) : (($signed((!(8'ha3))) ?
                      $unsigned((reg435 ? reg484 : reg624)) : reg593) ?
                  reg396[(4'hf):(4'hc)] : (|$signed((~reg228)))));
          if (reg484[(2'h3):(1'h0)])
            begin
              reg646 <= (reg605[(5'h1f):(5'h1e)] ?
                  reg415 : $signed((((reg595 ? (7'h54) : reg593) ?
                      $signed(reg447) : (~|reg453)) * reg629[(5'h15):(4'h9)])));
              reg648 <= (reg592[(2'h2):(1'h0)] <= (|$unsigned($signed(wire192))));
              reg649 <= reg588;
            end
          else
            begin
              reg647 = reg389[(2'h2):(2'h2)];
            end
          for (forvar650 = (1'h0); (forvar650 < (2'h2)); forvar650 = (forvar650 + (1'h1)))
            begin
              reg652 <= (($signed($unsigned(reg278[(1'h1):(1'h1)])) > $signed((8'hb9))) ?
                  (|wire192[(2'h2):(1'h1)]) : reg588[(1'h1):(1'h1)]);
            end
          if ((({$signed($signed(reg327))} || (+$signed((-reg210)))) ?
              reg430[(3'h7):(2'h3)] : reg606[(2'h3):(2'h2)]))
            begin
              reg653 <= reg268;
              reg654 <= (reg416[(4'h9):(4'h8)] ?
                  reg590[(4'h9):(4'h8)] : ($unsigned($unsigned({reg302,
                          reg237,
                          reg460})) ?
                      (((^reg623) & (reg607 ^~ reg388)) ?
                          ((reg313 ?
                              (8'ha1) : reg642) ^~ $signed(reg589)) : (~$unsigned(reg438))) : $signed((reg638 ?
                          forvar598[(3'h5):(3'h4)] : reg503))));
              reg655 <= (~|reg248[(3'h5):(2'h2)]);
              reg656 = $unsigned($unsigned(($signed((reg483 ?
                      reg203 : reg343)) ?
                  reg642 : ((~&reg338) ?
                      $unsigned(reg639) : reg446[(2'h2):(1'h0)]))));
              reg657 <= reg609[(4'h9):(4'h9)];
              reg658 = reg509;
            end
          else
            begin
              reg653 <= $signed(((reg236 ~^ ($signed(reg492) == (reg648 || reg625))) * $signed((+reg639[(4'h9):(3'h4)]))));
              reg656 = $signed($unsigned((reg514[(5'h1c):(5'h1a)] & $signed((-reg414)))));
              reg657 <= reg490[(2'h2):(1'h0)];
              reg658 = (reg416[(1'h0):(1'h0)] < reg293[(3'h4):(1'h1)]);
              reg659 <= ($signed((-$signed(reg255[(2'h2):(1'h1)]))) ?
                  $unsigned($unsigned($unsigned(reg640[(4'h9):(1'h1)]))) : ((~&{(~|wire350),
                          $unsigned(reg278),
                          (~|reg635)}) ?
                      reg602 : $unsigned($signed({reg414}))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar660 = (1'h0); (forvar660 < (2'h3)); forvar660 = (forvar660 + (1'h1)))
        begin
          for (forvar661 = (1'h0); (forvar661 < (1'h1)); forvar661 = (forvar661 + (1'h1)))
            begin
              reg662 = ((~|(((reg472 ?
                  reg371 : reg502) | (reg655 ^ (8'hbe))) >>> ((~&reg319) != $unsigned(reg445)))) >= $signed(reg429[(2'h2):(1'h0)]));
              reg663 <= $unsigned(reg312[(3'h6):(3'h5)]);
              reg664 <= reg218;
              reg665 = (^~reg205[(3'h5):(3'h5)]);
              reg666 = $unsigned(((({(8'hb1), (7'h57)} ?
                  $unsigned(wire192) : (reg424 ?
                      reg359 : reg509)) >= ($signed(reg339) <= $signed(reg343))) + ((wire193 != (~&reg645)) ?
                  (reg606 <= $unsigned(reg307)) : (!$signed(reg393)))));
              reg667 <= (~&$signed(reg228));
              reg668 = ((-reg587[(4'he):(4'hb)]) + (|$signed((^$signed(reg511)))));
            end
          reg669 <= ({(8'hac)} > {(reg258 ?
                  reg258[(1'h0):(1'h0)] : (!reg321[(1'h0):(1'h0)])),
              $unsigned((reg502 ? reg610 : (reg653 ? reg339 : reg320))),
              (7'h44)});
          for (forvar670 = (1'h0); (forvar670 < (2'h3)); forvar670 = (forvar670 + (1'h1)))
            begin
              reg671 <= reg421;
              reg672 <= $signed(((reg470 ?
                      (reg320[(5'h1b):(5'h1a)] ?
                          $unsigned(reg649) : (reg327 | (8'hb4))) : (|wire195)) ?
                  ((&(|reg259)) ?
                      reg299 : ($unsigned((7'h53)) ^~ $signed(wire195))) : ((((7'h56) ?
                          reg386 : reg345) ?
                      reg287[(5'h15):(4'h9)] : reg245) || (+(reg462 <= reg366)))));
              reg673 <= reg249;
              reg674 <= $signed($unsigned((((~|(8'ha1)) ?
                  (&reg472) : (reg657 ^~ reg610)) | (~^$unsigned(reg203)))));
              reg675 <= $signed($signed(($signed((~reg618)) ^~ reg496[(4'hb):(3'h5)])));
              reg676 = reg270;
              reg677 = $signed(reg346);
            end
          reg678 <= $unsigned((reg462[(3'h5):(2'h2)] ?
              ((reg208[(1'h1):(1'h0)] ~^ (~(7'h53))) & $unsigned(reg616)) : reg203));
          for (forvar679 = (1'h0); (forvar679 < (1'h0)); forvar679 = (forvar679 + (1'h1)))
            begin
              reg680 = $unsigned($signed((!((^~(7'h42)) && $signed(reg662)))));
              reg681 = ($signed($unsigned(reg299)) > $signed((reg515[(1'h1):(1'h0)] & $signed(((8'hbb) ?
                  reg268 : reg666)))));
              reg682 = ((!$unsigned(((^reg263) ^~ (!reg346)))) ?
                  (reg316[(3'h4):(1'h0)] <= (7'h4b)) : $signed({{(^~reg316),
                          $signed(reg591),
                          (~|(8'hb5))},
                      (~&$unsigned(reg501))}));
              reg683 <= (8'hb4);
              reg684 = (|reg512[(4'ha):(1'h0)]);
            end
          reg685 = ($signed(((-reg468) ? reg256[(2'h2):(2'h2)] : (8'hbe))) ?
              (!(({reg430, reg667} ?
                      (reg227 ? reg515 : reg612) : (reg654 ? reg638 : reg669)) ?
                  reg606 : ((reg641 ? (8'ha3) : reg330) ?
                      (|reg639) : (reg300 ?
                          (8'hbc) : reg472)))) : (reg675[(1'h0):(1'h0)] >>> ((reg339[(3'h6):(3'h5)] * (reg265 ?
                  reg494 : reg330)) < $signed({reg225, reg681}))));
          if ($signed((+$unsigned(reg606[(2'h2):(2'h2)]))))
            begin
              reg686 = (7'h40);
              reg687 = $signed($signed((+(reg668 ?
                  {reg683, reg446, reg592} : (wire350 || reg639)))));
            end
          else
            begin
              reg688 <= reg256;
              reg689 <= ((!$signed($unsigned($unsigned((8'ha2))))) ?
                  (reg682[(4'h9):(3'h6)] || reg228[(4'hd):(1'h1)]) : forvar670[(3'h4):(2'h3)]);
              reg690 = $unsigned(((((+reg373) ~^ $signed(reg284)) ?
                  $signed($signed(reg436)) : $unsigned((reg396 > reg447))) || (reg258[(2'h2):(1'h1)] ?
                  (-((8'h9f) * reg327)) : ((-reg307) ?
                      reg650 : $signed(reg245)))));
            end
        end
      reg691 = ((reg453[(1'h1):(1'h1)] || $unsigned($unsigned((reg674 ?
          reg593 : reg634)))) >>> $signed(reg634));
      if ($signed(forvar670))
        begin
          if ({{reg592}, reg210[(2'h2):(2'h2)]})
            begin
              reg692 = reg480;
            end
          else
            begin
              reg692 = (7'h53);
              reg693 <= (^~reg593);
              reg694 = reg496;
              reg695 = $signed(($signed(reg460[(3'h6):(3'h5)]) ?
                  $signed($signed($unsigned(reg668))) : $unsigned(reg201)));
              reg696 <= reg273[(4'h9):(3'h6)];
              reg697 = reg675[(4'ha):(3'h7)];
              reg698 <= {reg676,
                  ((reg645 ?
                          reg345 : ((7'h49) ?
                              (reg421 >= wire190) : (!reg293))) ?
                      (((reg483 >>> reg687) >>> reg618[(3'h7):(2'h3)]) != ((^~reg343) ?
                          $unsigned(reg693) : (~reg681))) : {{((8'hb5) & reg462),
                              $signed(wire516)},
                          $unsigned((reg624 ? reg689 : reg624))}),
                  {{reg493,
                          ($signed(reg245) ?
                              reg493 : (reg686 ? reg255 : reg617)),
                          ($signed((7'h56)) >> $unsigned(reg447))},
                      $signed($unsigned(reg634))}};
            end
          if ((&(7'h53)))
            begin
              reg699 <= reg503;
              reg700 <= ($unsigned(reg278[(5'h1f):(4'hb)]) == ((!(~^{reg341,
                      reg269,
                      reg312})) ?
                  {reg205[(3'h4):(1'h0)]} : (+reg502[(4'ha):(4'h9)])));
              reg701 = ($signed(reg366[(4'h8):(3'h6)]) ?
                  $unsigned({$signed((reg494 << reg415)),
                      (7'h44)}) : {($signed({reg335}) ?
                          $unsigned(reg635[(3'h4):(2'h3)]) : {$unsigned(reg210),
                              (-reg700),
                              $signed(reg430)})});
              reg702 <= reg515[(4'h8):(4'h8)];
              reg703 <= $unsigned($unsigned((~&$unsigned($unsigned(reg434)))));
              reg704 <= (+reg208[(1'h1):(1'h0)]);
              reg705 <= ((^$unsigned((-$signed((8'ha1))))) == reg503[(5'h10):(5'h10)]);
            end
          else
            begin
              reg701 = {{(+$unsigned((reg600 > reg509))),
                      {reg671, (reg513[(1'h1):(1'h0)] >= (reg619 | reg444))},
                      (reg673 ?
                          $signed((reg389 ?
                              reg302 : reg659)) : ({reg698} || reg513))},
                  ($signed((!$unsigned(reg362))) ? (7'h45) : (8'hb6))};
              reg702 <= $signed(reg694[(3'h6):(1'h0)]);
              reg703 <= reg320;
              reg706 = reg199[(5'h15):(2'h3)];
              reg707 <= reg686;
              reg708 <= ($signed(reg483[(1'h0):(1'h0)]) ?
                  (~&$unsigned((~$signed(reg701)))) : (($unsigned(((7'h47) ?
                      reg364 : reg435)) <<< $unsigned((reg687 * reg646))) != reg203[(5'h11):(3'h4)]));
              reg709 <= (~^$unsigned((|($unsigned((8'ha4)) ?
                  (~reg591) : (~&reg389)))));
            end
          reg710 = $signed($signed(reg268[(2'h3):(1'h0)]));
          if ((~&($unsigned(reg600) ^ reg699[(4'he):(4'h9)])))
            begin
              reg711 = (&$unsigned(reg360));
              reg712 = ($signed(reg512[(5'h15):(4'hb)]) ?
                  (reg430[(1'h1):(1'h1)] ?
                      (reg604[(5'h13):(1'h1)] ?
                          ($signed(reg667) ^~ reg702[(3'h6):(1'h1)]) : reg494) : (reg376[(1'h1):(1'h0)] ?
                          (reg338 ?
                              $unsigned(reg456) : (|reg203)) : $unsigned($signed(reg360)))) : {($signed($signed(reg228)) << ((&reg475) ?
                          (~reg512) : $signed(reg255)))});
            end
          else
            begin
              reg711 = reg677[(5'h12):(5'h11)];
              reg713 <= {reg307[(3'h6):(2'h3)], {$signed(reg273)}};
              reg714 = reg319[(3'h4):(1'h0)];
              reg715 = $signed($signed(reg402));
            end
          reg716 = (^$signed($unsigned(($signed((8'haa)) >= reg610[(2'h2):(1'h0)]))));
        end
      else
        begin
          reg692 = (!(reg667[(1'h0):(1'h0)] && {(reg313 + $signed((7'h43)))}));
          reg693 <= $unsigned(reg232[(1'h0):(1'h0)]);
        end
    end
  assign wire717 = $unsigned($signed({(((8'ha5) <= reg386) ?
                           $signed(reg438) : {reg265, reg591}),
                       (~(reg689 <= reg704))}));
  assign wire718 = ($unsigned((8'ha6)) >>> wire584);
  always
    @(posedge clk) begin
      reg719 = reg468[(4'he):(4'hb)];
      reg720 = reg446;
      reg721 = $signed($unsigned($signed(reg616[(2'h2):(1'h0)])));
      for (forvar722 = (1'h0); (forvar722 < (3'h4)); forvar722 = (forvar722 + (1'h1)))
        begin
          reg723 = $unsigned({(~(+$unsigned(wire195)))});
          reg724 <= reg434;
          if ((&reg678[(1'h0):(1'h0)]))
            begin
              reg725 = reg343[(4'ha):(3'h5)];
              reg726 <= (|$signed(reg263));
              reg727 <= ($unsigned((8'hb5)) ?
                  (reg646[(3'h6):(3'h5)] > reg664) : {reg225,
                      reg284[(2'h3):(2'h2)],
                      reg376});
              reg728 <= (&$signed($signed((+(-(8'ha5))))));
              reg729 = $unsigned(($signed(reg659) && (8'hba)));
              reg730 <= reg389;
              reg731 <= $unsigned(($unsigned(reg230[(4'hb):(3'h7)]) >>> ((!(7'h49)) ?
                  ($unsigned((7'h4d)) <= reg720[(4'h8):(3'h5)]) : {{reg649,
                          reg612,
                          reg688}})));
            end
          else
            begin
              reg726 <= $signed(((!(&$unsigned(reg341))) ?
                  ({reg597[(1'h0):(1'h0)],
                          $signed(reg316),
                          (reg698 ? reg726 : reg468)} ?
                      ($signed(reg434) == {reg713,
                          reg327,
                          reg619}) : reg445) : {reg511[(5'h13):(3'h6)]}));
            end
          for (forvar732 = (1'h0); (forvar732 < (1'h0)); forvar732 = (forvar732 + (1'h1)))
            begin
              reg733 = $unsigned(wire193[(2'h2):(1'h1)]);
              reg734 <= reg447;
              reg735 = ($signed($signed($unsigned($signed(reg484)))) ?
                  (reg362[(2'h2):(1'h0)] * reg338) : (^~(reg653[(3'h4):(1'h0)] <<< (reg346 ?
                      (wire192 ? reg341 : reg225) : $signed((8'hbc))))));
              reg736 <= reg245[(5'h12):(3'h7)];
              reg737 = reg435;
              reg738 = (~($signed($signed($signed(wire190))) < $signed(($unsigned(reg429) == reg388[(2'h2):(2'h2)]))));
              reg739 = $unsigned($unsigned((^~{$unsigned(reg730), reg208})));
            end
          for (forvar740 = (1'h0); (forvar740 < (1'h1)); forvar740 = (forvar740 + (1'h1)))
            begin
              reg741 <= $unsigned((~^(((reg237 ?
                      reg256 : reg491) ~^ (reg318 <= reg280)) ?
                  $unsigned((7'h56)) : $signed(((8'hb4) ? reg513 : reg429)))));
              reg742 <= (reg399[(5'h14):(5'h10)] ?
                  $signed((&reg735[(1'h1):(1'h0)])) : reg238);
            end
        end
      for (forvar743 = (1'h0); (forvar743 < (3'h6)); forvar743 = (forvar743 + (1'h1)))
        begin
          reg744 <= reg341[(3'h4):(1'h1)];
          reg745 <= ($signed($signed(reg483)) ?
              (($unsigned(((8'hbf) ^~ reg201)) << (reg307 || reg672[(3'h7):(1'h1)])) ?
                  $signed((!$unsigned((8'h9f)))) : $signed($unsigned({reg383}))) : {$unsigned($unsigned($unsigned(reg311))),
                  reg602,
                  $unsigned((reg269 ? {reg373} : (reg652 ? reg737 : reg227)))});
          for (forvar746 = (1'h0); (forvar746 < (2'h2)); forvar746 = (forvar746 + (1'h1)))
            begin
              reg747 <= (7'h45);
              reg748 = (~(reg744[(2'h2):(1'h0)] + ($signed((reg678 - wire193)) * ((wire194 ?
                  reg327 : (7'h51)) && (wire718 == reg475)))));
              reg749 = (reg399[(1'h1):(1'h1)] > reg341[(2'h3):(1'h1)]);
              reg750 <= (((-reg700[(3'h4):(2'h2)]) ?
                  $unsigned((reg208[(2'h2):(1'h1)] <= $signed(reg227))) : $signed(({reg232} ?
                      ((8'haf) >>> reg671) : (8'ha4)))) == $signed(reg613));
              reg751 = ((~^$unsigned({$signed(reg468),
                  {(7'h43)},
                  reg696[(2'h2):(1'h0)]})) && (~&(((wire717 << reg649) || $signed(reg491)) ?
                  (((8'h9d) << reg700) ^~ (reg386 ?
                      (8'h9e) : reg228)) : reg276)));
              reg752 = {(|$unsigned(reg490[(2'h2):(1'h1)])),
                  reg300,
                  (reg430[(5'h11):(5'h10)] ?
                      $unsigned({$unsigned(reg616),
                          reg249}) : (!$unsigned($signed(forvar740))))};
              reg753 = $unsigned(reg592);
            end
        end
    end
  assign wire754 = reg438[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg755 = (!(~(reg744 | ((reg634 >> reg403) & (~&reg659)))));
      for (forvar756 = (1'h0); (forvar756 < (2'h3)); forvar756 = (forvar756 + (1'h1)))
        begin
          reg757 <= (^($unsigned((-{(8'hac), reg597, reg359})) <<< (7'h4e)));
          reg758 = $unsigned((reg472[(3'h4):(1'h0)] >> $signed(reg402[(4'he):(4'he)])));
        end
      for (forvar759 = (1'h0); (forvar759 < (1'h1)); forvar759 = (forvar759 + (1'h1)))
        begin
          reg760 <= $signed(reg707[(1'h0):(1'h0)]);
          for (forvar761 = (1'h0); (forvar761 < (1'h0)); forvar761 = (forvar761 + (1'h1)))
            begin
              reg762 <= $signed((reg602[(4'ha):(2'h2)] ?
                  (~^((|(7'h58)) ?
                      $signed((8'hb9)) : {reg338})) : $signed(($unsigned(reg602) | (reg316 ?
                      reg689 : (8'ha2))))));
            end
          reg763 <= ((reg259 ?
                  $unsigned(reg731[(4'h8):(4'h8)]) : $signed($signed((8'h9f)))) ?
              $signed((|(reg199 & $signed(reg429)))) : {((reg509 ?
                          (^reg760) : $signed((7'h47))) ?
                      reg434[(5'h13):(4'h8)] : (+(~^wire194))),
                  (!((reg320 ? reg496 : reg730) ?
                      $signed(reg365) : reg713[(3'h7):(1'h0)])),
                  reg338[(2'h2):(1'h0)]});
          for (forvar764 = (1'h0); (forvar764 < (3'h5)); forvar764 = (forvar764 + (1'h1)))
            begin
              reg765 = ((($signed(reg312[(3'h4):(3'h4)]) ?
                      {$unsigned(reg259),
                          (reg321 ? reg636 : reg446),
                          $signed(reg726)} : $signed(reg620[(3'h6):(3'h6)])) >> (|(reg610[(4'hd):(2'h2)] | reg393))) ?
                  reg727 : ($signed($unsigned(((7'h4e) ? reg359 : wire190))) ?
                      {(reg652 ?
                              {reg734,
                                  wire192} : $signed(reg515))} : (reg256[(3'h5):(3'h5)] ?
                          ((~&reg616) ?
                              (reg389 ?
                                  forvar759 : reg210) : $signed(reg338)) : $signed($signed((8'ha5))))));
            end
          for (forvar766 = (1'h0); (forvar766 < (2'h2)); forvar766 = (forvar766 + (1'h1)))
            begin
              reg767 <= (~{$unsigned(reg273[(4'hd):(3'h6)]),
                  $unsigned($unsigned({reg470}))});
            end
          for (forvar768 = (1'h0); (forvar768 < (3'h4)); forvar768 = (forvar768 + (1'h1)))
            begin
              reg769 <= reg231[(3'h7):(2'h2)];
              reg770 = $unsigned({$signed(($signed(reg258) ?
                      (reg227 != (8'hb6)) : reg474)),
                  ((^~reg243) ?
                      (reg339 < reg245) : ((!reg675) ?
                          $signed(reg339) : (|reg313)))});
              reg771 = $signed($unsigned(reg639));
            end
        end
      if ($unsigned(reg227[(4'ha):(3'h4)]))
        begin
          if (reg299)
            begin
              reg772 = ((|reg638[(3'h4):(1'h0)]) ?
                  {(($unsigned(reg674) ? $signed(reg693) : (8'hbe)) ?
                          reg493[(5'h16):(4'he)] : $signed((reg704 <= reg435))),
                      (reg341[(3'h6):(3'h6)] ?
                          (^reg667) : {reg655})} : reg699[(1'h0):(1'h0)]);
              reg773 <= $unsigned(($signed($unsigned({reg302})) ?
                  (+{$signed((8'hbd)), (reg403 ? reg770 : reg704)}) : reg610));
              reg774 <= reg284;
              reg775 <= reg762[(3'h7):(2'h3)];
              reg776 <= $unsigned(reg339[(4'h8):(3'h7)]);
            end
          else
            begin
              reg772 = ((((~&$signed(reg371)) ^~ reg664[(5'h15):(5'h14)]) ?
                      reg273 : reg511[(5'h16):(5'h11)]) ?
                  (~|$unsigned(reg338[(1'h0):(1'h0)])) : reg745);
              reg773 <= (((!reg421[(3'h6):(2'h2)]) ?
                      ((-$signed((7'h4e))) ?
                          $signed($signed((7'h44))) : reg724) : ((&$unsigned(reg667)) ?
                          (+$signed(reg460)) : (^~$signed(reg388)))) ?
                  (8'hb3) : $signed(((^(reg468 ? reg236 : reg589)) ?
                      $unsigned($unsigned(reg430)) : (7'h4e))));
            end
          if ($signed($unsigned(($unsigned({reg245,
              reg398,
              reg203}) | ((!reg203) ? (&reg398) : reg365)))))
            begin
              reg777 = $unsigned((+$unsigned(((reg370 - reg772) > $unsigned(reg627)))));
            end
          else
            begin
              reg778 <= $unsigned((reg480[(4'he):(3'h7)] || {({reg474,
                      wire754,
                      reg705} >> (reg734 ? reg505 : reg256))}));
              reg779 <= $signed({$unsigned({$unsigned((7'h43)), reg343}),
                  (~&reg330[(1'h0):(1'h0)])});
              reg780 = {(reg263 ? reg320 : (^reg273))};
              reg781 <= reg727[(3'h7):(3'h7)];
              reg782 <= reg238[(1'h1):(1'h1)];
              reg783 <= reg613[(4'hd):(1'h1)];
              reg784 = ($unsigned(((7'h4c) == forvar759)) > ((-((reg483 ?
                      reg659 : reg414) && {(8'h9d)})) ?
                  reg587[(5'h11):(4'he)] : reg514[(4'h8):(2'h3)]));
            end
          reg785 <= reg430;
          if (reg726)
            begin
              reg786 = wire584[(1'h0):(1'h0)];
              reg787 <= $signed(((|($signed(reg709) ?
                      $unsigned(reg675) : reg480[(4'he):(2'h2)])) ?
                  $signed(((reg434 >= reg494) ?
                      (reg403 > reg639) : ((8'hba) && reg627))) : (~&$unsigned((reg238 >> reg236)))));
              reg788 = $unsigned((~&{(^reg513)}));
              reg789 <= (^~reg414);
              reg790 <= ($signed(reg203) ?
                  (+($unsigned((reg742 ?
                      reg699 : (8'ha8))) || (!(-reg713)))) : reg683);
            end
          else
            begin
              reg787 <= (8'ha5);
              reg789 <= reg415;
              reg791 = reg652;
              reg792 = ({{{$unsigned((8'ha3)), $unsigned(reg507)}},
                      $unsigned($unsigned(((8'hb2) ? reg787 : (7'h52))))} ?
                  reg779[(5'h14):(5'h10)] : ((7'h43) ?
                      (reg453[(4'hb):(3'h4)] ^ (reg237[(2'h3):(1'h0)] ^ {reg709,
                          reg276})) : (~&((&wire192) >>> reg683[(2'h2):(2'h2)]))));
              reg793 <= (reg338 >> $unsigned((reg742[(2'h2):(1'h0)] ?
                  $unsigned(reg208) : $signed((reg252 <= reg612)))));
              reg794 = reg667;
              reg795 <= $unsigned(((8'hae) >>> (reg793[(3'h7):(2'h2)] >= reg243[(3'h6):(1'h1)])));
            end
          reg796 <= reg693[(4'hf):(4'hd)];
          reg797 = $unsigned((7'h57));
          if ($signed((((^~{reg776}) ?
                  (~^(reg468 ? reg484 : (8'h9c))) : (wire192 >> reg383)) ?
              $unsigned(reg284[(1'h0):(1'h0)]) : ({reg760,
                  (&reg398),
                  reg512} >> {reg440, $signed(reg388)}))))
            begin
              reg798 <= {reg501[(4'hb):(3'h7)],
                  {$signed($unsigned(reg389[(2'h3):(2'h2)]))}};
              reg799 = {(~(reg429[(3'h6):(3'h4)] != reg268[(3'h5):(1'h1)]))};
              reg800 = reg318;
            end
          else
            begin
              reg798 <= $unsigned(({reg502[(4'hf):(4'hf)],
                  (reg376[(4'hc):(1'h1)] ? (-reg635) : (reg434 && reg393)),
                  (reg468 ^ (reg225 != reg770))} ^ reg654[(2'h3):(1'h1)]));
              reg799 = $signed($unsigned(($signed((^~reg726)) | {$signed(reg201)})));
              reg800 = $unsigned(reg779[(4'he):(3'h5)]);
            end
        end
      else
        begin
          for (forvar772 = (1'h0); (forvar772 < (1'h0)); forvar772 = (forvar772 + (1'h1)))
            begin
              reg777 = (-reg345);
            end
          for (forvar778 = (1'h0); (forvar778 < (3'h6)); forvar778 = (forvar778 + (1'h1)))
            begin
              reg779 <= $unsigned(($signed(reg683) ?
                  wire190[(2'h3):(1'h1)] : reg657[(5'h16):(5'h11)]));
              reg780 = {(8'hb8),
                  reg424[(3'h5):(1'h1)],
                  (reg312 <= (!(-{reg424, reg648})))};
              reg784 = ($signed($signed(reg360)) > reg243);
              reg786 = {wire190, $signed(reg745)};
              reg787 <= $unsigned($signed(reg208));
              reg789 <= (({((reg755 ?
                              (8'ha3) : reg798) - forvar761[(1'h1):(1'h1)]),
                          $unsigned((|reg779))} ?
                      reg635 : (reg319[(1'h0):(1'h0)] ?
                          (^~$signed(reg797)) : (wire193[(4'hb):(1'h0)] ?
                              reg511[(4'ha):(1'h0)] : (~^reg634)))) ?
                  (((~|(!reg318)) ?
                      ({reg415} ?
                          reg243[(4'hc):(3'h6)] : $signed(reg772)) : $unsigned((reg293 || reg365))) >>> (($signed(reg373) > $signed(reg652)) != reg199[(5'h14):(4'h9)])) : reg667[(1'h0):(1'h0)]);
            end
          reg790 <= reg776;
          if ($signed((+$unsigned($unsigned(reg231)))))
            begin
              reg793 <= ((((~|(reg671 <<< reg312)) ?
                  (reg231 ^~ reg284) : $signed(((8'ha2) ?
                      reg774 : reg415))) | reg403[(5'h16):(4'he)]) ~^ ((~(~reg654[(2'h3):(2'h2)])) * $signed(((reg515 - (7'h56)) || $signed(reg293)))));
              reg794 = reg678[(1'h1):(1'h0)];
              reg797 = (((&(8'hb5)) < $unsigned($unsigned(reg324))) << {$signed(($unsigned(reg730) == reg663[(1'h1):(1'h0)]))});
              reg798 <= $signed(reg366[(2'h3):(2'h3)]);
              reg799 = (|$signed(reg345[(4'h8):(3'h7)]));
              reg801 <= (^((reg470[(4'hd):(4'h9)] > $signed(((7'h4d) ?
                  reg783 : reg471))) - reg244[(5'h14):(4'hc)]));
            end
          else
            begin
              reg791 = $signed(reg783);
              reg793 <= (^reg703);
              reg795 <= reg781[(2'h3):(2'h2)];
              reg797 = (reg707 | $signed($signed(($unsigned(reg338) ?
                  reg324 : $unsigned(reg421)))));
              reg799 = reg312;
              reg800 = reg606[(2'h3):(1'h1)];
              reg802 = (reg617 ~^ (~&(reg646 ?
                  {$unsigned(reg612),
                      reg371,
                      reg610[(4'hf):(1'h1)]} : $unsigned(wire350))));
            end
          if ((7'h50))
            begin
              reg803 <= $signed(((^~reg446[(3'h6):(3'h5)]) ?
                  (7'h55) : (8'hac)));
              reg804 = ({($signed($unsigned(reg653)) ?
                          (|reg456[(3'h5):(1'h1)]) : reg591)} ?
                  $unsigned($signed(forvar764)) : {$signed(($signed(reg727) ?
                          (7'h4f) : $unsigned(reg589))),
                      (~(&reg403)),
                      (&reg509)});
              reg805 <= (reg501[(3'h7):(3'h7)] ?
                  (reg456 ?
                      ($signed($signed(reg776)) >= reg627[(3'h7):(3'h7)]) : $unsigned(($unsigned(reg258) + reg236))) : $unsigned(reg249));
              reg806 = reg514[(4'hf):(3'h4)];
              reg807 = reg765[(1'h1):(1'h0)];
            end
          else
            begin
              reg803 <= (reg208 ? reg663 : {wire351[(5'h13):(5'h12)]});
              reg805 <= $unsigned($unsigned($unsigned(((reg657 ~^ reg781) << {reg512,
                  (7'h4a)}))));
              reg808 <= $unsigned((~^(reg744 < (((7'h4f) - reg218) <= $unsigned((8'h9c))))));
              reg809 <= (($signed($signed(reg434)) <= reg804) | $unsigned(wire754));
              reg810 <= reg806[(4'h9):(3'h5)];
            end
        end
      if ($signed($unsigned($signed(reg741))))
        begin
          if (reg613[(1'h1):(1'h1)])
            begin
              reg811 <= (reg373[(4'hc):(3'h4)] != ($signed($unsigned($signed(reg265))) ?
                  $signed((&(^reg797))) : reg430[(3'h7):(3'h4)]));
              reg812 = $unsigned(reg742);
            end
          else
            begin
              reg812 = (^~$signed(reg702));
              reg813 <= (~|reg245[(5'h10):(1'h1)]);
            end
          for (forvar814 = (1'h0); (forvar814 < (1'h0)); forvar814 = (forvar814 + (1'h1)))
            begin
              reg815 <= $unsigned(((+$unsigned(reg728[(4'hb):(2'h3)])) + reg287[(4'hc):(2'h3)]));
              reg816 = $unsigned($signed($unsigned((~^{forvar761, reg724}))));
              reg817 = reg269;
            end
          for (forvar818 = (1'h0); (forvar818 < (2'h3)); forvar818 = (forvar818 + (1'h1)))
            begin
              reg819 = reg236[(3'h4):(3'h4)];
              reg820 = reg318[(2'h3):(2'h2)];
            end
          if ({$signed(((~|$signed(reg780)) != reg607)),
              (~&$unsigned((reg819[(2'h3):(1'h1)] ^~ $unsigned(reg231)))),
              $unsigned(reg770)})
            begin
              reg821 = reg688;
              reg822 = $signed({reg728, reg593, (!reg456[(4'hf):(4'he)])});
              reg823 = $unsigned((!$unsigned(($signed((8'hae)) ?
                  $unsigned(wire351) : (^~reg370)))));
              reg824 = reg727;
              reg825 = ($unsigned((($signed(forvar814) == (reg284 ?
                      reg493 : reg624)) ?
                  reg230[(4'h8):(1'h1)] : $signed(reg446))) ~^ reg793[(2'h2):(1'h0)]);
              reg826 = reg216[(4'hc):(4'h8)];
              reg827 <= {(($unsigned($signed(reg813)) <= $unsigned(reg365[(1'h1):(1'h0)])) ^ (((wire190 ?
                          reg773 : (8'ha1)) ^~ (&reg815)) ?
                      $unsigned($unsigned(reg589)) : (&(8'hb1))))};
            end
          else
            begin
              reg821 = reg215;
              reg822 = {$signed($unsigned((-(wire193 ~^ reg696)))),
                  (~^$unsigned(((^~reg817) ^ $signed(reg591))))};
              reg827 <= $unsigned(reg362);
            end
          if (reg373)
            begin
              reg828 <= (reg778 * reg606);
            end
          else
            begin
              reg828 <= (forvar772[(5'h11):(4'hf)] ?
                  (~(((|reg809) ? $unsigned(reg341) : (7'h48)) ?
                      $unsigned((^~reg511)) : ($unsigned(reg243) || reg445[(4'he):(3'h7)]))) : {{(reg635[(1'h0):(1'h0)] ?
                              $signed(reg480) : (reg788 * reg501)),
                          $unsigned((8'hb5))},
                      ((&$signed(reg231)) ?
                          {$unsigned(reg819),
                              reg648[(3'h4):(2'h3)],
                              (reg763 | reg765)} : $unsigned((reg709 << reg507))),
                      $unsigned(($unsigned(reg826) + reg700[(3'h5):(2'h3)]))});
              reg829 = (^~(^~({{reg210}, $unsigned(reg616), (!reg365)} ?
                  reg789[(5'h1a):(5'h13)] : ({reg364, wire717} ?
                      (~^reg649) : reg483[(4'hf):(4'he)]))));
              reg830 = $unsigned(($unsigned(({reg646,
                  (8'hbd),
                  reg365} > $unsigned(reg269))) || reg258));
              reg831 = $unsigned($unsigned($signed((7'h45))));
              reg832 <= $unsigned(reg263);
              reg833 <= $unsigned($unsigned((reg786 || $signed((reg789 ?
                  (8'hac) : (8'haa))))));
              reg834 <= ((reg231[(4'hb):(1'h0)] ?
                  ((~reg341[(4'h9):(3'h7)]) ?
                      $signed((7'h4d)) : ($unsigned(reg597) ^ reg283[(3'h4):(2'h3)])) : $unsigned((~(reg822 ?
                      reg709 : reg376)))) + ($unsigned($unsigned(reg302)) ?
                  reg652[(4'ha):(3'h4)] : ($signed((reg237 ?
                      reg793 : reg809)) >> ($signed(reg828) ?
                      (|reg635) : $signed(forvar761)))));
            end
        end
      else
        begin
          for (forvar811 = (1'h0); (forvar811 < (3'h6)); forvar811 = (forvar811 + (1'h1)))
            begin
              reg812 = (reg312[(3'h5):(3'h5)] + $unsigned(reg300));
              reg814 = reg324;
              reg816 = (reg826 >> ((+$signed($unsigned(reg218))) - reg804[(3'h4):(1'h1)]));
              reg818 <= reg232;
              reg819 = $unsigned($unsigned((8'hbf)));
              reg820 = reg273[(5'h15):(2'h3)];
              reg827 <= $signed($unsigned($unsigned(reg708)));
            end
          reg828 <= $unsigned(($signed((+$signed((7'h4d)))) && reg825[(3'h5):(2'h2)]));
          for (forvar829 = (1'h0); (forvar829 < (3'h4)); forvar829 = (forvar829 + (1'h1)))
            begin
              reg832 <= $signed($unsigned((((|reg265) ?
                      $unsigned((8'hb1)) : {reg415, reg444, reg813}) ?
                  reg199[(3'h5):(2'h3)] : reg750)));
              reg835 = ($signed(reg318) > ($unsigned(reg414) ?
                  $signed((reg430[(5'h14):(4'hf)] ^ ((7'h54) > reg484))) : ($unsigned({reg829,
                          reg376}) ?
                      (reg208[(1'h1):(1'h1)] >= reg339) : wire192)));
              reg836 = (~reg252);
              reg837 <= {{$signed((!(reg362 ? reg444 : reg728))),
                      (reg255[(3'h4):(2'h3)] ^ reg675[(3'h5):(2'h2)]),
                      reg757[(4'hc):(1'h0)]}};
              reg838 = $signed(reg678);
            end
        end
      reg839 <= forvar814[(3'h4):(2'h2)];
    end
  always
    @(posedge clk) begin
      if (reg747)
        begin
          if (reg650[(5'h14):(4'hf)])
            begin
              reg840 = ($signed(({(&(8'haf)), reg833[(5'h14):(4'hb)]} ?
                  reg655[(1'h0):(1'h0)] : $signed($signed(reg620)))) ^~ reg839);
              reg841 <= $unsigned($signed(reg205));
              reg842 <= {(~|reg650), reg727};
              reg843 = ((((7'h4d) > $signed($signed(wire351))) ?
                      $unsigned((reg511[(5'h10):(4'hb)] ?
                          (reg834 ?
                              reg339 : (7'h55)) : $signed(reg362))) : $signed(wire194[(5'h17):(5'h16)])) ?
                  {$signed(((reg364 | reg592) ?
                          $signed(reg655) : (reg386 && reg787))),
                      $unsigned(reg703[(3'h4):(2'h2)]),
                      (8'hae)} : ({(~|reg776[(3'h6):(2'h3)])} <= $unsigned($unsigned(reg705))));
              reg844 <= reg258;
              reg845 = (({reg724[(4'hd):(3'h7)]} ?
                  (((reg429 ^~ (8'hb5)) ^~ reg511) ?
                      (~|(~^reg445)) : ($unsigned(reg698) - (reg243 ^ reg302))) : reg813) != $signed((!reg474)));
              reg846 <= (^~reg741[(5'h11):(4'ha)]);
            end
          else
            begin
              reg840 = (&reg839[(2'h2):(2'h2)]);
              reg843 = reg270[(4'ha):(1'h1)];
            end
          for (forvar847 = (1'h0); (forvar847 < (2'h3)); forvar847 = (forvar847 + (1'h1)))
            begin
              reg848 = ($unsigned(($signed((reg335 ?
                      (7'h58) : reg345)) >= {((8'hb2) * reg339)})) ?
                  ((+$signed((~reg502))) ?
                      (~^$signed(reg440)) : (reg402 <<< $signed($signed(reg744)))) : ($unsigned($unsigned($signed(reg696))) ?
                      reg287 : (({reg762} ? reg474 : reg774) || reg199)));
              reg849 <= (~|reg655[(1'h0):(1'h0)]);
              reg850 <= ((reg769[(3'h4):(2'h2)] ?
                      $signed($signed((+reg430))) : (((wire516 >= reg654) ?
                          (reg438 * reg429) : $unsigned((7'h52))) ~^ reg597)) ?
                  $unsigned($unsigned($signed((reg793 ?
                      reg789 : reg769)))) : (reg259 ?
                      (reg245 ?
                          (wire195 ?
                              (reg283 ?
                                  reg338 : reg648) : $signed(reg671)) : (~^$unsigned(reg641))) : $signed($unsigned((~reg688)))));
              reg851 = (reg359[(1'h0):(1'h0)] ^~ $unsigned((reg471[(2'h3):(2'h3)] ?
                  (8'h9f) : ($signed(reg774) ?
                      (reg796 && reg653) : $unsigned((8'hb3))))));
            end
          reg852 = $unsigned($unsigned({($signed(reg779) - reg810)}));
          reg853 <= (reg505[(2'h2):(2'h2)] + $unsigned((wire754 ?
              (~|$signed(wire351)) : ((8'haa) ^~ (reg283 || reg785)))));
        end
      else
        begin
          reg841 <= reg321[(4'hc):(4'h8)];
          for (forvar842 = (1'h0); (forvar842 < (1'h0)); forvar842 = (forvar842 + (1'h1)))
            begin
              reg843 = $unsigned((^reg674));
              reg844 <= $signed(reg339);
              reg845 = $unsigned($signed(reg673[(2'h2):(1'h1)]));
            end
          if ($unsigned((7'h54)))
            begin
              reg846 <= reg232[(1'h1):(1'h0)];
              reg847 <= $signed((|($unsigned((~^reg424)) | reg709)));
              reg848 = ((+(~&reg648)) ?
                  (($signed(reg255[(3'h6):(2'h2)]) ?
                      reg818[(5'h1f):(5'h1e)] : (^(8'h9d))) >> (8'ha3)) : reg700[(3'h4):(3'h4)]);
              reg849 <= reg501;
            end
          else
            begin
              reg846 <= (|$unsigned(reg843[(4'h9):(3'h6)]));
              reg848 = reg346;
              reg849 <= reg848;
            end
        end
      reg854 = (~&reg360);
      for (forvar855 = (1'h0); (forvar855 < (3'h4)); forvar855 = (forvar855 + (1'h1)))
        begin
          if (reg435)
            begin
              reg856 <= reg793;
              reg857 = ($unsigned(wire717[(2'h2):(1'h0)]) ?
                  reg414[(1'h1):(1'h0)] : (reg704[(3'h5):(1'h0)] ?
                      {reg657[(4'hd):(3'h5)]} : (!(reg276 ?
                          (-reg627) : forvar842[(4'h9):(3'h6)]))));
              reg858 <= reg319[(2'h2):(1'h1)];
              reg859 <= (reg837[(1'h0):(1'h0)] ?
                  (&$signed($signed((reg470 ?
                      reg471 : reg470)))) : ($signed($unsigned($signed((8'hab)))) ?
                      reg844[(1'h1):(1'h1)] : $unsigned($signed($unsigned(reg699)))));
              reg860 = (~&$signed($unsigned(($unsigned(reg503) ?
                  reg316 : $signed((7'h41))))));
            end
          else
            begin
              reg856 <= reg639[(3'h5):(3'h5)];
              reg857 = (reg813 ~^ {reg341[(4'h9):(2'h2)],
                  $signed(($signed(reg403) ? (reg627 - reg704) : (^reg218)))});
              reg860 = {((({(7'h4c)} ? reg818 : reg276) << (reg616 ?
                      (reg648 ?
                          reg244 : reg775) : (~|reg421))) && $signed({$unsigned(reg218),
                      $unsigned(reg592)})),
                  $unsigned((8'hb2)),
                  reg828[(4'h9):(3'h7)]};
              reg861 = (~(reg230 ?
                  (~({(7'h4a), reg512, reg265} << (&reg760))) : (^reg750)));
            end
          reg862 = (wire717 << $unsigned((~&((8'hb6) >= (reg776 ?
              (7'h4e) : reg674)))));
          if ((reg808[(4'h8):(2'h3)] <<< $unsigned((&(-(&reg861))))))
            begin
              reg863 <= $unsigned((reg502 ^ reg736[(1'h0):(1'h0)]));
              reg864 <= (+reg650[(3'h5):(1'h1)]);
              reg865 = (^(^reg462));
              reg866 <= ($signed($signed($signed({reg474, reg256, reg843}))) ?
                  $unsigned({((8'ha2) ?
                          (reg435 ? reg483 : reg302) : $unsigned(reg773)),
                      (reg750 * (reg675 || (7'h40))),
                      ((~&reg678) ?
                          reg592[(1'h1):(1'h1)] : (~|reg619))}) : (((~^$unsigned(reg741)) ^ (reg494[(2'h2):(1'h1)] ?
                      forvar855[(5'h1b):(4'h8)] : reg587)) >> reg645[(2'h3):(2'h3)]));
              reg867 = (^~$unsigned($signed((!reg850))));
              reg868 = reg396;
            end
          else
            begin
              reg865 = $signed({($unsigned((~|reg273)) >= $unsigned((reg366 ?
                      reg760 : reg283))),
                  (($unsigned(reg709) ?
                      (forvar842 ?
                          forvar842 : reg678) : (reg338 <<< (8'hb3))) - {(reg842 ?
                          reg319 : reg509),
                      {reg619, reg664, reg600}}),
                  reg365[(4'h8):(3'h5)]});
              reg866 <= (|$signed($signed(($unsigned(reg730) | $signed(reg844)))));
              reg867 = reg851;
            end
          for (forvar869 = (1'h0); (forvar869 < (2'h2)); forvar869 = (forvar869 + (1'h1)))
            begin
              reg870 <= {(reg256 ?
                      $signed(($unsigned(reg509) ?
                          (reg775 < (7'h46)) : (~|reg293))) : $unsigned(($unsigned(reg724) ?
                          reg396[(3'h7):(3'h7)] : (^reg416)))),
                  reg767[(1'h0):(1'h0)],
                  $unsigned(reg843)};
              reg871 <= (reg446 >= $unsigned(reg480[(3'h5):(3'h5)]));
              reg872 <= $signed((7'h40));
              reg873 = $unsigned($signed(((8'hb2) ?
                  (~^$signed(reg238)) : reg674[(1'h0):(1'h0)])));
              reg874 <= (8'hb3);
              reg875 = reg818;
            end
          for (forvar876 = (1'h0); (forvar876 < (3'h4)); forvar876 = (forvar876 + (1'h1)))
            begin
              reg877 = reg335[(1'h1):(1'h0)];
              reg878 <= reg689;
              reg879 <= reg210;
              reg880 <= (reg373[(4'ha):(1'h1)] > reg462);
              reg881 <= $unsigned(($unsigned(reg341[(3'h6):(2'h3)]) ?
                  (~&$unsigned(((8'ha7) <<< (7'h57)))) : $unsigned(($signed(reg227) ^~ {reg763,
                      reg655,
                      reg663}))));
              reg882 = ($unsigned($unsigned(reg453)) ^ (7'h4f));
              reg883 = (^reg434);
            end
        end
      reg884 <= reg653;
      reg885 = reg667;
      reg886 = reg648[(2'h3):(1'h0)];
      for (forvar887 = (1'h0); (forvar887 < (1'h1)); forvar887 = (forvar887 + (1'h1)))
        begin
          for (forvar888 = (1'h0); (forvar888 < (1'h1)); forvar888 = (forvar888 + (1'h1)))
            begin
              reg889 <= (reg745 >>> reg238[(2'h2):(1'h1)]);
              reg890 = (~&((reg645 ?
                      (((7'h55) * (8'hbb)) ?
                          reg837 : (reg512 ? reg655 : reg730)) : ((reg276 ?
                          reg255 : (8'ha6)) < (~^(8'hab)))) ?
                  (reg618[(1'h0):(1'h0)] ?
                      reg593 : (((7'h40) == reg742) ?
                          reg878 : (!reg346))) : (8'ha1)));
              reg891 <= reg307[(4'h8):(2'h3)];
              reg892 <= reg335;
              reg893 = (!reg683[(1'h1):(1'h1)]);
              reg894 = reg616;
              reg895 <= (8'h9d);
            end
        end
    end
  module896 #() modinst1495 (wire1494, clk, reg683, reg750, reg638, reg468);
  always
    @(posedge clk) begin
      for (forvar1496 = (1'h0); (forvar1496 < (3'h6)); forvar1496 = (forvar1496 + (1'h1)))
        begin
          reg1497 <= reg316;
          for (forvar1498 = (1'h0); (forvar1498 < (1'h1)); forvar1498 = (forvar1498 + (1'h1)))
            begin
              reg1499 = reg619;
              reg1500 <= $signed((~reg693[(5'h10):(1'h0)]));
              reg1501 <= ((reg199 & {($signed(reg299) ?
                          ((8'hbe) > (8'hbb)) : (~|reg783))}) ?
                  $unsigned(reg635) : ($unsigned(((^~reg256) ?
                          (reg808 ? (7'h51) : reg293) : $unsigned((7'h4d)))) ?
                      $signed($unsigned($signed((7'h40)))) : (^reg744[(3'h6):(1'h0)])));
              reg1502 = reg507;
            end
        end
      reg1503 = reg493[(5'h14):(4'h9)];
      if ((+reg492))
        begin
          for (forvar1504 = (1'h0); (forvar1504 < (1'h1)); forvar1504 = (forvar1504 + (1'h1)))
            begin
              reg1505 = reg364;
              reg1506 = (&$signed(reg853[(4'h8):(1'h0)]));
              reg1507 <= (8'hb3);
              reg1508 <= ($signed(((~&$signed(reg801)) * $unsigned({reg837,
                      reg624}))) ?
                  ($unsigned(reg745[(3'h6):(3'h4)]) ?
                      (7'h48) : ({reg244, (~reg232)} ^~ ($unsigned(wire1494) ?
                          (+reg636) : (^(8'hae))))) : $unsigned((reg604[(4'he):(1'h1)] & reg474)));
              reg1509 = (~^((~($unsigned(reg513) ?
                      (reg833 || (7'h4b)) : (7'h4a))) ?
                  (~&($unsigned(reg702) ~^ $unsigned(wire194))) : reg440));
              reg1510 = reg757[(4'h9):(4'h8)];
            end
          reg1511 = $signed(reg593[(4'hd):(3'h5)]);
          reg1512 = reg388[(3'h7):(2'h3)];
          reg1513 = ((reg726[(4'hd):(3'h4)] > ($signed($signed(reg388)) ?
              reg773 : reg472)) ^ reg468);
          for (forvar1514 = (1'h0); (forvar1514 < (1'h0)); forvar1514 = (forvar1514 + (1'h1)))
            begin
              reg1515 = (~&reg703);
              reg1516 <= (({reg268,
                  (reg795 ^ $signed((7'h51)))} <= $unsigned(reg483[(1'h0):(1'h0)])) ~^ (-(^(reg484[(2'h3):(2'h2)] <<< reg675[(1'h1):(1'h0)]))));
              reg1517 <= (8'hbe);
            end
        end
      else
        begin
          for (forvar1504 = (1'h0); (forvar1504 < (3'h4)); forvar1504 = (forvar1504 + (1'h1)))
            begin
              reg1507 <= reg330;
              reg1509 = $unsigned(((^~$unsigned((reg779 ?
                  reg672 : reg255))) ^ ((7'h44) < reg779)));
              reg1514 <= reg389;
              reg1516 <= reg683[(4'h9):(1'h0)];
              reg1517 <= $unsigned((reg424 == reg744));
              reg1518 = ((8'ha7) >= ({$unsigned({reg837, (8'ha7)}),
                  $signed($signed(reg259))} >> reg316));
              reg1519 = reg245[(4'hc):(3'h7)];
            end
          if ($unsigned({(+reg884),
              $signed((~(reg798 ? reg776 : reg616))),
              reg472}))
            begin
              reg1520 = $signed((~|reg460[(3'h4):(1'h0)]));
            end
          else
            begin
              reg1520 = reg1501[(5'h1d):(5'h16)];
              reg1521 = ($signed({reg471}) > $signed(reg593));
              reg1522 = reg237[(3'h5):(2'h3)];
            end
          if (reg809[(4'he):(1'h0)])
            begin
              reg1523 <= (reg370[(5'h12):(4'he)] - (reg494[(5'h1f):(1'h0)] ^ ($unsigned($unsigned(reg502)) <= (~reg664))));
            end
          else
            begin
              reg1523 <= (reg610 ~^ $unsigned((((~&reg853) >>> (~|reg244)) * $unsigned((~|reg787)))));
              reg1524 <= ((($signed($unsigned(reg1508)) != (~$signed(reg891))) && reg727) & (reg856 || (8'ha6)));
              reg1525 <= reg434[(5'h19):(4'he)];
            end
          for (forvar1526 = (1'h0); (forvar1526 < (2'h3)); forvar1526 = (forvar1526 + (1'h1)))
            begin
              reg1527 <= ($signed($signed((~&reg839))) >> (((|{reg331}) - (~|reg474[(5'h15):(4'hb)])) * $unsigned(reg849[(4'hb):(2'h2)])));
              reg1528 <= reg607;
              reg1529 <= $signed(reg393[(4'hd):(4'hc)]);
              reg1530 = ($signed((~|($signed(reg1500) >> (reg483 ?
                  (8'ha5) : reg1506)))) <<< $unsigned((|(+$unsigned(reg429)))));
              reg1531 = ($unsigned(((!$signed(reg602)) ?
                  ((reg815 ? reg365 : reg228) ?
                      {reg879, reg416} : reg225) : (reg757 ?
                      reg610 : $unsigned((7'h55))))) | $unsigned(($unsigned(reg346) ?
                  {reg704[(4'ha):(2'h3)]} : $signed($signed(reg849)))));
              reg1532 <= $unsigned($unsigned({reg619[(4'h9):(4'h9)]}));
            end
        end
      if (reg276[(3'h4):(2'h2)])
        begin
          reg1533 <= ((|$signed((8'hae))) ?
              $unsigned((($unsigned(reg762) ?
                      $signed(reg359) : (reg435 << reg490)) ?
                  ((8'h9c) ?
                      $signed(reg364) : (^~reg1513)) : (!$unsigned(wire193)))) : ($signed((8'hb2)) ^~ (+reg511[(4'hb):(3'h7)])));
          reg1534 <= ({reg808[(3'h4):(3'h4)], (&reg203)} ?
              {(reg460 ? reg514[(5'h18):(3'h5)] : $unsigned((+reg507))),
                  $signed($unsigned((reg389 | reg263)))} : (8'hbf));
          reg1535 = {((^~{reg672,
                      (wire516 ? reg704 : reg648),
                      {reg1523, reg345}}) ?
                  ({forvar1504[(4'hb):(1'h1)]} ?
                      ((reg850 ~^ reg834) + $signed(forvar1498)) : reg238[(2'h2):(2'h2)]) : reg785),
              ($unsigned((-reg783[(4'hf):(3'h4)])) ?
                  ((-(^reg809)) ?
                      (~^(-reg1525)) : (8'ha5)) : $unsigned($signed($signed(reg731)))),
              (reg399[(1'h0):(1'h0)] <= (+(8'hbb)))};
        end
      else
        begin
          reg1535 = ((reg782 || $unsigned(($signed(reg773) >= reg364[(2'h3):(1'h0)]))) ?
              (8'haa) : {reg728,
                  $unsigned((reg734[(5'h15):(2'h3)] >= $unsigned(reg343)))});
        end
      for (forvar1536 = (1'h0); (forvar1536 < (2'h3)); forvar1536 = (forvar1536 + (1'h1)))
        begin
          if (reg345)
            begin
              reg1537 <= $unsigned($unsigned(wire193));
            end
          else
            begin
              reg1538 = reg268;
              reg1539 <= (($unsigned((~^(|reg232))) ?
                      $unsigned(({wire193, reg1532, reg1505} ?
                          (forvar1504 ?
                              reg324 : reg813) : reg597[(1'h0):(1'h0)])) : ($unsigned($signed(reg414)) * (~^(reg703 ?
                          reg745 : reg1499)))) ?
                  reg859 : $unsigned((reg373 <= $unsigned((wire193 <<< (8'hb2))))));
              reg1540 = {$unsigned($unsigned({$unsigned(reg613),
                      $signed(reg655),
                      reg365}))};
              reg1541 = {$unsigned((reg880 >>> reg258))};
            end
          for (forvar1542 = (1'h0); (forvar1542 < (2'h3)); forvar1542 = (forvar1542 + (1'h1)))
            begin
              reg1543 = (~&$signed((+(!$unsigned(reg338)))));
              reg1544 <= $signed(reg362);
            end
          reg1545 = reg490[(2'h2):(2'h2)];
          reg1546 = $signed({reg273[(3'h7):(2'h2)], wire754[(3'h4):(2'h2)]});
          if (($signed((reg307[(4'hf):(1'h0)] ^~ reg300[(2'h3):(1'h1)])) ~^ ({(8'hbd),
              ((reg757 ? (7'h55) : reg702) ?
                  reg657[(5'h11):(4'hb)] : (reg371 > reg255)),
              ($unsigned(reg388) ?
                  $signed(reg591) : (|reg832))} & (reg774[(5'h12):(3'h6)] ^ reg760))))
            begin
              reg1547 = (($signed(((reg769 ? reg762 : reg673) & {reg671,
                      (7'h56),
                      reg1508})) || (($signed(reg776) ?
                          (|reg699) : (reg300 != reg613)) ?
                      $unsigned((|(8'hbd))) : (reg801[(3'h6):(3'h5)] ^~ (reg512 < reg1522)))) ?
                  ((((8'ha9) <<< (^~(7'h45))) ?
                          ((~|reg762) & $signed((8'had))) : reg475) ?
                      reg360[(3'h7):(1'h1)] : $unsigned({reg273[(2'h3):(2'h2)],
                          (reg778 ? reg892 : reg307),
                          reg453[(4'hd):(4'ha)]})) : $signed(reg655[(2'h2):(1'h1)]));
              reg1548 <= ({reg227[(4'h8):(3'h6)],
                      ($unsigned(reg414[(1'h0):(1'h0)]) > reg1519[(1'h1):(1'h0)])} ?
                  reg664[(4'hb):(3'h5)] : $signed((&reg1546[(5'h17):(4'h9)])));
              reg1549 <= {$unsigned((~^{(reg1517 ? reg856 : (7'h49)),
                      $signed(forvar1504)})),
                  ((~&$unsigned(((8'ha4) ?
                      reg726 : reg1509))) || ($unsigned($unsigned(reg828)) ?
                      ((~reg330) ^ (~^wire718)) : $signed(reg874))),
                  reg245[(2'h3):(2'h2)]};
              reg1550 <= wire191[(4'hb):(2'h2)];
              reg1551 <= (reg815[(5'h13):(4'hf)] >>> (~^$signed(reg371[(4'ha):(3'h6)])));
              reg1552 <= {reg607[(4'hc):(3'h7)],
                  (((^reg1545[(3'h6):(3'h6)]) ?
                      ((~^(8'hb2)) ?
                          (~reg592) : (7'h47)) : (+$signed(wire717))) != ({(!(7'h58))} >>> reg256[(2'h3):(1'h0)]))};
            end
          else
            begin
              reg1548 <= $unsigned($signed((+$signed(reg438[(2'h3):(1'h1)]))));
              reg1553 = reg789[(4'hb):(1'h0)];
              reg1554 <= reg782[(1'h1):(1'h0)];
            end
        end
      if ($signed(reg675[(4'h9):(3'h7)]))
        begin
          if (reg218[(4'hb):(3'h5)])
            begin
              reg1555 <= $unsigned(reg673[(1'h0):(1'h0)]);
              reg1556 = $signed(((((reg434 ^ wire191) ~^ $signed(reg1541)) && (&((8'hb5) * reg1547))) ^ forvar1504));
              reg1557 = $unsigned((reg318[(2'h3):(2'h3)] ?
                  $unsigned(reg511[(4'he):(4'hb)]) : reg258));
              reg1558 <= (reg844 ?
                  $signed(reg864) : ($signed(reg203) < (((8'hb1) <<< $signed(reg513)) ?
                      reg414 : ((8'ha3) >>> (reg327 ? reg813 : reg346)))));
              reg1559 <= ({$signed(reg778),
                      $unsigned((reg345 ?
                          (reg669 ? reg850 : reg832) : $signed((8'hbe))))} ?
                  $signed($unsigned($signed((reg468 ?
                      reg1529 : reg471)))) : ($signed(reg744[(2'h2):(2'h2)]) ?
                      {$unsigned(((8'ha6) ? reg231 : (7'h47))),
                          ((~|reg1557) ^ (forvar1514 ? (8'ha6) : reg810)),
                          $signed((reg663 << reg278))} : reg513));
              reg1560 <= forvar1498;
              reg1561 = {(reg265[(1'h1):(1'h1)] ?
                      $signed($unsigned(reg762[(4'hd):(4'hd)])) : reg895[(3'h5):(3'h5)]),
                  reg604};
            end
          else
            begin
              reg1556 = reg785;
              reg1557 = (^~$signed((|reg879)));
              reg1558 <= (reg430 != reg1505[(2'h2):(2'h2)]);
              reg1559 <= ((reg636 ?
                      (((~|reg895) ? $signed((8'h9e)) : {reg345}) ?
                          reg398[(1'h0):(1'h0)] : $unsigned((7'h4c))) : (($signed(reg859) <<< (reg280 ~^ reg225)) ?
                          ($signed((8'ha2)) != (~|reg727)) : $signed({reg388,
                              reg208}))) ?
                  (reg1499[(2'h3):(2'h3)] ?
                      $signed($signed(reg1530[(3'h4):(2'h2)])) : $signed($signed(reg273[(4'hb):(4'hb)]))) : $signed((reg243 >> $unsigned($signed(reg1507)))));
              reg1561 = (reg727 + reg602);
              reg1562 <= (~reg343);
            end
          reg1563 <= ((&reg1497[(5'h13):(3'h5)]) ^~ (~(($unsigned(reg833) ?
                  {(8'ha3), reg300, (8'ha2)} : $signed(wire584)) ?
              $signed(reg511) : ($unsigned(reg1515) ?
                  reg490 : (reg891 == forvar1526)))));
          for (forvar1564 = (1'h0); (forvar1564 < (3'h6)); forvar1564 = (forvar1564 + (1'h1)))
            begin
              reg1565 = reg1512[(3'h4):(1'h0)];
              reg1566 <= reg648[(2'h3):(2'h2)];
              reg1567 = ((reg808 ?
                      (forvar1514 ^~ {(reg1534 ^ reg475)}) : (~&reg1517)) ?
                  $unsigned((reg1531 ?
                      $signed(((7'h49) ?
                          reg892 : reg471)) : (reg1528[(2'h2):(1'h0)] <<< reg507[(4'hb):(3'h7)]))) : $unsigned($unsigned((~|(&reg491)))));
            end
          reg1568 = $signed(((reg244 + reg435) ?
              reg502[(5'h13):(2'h3)] : reg880));
          for (forvar1569 = (1'h0); (forvar1569 < (2'h3)); forvar1569 = (forvar1569 + (1'h1)))
            begin
              reg1570 = reg1538;
              reg1571 <= $signed(reg853);
              reg1572 <= $signed((($unsigned(((7'h4c) ?
                      reg747 : reg700)) ^~ {reg1563[(4'h8):(2'h3)]}) ?
                  ({reg373[(4'he):(1'h0)],
                      (reg343 ? reg1499 : reg674),
                      $signed(reg430)} << ($unsigned(reg892) <<< reg809[(4'ha):(1'h1)])) : {(!$signed(reg1507))}));
              reg1573 = reg593;
              reg1574 = (~&reg1530[(3'h7):(2'h3)]);
            end
          reg1575 <= (^$signed(((^{reg635,
              (8'hbd)}) >> reg1555[(5'h12):(2'h3)])));
          if ((reg430 ~^ reg338))
            begin
              reg1576 <= {(reg745[(2'h2):(1'h0)] - (|$unsigned({reg815,
                      reg1522,
                      reg1512}))),
                  reg317};
              reg1577 <= {$signed(($signed((&reg707)) || ((reg639 ?
                          reg1505 : reg327) ?
                      (reg311 >= reg881) : (&reg674))))};
              reg1578 <= ({($signed((+(7'h4d))) << (+reg273)),
                      {{(reg447 < reg763), reg346[(2'h3):(1'h1)]},
                          reg440[(3'h4):(1'h0)],
                          (-$signed(forvar1536))}} ?
                  reg1576 : $signed($signed(($unsigned(reg511) & (!(8'hbe))))));
            end
          else
            begin
              reg1579 = (reg1550 ?
                  (~$signed(reg398[(3'h5):(3'h5)])) : $unsigned({($unsigned(reg1517) && (reg1530 ?
                          reg249 : reg270)),
                      $signed((~|reg698)),
                      $unsigned($signed(reg618))}));
              reg1580 <= (|(~|(~&(7'h51))));
            end
        end
      else
        begin
          reg1556 = reg1577;
          reg1557 = (reg210 ?
              {((reg199[(5'h1a):(4'ha)] ? $signed(reg255) : reg674) ?
                      reg1560[(3'h4):(2'h3)] : $signed({reg480,
                          reg444,
                          reg874})),
                  (reg1510 ^ (reg203[(4'h9):(1'h0)] ?
                      (reg616 >>> reg501) : (reg858 > reg591)))} : $signed((|(reg652[(5'h10):(4'hc)] ?
                  (reg1523 ? (8'hb2) : (8'h9e)) : reg318))));
        end
    end
  always
    @(posedge clk) begin
      reg1581 = ($signed(($signed($signed(reg810)) ?
              $unsigned($unsigned(reg278)) : ({(8'h9c)} ?
                  reg798[(3'h6):(2'h2)] : $unsigned(reg258)))) ?
          (((~^(reg503 || reg1555)) ?
                  $signed({reg652, reg871}) : $signed({reg230})) ?
              reg589 : reg280[(4'hc):(4'hb)]) : $signed(reg880));
      reg1582 = {({(~|((7'h40) << reg787))} && {reg892[(3'h5):(3'h4)],
              reg299})};
      reg1583 <= wire195[(3'h6):(2'h3)];
      reg1584 <= $unsigned(reg362[(4'ha):(4'ha)]);
      for (forvar1585 = (1'h0); (forvar1585 < (1'h0)); forvar1585 = (forvar1585 + (1'h1)))
        begin
          reg1586 <= $unsigned({($signed(reg232) ?
                  reg293 : $signed((reg811 >> reg785))),
              ($unsigned($unsigned((8'hb9))) >> (~&$unsigned(reg827)))});
          if ($signed((~^$signed(reg713[(3'h4):(3'h4)]))))
            begin
              reg1587 <= $unsigned($signed((-((reg312 & (7'h52)) <<< $unsigned(reg1578)))));
              reg1588 = reg496[(1'h1):(1'h0)];
              reg1589 <= ((~|(reg837 ?
                      {(|reg879), (8'h9e)} : (((7'h51) - reg474) ?
                          (^~reg231) : reg365))) ?
                  {$unsigned((-reg734[(5'h15):(4'ha)])),
                      reg318[(3'h5):(1'h0)]} : (&(reg1566 == (reg689 ?
                      reg365[(3'h5):(1'h1)] : $unsigned(reg386)))));
              reg1590 = ({{$signed($unsigned(reg300))},
                  $unsigned($unsigned(reg874))} || ({$unsigned((~&reg484))} ?
                  $unsigned(($unsigned(reg624) ?
                      reg810 : (~^(8'hbc)))) : reg1572));
              reg1591 <= reg832[(5'h1d):(3'h5)];
              reg1592 = ((!(reg619 ^ reg699)) || {$unsigned(reg434)});
              reg1593 = (~(!$unsigned(($signed(reg646) ?
                  (reg273 != (7'h52)) : (~&reg648)))));
            end
          else
            begin
              reg1588 = $unsigned($signed($unsigned(((reg364 + reg1550) ?
                  $signed(reg796) : (reg671 ? reg238 : reg1575)))));
              reg1589 <= ($unsigned(reg1533[(3'h4):(2'h3)]) <= ({(!(reg252 ~^ reg803)),
                  $signed($signed(reg1529)),
                  ((~^reg892) ?
                      reg606 : (reg472 ?
                          reg760 : reg730))} <<< $unsigned({(reg386 ?
                      reg480 : reg388)})));
              reg1590 = $signed({($signed($unsigned(reg671)) ?
                      ((~reg1562) ?
                          $unsigned(reg1562) : (reg430 | (7'h50))) : (~&$signed(reg360)))});
              reg1592 = {{(((reg846 ?
                              wire191 : reg199) > reg228[(2'h3):(2'h2)]) ?
                          {reg827[(3'h6):(1'h0)]} : reg646[(4'hf):(4'h9)]),
                      (!$unsigned({wire584}))},
                  {$signed((-(~^wire193)))}};
              reg1593 = (reg273[(5'h10):(2'h2)] ?
                  reg734 : ((reg341 >> $unsigned(reg1533[(5'h11):(2'h2)])) ?
                      (~|$signed((&forvar1585))) : (^((reg1533 ~^ reg863) << (8'hbe)))));
              reg1594 <= (+reg607);
            end
          for (forvar1595 = (1'h0); (forvar1595 < (3'h5)); forvar1595 = (forvar1595 + (1'h1)))
            begin
              reg1596 <= reg424;
              reg1597 = $signed((^(reg760 + $signed((reg657 ?
                  reg231 : (8'hac))))));
              reg1598 <= (reg436 && {($signed({reg597,
                      reg696}) >> (|(-reg362)))});
              reg1599 <= $unsigned($signed((((reg1587 >> (8'ha3)) ?
                      (reg655 < (8'hb6)) : (~&reg654)) ?
                  (reg853[(4'hc):(3'h4)] ?
                      (wire584 << reg1516) : ((8'hb0) ?
                          (8'hab) : reg218)) : (wire351[(5'h14):(3'h7)] & $signed((8'hb5))))));
              reg1600 <= ((({(!reg624),
                      $unsigned(reg462)} & {reg1576[(3'h6):(2'h3)],
                      (reg895 && reg1599)}) ?
                  reg460[(3'h7):(1'h0)] : $unsigned({(reg243 ?
                          reg330 : reg1586),
                      (7'h41),
                      reg316})) && ($unsigned(reg762) ?
                  (&{(reg745 << reg1534), $unsigned(reg1525)}) : reg785));
            end
          reg1601 = $unsigned(((($signed(reg866) & reg645) ?
              {(reg892 ?
                      (7'h54) : (7'h4a))} : reg713) ~^ reg491[(1'h1):(1'h0)]));
          for (forvar1602 = (1'h0); (forvar1602 < (3'h5)); forvar1602 = (forvar1602 + (1'h1)))
            begin
              reg1603 <= reg502[(3'h7):(2'h3)];
              reg1604 <= (~reg237[(1'h0):(1'h0)]);
              reg1605 <= (reg453[(3'h7):(1'h0)] > $signed(reg515[(2'h3):(2'h2)]));
              reg1606 <= reg850;
              reg1607 <= {(~|(((reg713 ^ (8'hb7)) ?
                          (reg879 >> reg331) : reg736[(3'h6):(2'h2)]) ?
                      $signed($unsigned(reg779)) : $signed((reg1572 >> (8'ha7)))))};
            end
          if (($signed(((^(reg343 ?
                  wire190 : reg316)) > reg199[(2'h3):(2'h2)])) ?
              ({reg468} ?
                  $signed((-{(8'hb3)})) : $unsigned({$signed(reg393),
                      $unsigned(reg889),
                      (reg330 ~^ reg474)})) : ((+$unsigned((reg1500 <= (8'hb4)))) <= reg256[(5'h1c):(4'ha)])))
            begin
              reg1608 = (|reg245);
            end
          else
            begin
              reg1609 <= {(($unsigned((reg672 ? reg744 : reg199)) ?
                          {$signed(reg1593),
                              reg1528,
                              forvar1595[(4'ha):(1'h0)]} : ($signed(reg779) ?
                              (reg606 < reg844) : (~&reg494))) ?
                      $unsigned({reg338[(2'h2):(2'h2)],
                          reg255[(2'h2):(1'h0)]}) : {(wire192 + (reg847 != reg597)),
                          $signed((7'h4d))}),
                  reg1593[(1'h0):(1'h0)]};
              reg1610 <= $unsigned(reg484[(1'h1):(1'h0)]);
              reg1611 = ($unsigned($unsigned(((reg335 ^ reg501) ?
                      (^~reg1571) : reg859))) ?
                  $unsigned((^~((reg736 ?
                      reg607 : reg808) && $unsigned(reg483)))) : reg734);
              reg1612 <= $signed((8'hbd));
            end
        end
    end
  assign wire1613 = ((+reg1534) && (+wire192));
  always
    @(posedge clk) begin
      if (((reg491[(2'h2):(2'h2)] ?
          $signed($unsigned($unsigned(reg312))) : reg1529[(3'h4):(2'h2)]) << ({((reg795 ?
                  reg589 : (8'ha9)) << (reg769 ? (8'haa) : reg276)),
              $unsigned($unsigned((7'h50))),
              $signed((reg815 || reg398))} ?
          $signed(reg1609[(1'h1):(1'h1)]) : reg774)))
        begin
          if ((reg779 & $signed(reg366)))
            begin
              reg1614 <= (reg828[(5'h12):(1'h1)] ?
                  ($unsigned(reg1607[(5'h15):(5'h12)]) << reg496[(5'h17):(1'h1)]) : reg1600);
              reg1615 <= reg1559[(3'h6):(3'h6)];
              reg1616 = $signed(reg245[(2'h2):(2'h2)]);
              reg1617 <= (-(~{{(reg445 ~^ reg462), {reg1501, reg616}},
                  (~(reg1600 ? reg256 : reg1532))}));
              reg1618 <= $signed((~&{(|reg837[(4'hf):(4'he)])}));
            end
          else
            begin
              reg1616 = (($unsigned({(reg672 ? reg1562 : reg346),
                          (reg635 ? reg874 : reg1528),
                          (reg299 ^~ reg673)}) ?
                      reg424[(4'ha):(4'ha)] : {$unsigned((wire192 - (8'hb7)))}) ?
                  $signed(reg460[(2'h2):(1'h1)]) : reg809);
              reg1619 = (~^{reg1580});
              reg1620 <= $unsigned($unsigned((reg480[(4'hf):(4'h9)] == $signed(reg472))));
              reg1621 <= ($unsigned(({(reg879 ? reg509 : (8'ha0)),
                          (reg604 != reg1532)} ?
                      reg346[(3'h4):(2'h3)] : $signed(reg593))) ?
                  (~|$unsigned(reg383[(5'h1f):(4'hb)])) : reg398[(3'h7):(1'h1)]);
            end
          reg1622 = $unsigned($signed({(-reg1600),
              $signed(reg597[(2'h2):(1'h0)]),
              ((reg1548 ? reg493 : reg237) < reg312)}));
          for (forvar1623 = (1'h0); (forvar1623 < (3'h6)); forvar1623 = (forvar1623 + (1'h1)))
            begin
              reg1624 = {((~^reg744) >= {wire195[(3'h6):(2'h2)],
                      ((7'h42) ?
                          (reg1576 ? reg610 : reg1614) : {reg430,
                              (7'h40),
                              reg511}),
                      $signed({reg1618, reg750, reg287})}),
                  $unsigned((8'hb0))};
              reg1625 = (8'hae);
              reg1626 = reg783;
              reg1627 <= (reg832 ?
                  $unsigned({(^~reg399)}) : (reg515[(1'h1):(1'h0)] ?
                      (~^((&reg514) ? $signed(reg1558) : (~reg589))) : reg587));
              reg1628 = reg320;
              reg1629 = (~|($unsigned(reg339) ^ reg453));
              reg1630 = (&{((reg674 ?
                      $signed(reg895) : reg484[(3'h5):(1'h0)]) || $signed((reg1599 >= reg388))),
                  $unsigned(reg813[(3'h7):(2'h3)])});
            end
          for (forvar1631 = (1'h0); (forvar1631 < (2'h2)); forvar1631 = (forvar1631 + (1'h1)))
            begin
              reg1632 <= ((+reg389[(1'h1):(1'h0)]) ?
                  reg373[(4'hb):(4'ha)] : reg227[(3'h6):(1'h1)]);
              reg1633 = (((((~&reg321) >= $unsigned(reg343)) == (reg462 == reg592)) ~^ reg884[(4'hb):(2'h3)]) ?
                  $signed($unsigned($unsigned((reg1562 ?
                      (8'ha0) : reg1591)))) : (-reg203[(3'h5):(2'h3)]));
            end
          for (forvar1634 = (1'h0); (forvar1634 < (3'h5)); forvar1634 = (forvar1634 + (1'h1)))
            begin
              reg1635 = $signed($signed(((^$signed(reg1596)) ^ reg769)));
              reg1636 <= (~&(reg659 && {$unsigned((reg1596 ? reg833 : reg643)),
                  {reg210[(2'h2):(2'h2)]},
                  reg671}));
            end
          if ((+(reg742[(1'h0):(1'h0)] ? reg245 : reg889[(3'h4):(2'h3)])))
            begin
              reg1637 <= reg434;
              reg1638 = ($unsigned($signed(reg1605[(5'h19):(2'h2)])) <= $signed(reg1600));
            end
          else
            begin
              reg1637 <= $signed(reg745);
              reg1638 = (((reg600[(2'h3):(2'h2)] ^ reg1604) ^ $unsigned((~{reg742,
                  wire717}))) < $signed((reg440 - {(reg238 ? reg1617 : reg785),
                  (7'h47),
                  reg1599})));
              reg1639 = ((reg778 ^ (!$unsigned(reg435[(3'h4):(2'h3)]))) ^ reg645);
              reg1640 = reg265[(1'h0):(1'h0)];
            end
          for (forvar1641 = (1'h0); (forvar1641 < (3'h4)); forvar1641 = (forvar1641 + (1'h1)))
            begin
              reg1642 = (7'h46);
              reg1643 <= {reg403[(4'h8):(3'h4)]};
              reg1644 <= reg462;
              reg1645 = reg1549[(3'h6):(1'h1)];
              reg1646 <= $signed(reg837[(4'h8):(2'h2)]);
              reg1647 <= $signed((~((reg1642[(5'h13):(5'h11)] ?
                  $signed(reg316) : {(7'h4c)}) <= (^~reg741[(4'hb):(2'h2)]))));
              reg1648 = ((~^(reg313 ?
                      (!reg745) : (reg787[(3'h7):(3'h6)] * $signed(reg300)))) ?
                  ((&$signed({reg850, reg268, reg597})) ?
                      $signed(($signed(reg789) ?
                          reg1587[(2'h2):(2'h2)] : {(7'h4f),
                              (8'hbe)})) : reg256) : forvar1641[(2'h2):(1'h1)]);
            end
        end
      else
        begin
          for (forvar1614 = (1'h0); (forvar1614 < (1'h1)); forvar1614 = (forvar1614 + (1'h1)))
            begin
              reg1616 = (8'hb0);
            end
          reg1619 = reg672[(5'h11):(3'h7)];
          reg1620 <= reg704;
        end
      reg1649 <= reg842;
      for (forvar1650 = (1'h0); (forvar1650 < (1'h1)); forvar1650 = (forvar1650 + (1'h1)))
        begin
          if ($unsigned($signed(reg707)))
            begin
              reg1651 <= $signed($signed($signed(($signed((7'h48)) && (~^(8'hb6))))));
              reg1652 = $unsigned((reg330[(3'h4):(2'h2)] ?
                  $unsigned($unsigned(reg1639)) : {reg858[(3'h7):(3'h6)],
                      ((8'had) <<< $signed(reg252)),
                      {$unsigned(reg700)}}));
              reg1653 = reg1646[(1'h1):(1'h0)];
              reg1654 <= (({reg1551} ?
                      wire351[(4'hb):(4'ha)] : $signed(reg403[(5'h1a):(2'h3)])) ?
                  (-$signed(($signed((8'had)) ?
                      reg492 : $signed(reg249)))) : ($unsigned((|(reg592 ?
                      reg1629 : reg774))) * ($signed(reg1583[(2'h2):(1'h1)]) > $unsigned((reg1647 ?
                      reg206 : (8'haf))))));
            end
          else
            begin
              reg1651 <= $signed(reg1550);
              reg1654 <= {reg284, reg872};
              reg1655 <= reg359[(3'h4):(2'h2)];
              reg1656 = (({$unsigned($unsigned(reg280)),
                      ((reg627 ? reg341 : (8'hbb)) ?
                          (reg884 ? reg403 : (8'hbe)) : reg801),
                      $signed($signed(reg494))} >= {(~&(!reg416)),
                      $unsigned((+reg231)),
                      $unsigned((8'hab))}) ?
                  (reg726[(4'hd):(1'h1)] ?
                      {(reg435 ? (reg604 | reg511) : (-wire718)),
                          $signed((reg319 > reg672)),
                          $unsigned(((8'hae) ?
                              reg1558 : reg501))} : $unsigned($signed($unsigned(reg1527)))) : reg801);
              reg1657 <= {(8'hb4),
                  $unsigned($unsigned(({reg1639, reg199} ?
                      reg1572[(2'h2):(1'h1)] : (^reg1644)))),
                  $signed(reg1501[(2'h3):(2'h2)])};
              reg1658 <= reg1624;
              reg1659 = reg1599;
            end
          reg1660 = ((~^reg359) - $unsigned((~&reg1635)));
          for (forvar1661 = (1'h0); (forvar1661 < (3'h5)); forvar1661 = (forvar1661 + (1'h1)))
            begin
              reg1662 = (((~^$unsigned(reg828[(2'h3):(1'h1)])) ?
                  ((|(reg1533 == (8'hab))) ?
                      reg203[(3'h7):(3'h5)] : $signed((reg265 * reg313))) : reg1652[(4'he):(1'h0)]) & wire194);
              reg1663 = $unsigned($signed(reg801));
              reg1664 <= reg386[(2'h3):(1'h0)];
              reg1665 <= (+(wire195[(3'h4):(3'h4)] <= $signed(($signed(reg399) * $unsigned(forvar1650)))));
              reg1666 = $signed($unsigned($signed((~reg415[(4'hc):(3'h5)]))));
            end
          if (((reg263 ?
                  (-$unsigned(reg474)) : (((reg698 ?
                          (7'h50) : reg785) != reg483) ?
                      (|((8'ha4) > reg683)) : reg842[(5'h11):(1'h1)])) ?
              (8'hac) : ((^~{reg232}) & $unsigned(reg589[(3'h5):(2'h2)]))))
            begin
              reg1667 = $signed((reg1644[(3'h4):(3'h4)] + reg1645));
              reg1668 <= reg731[(4'hb):(4'ha)];
            end
          else
            begin
              reg1668 <= ($unsigned(($signed($unsigned(reg501)) ?
                      $signed($unsigned(reg1539)) : $signed((reg776 ?
                          (7'h50) : reg613)))) ?
                  (reg399[(4'hc):(2'h2)] >>> reg736) : (8'ha7));
              reg1669 = reg1596[(1'h0):(1'h0)];
              reg1670 <= ((-(reg311 ?
                      (~$signed(reg837)) : $unsigned((reg745 ?
                          reg1580 : (8'haa))))) ?
                  reg1533 : (reg779[(5'h13):(3'h6)] ?
                      (^~((reg616 ?
                          reg1616 : (8'h9f)) <= $signed((8'ha8)))) : (~$signed((reg1548 ?
                          reg646 : wire194)))));
            end
          reg1671 <= (|(+reg1617));
        end
      if (reg496)
        begin
          if ($signed(($signed(reg808[(3'h4):(1'h0)]) & (((reg1625 ?
                  reg1576 : wire1494) ~^ reg330) ?
              reg513[(1'h1):(1'h1)] : (7'h4d)))))
            begin
              reg1672 = {reg673,
                  ((({reg474} | wire351[(5'h11):(2'h3)]) ?
                      (~&$unsigned((7'h41))) : ($signed((7'h56)) ?
                          (reg331 ?
                              reg870 : reg1517) : $unsigned(reg779))) < $signed({{(7'h49)},
                      $unsigned(reg480)}))};
            end
          else
            begin
              reg1673 <= reg307[(1'h0):(1'h0)];
              reg1674 = reg373;
              reg1675 <= (+(reg1669[(5'h15):(4'h8)] ^~ ((7'h4a) ?
                  {(|reg781),
                      $signed(reg639),
                      (reg371 ? reg268 : (8'hb5))} : ({(7'h41),
                      reg416,
                      reg760} * (reg657 ? reg503 : (8'hb2))))));
            end
          for (forvar1676 = (1'h0); (forvar1676 < (3'h4)); forvar1676 = (forvar1676 + (1'h1)))
            begin
              reg1677 <= {reg1599,
                  (+reg1598[(2'h2):(1'h1)]),
                  (reg1607[(5'h19):(4'hd)] ?
                      {reg650[(4'ha):(3'h7)],
                          ({forvar1623} ?
                              (reg1637 ? reg1619 : reg1635) : (reg270 ?
                                  reg269 : reg1507)),
                          reg879[(5'h18):(3'h6)]} : reg728)};
            end
          reg1678 = ($signed({$signed((wire194 > reg1591)),
                  (reg470[(4'hf):(4'he)] << reg853[(1'h0):(1'h0)]),
                  (^reg763[(4'hd):(4'h8)])}) ?
              (^reg1525) : $unsigned({((^~reg484) ?
                      {reg1563, reg1655, (7'h43)} : (|reg210)),
                  ((reg1612 >> reg793) | ((8'hae) << reg1534)),
                  ($signed(reg484) - $signed(reg505))}));
          reg1679 <= ($unsigned($unsigned(reg884)) ?
              reg512[(4'he):(4'hc)] : {(&(!reg597))});
          reg1680 <= {(|reg724[(4'he):(3'h5)]), reg1616, {reg796}};
        end
      else
        begin
          reg1673 <= (((^~$signed((~|reg313))) ?
                  reg436[(4'he):(4'hd)] : forvar1634[(4'hd):(1'h0)]) ?
              (|((+$unsigned((8'hb3))) ?
                  reg809[(4'hd):(3'h7)] : ({(7'h48),
                      reg265,
                      reg255} << reg602))) : {{(^reg494),
                      (+reg773[(1'h0):(1'h0)])},
                  (reg744[(1'h1):(1'h0)] + ((wire351 >= reg359) ?
                      reg1667[(5'h1c):(5'h1b)] : $signed(reg726))),
                  (8'hb6)});
          for (forvar1674 = (1'h0); (forvar1674 < (3'h6)); forvar1674 = (forvar1674 + (1'h1)))
            begin
              reg1676 = reg1627[(5'h1c):(3'h7)];
              reg1677 <= reg750[(5'h1a):(4'h9)];
            end
          reg1679 <= reg1594;
          reg1681 = {reg1555};
          for (forvar1682 = (1'h0); (forvar1682 < (3'h5)); forvar1682 = (forvar1682 + (1'h1)))
            begin
              reg1683 <= reg1578[(2'h3):(2'h2)];
              reg1684 = (^reg597[(1'h0):(1'h0)]);
              reg1685 = (reg1645[(3'h4):(2'h2)] ?
                  $signed(($unsigned((~^reg1655)) ?
                      ({reg774} || ((7'h47) ?
                          reg872 : reg781)) : ((^reg782) <<< (reg884 ?
                          reg280 : forvar1634)))) : $unsigned((&($signed(reg1662) ?
                      $signed((8'haf)) : forvar1641[(3'h5):(3'h4)]))));
              reg1686 <= $unsigned($unsigned(reg798));
            end
          if (reg699[(3'h5):(3'h5)])
            begin
              reg1687 = $signed(((($signed(reg360) ?
                          $signed(reg866) : forvar1650) ?
                      ((~^reg1635) ? reg256 : $signed(reg430)) : reg335) ?
                  reg238 : ((&reg1681) || (!(reg210 ? (7'h4b) : reg783)))));
              reg1688 <= {reg345[(4'hd):(3'h4)]};
              reg1689 = $signed(reg1670);
              reg1690 <= (^$unsigned(reg880));
              reg1691 = reg654[(2'h2):(2'h2)];
              reg1692 = forvar1641[(3'h6):(3'h5)];
            end
          else
            begin
              reg1688 <= (reg864 ?
                  ($signed($unsigned($unsigned(reg1687))) ?
                      $signed($signed((^~reg299))) : ((~(8'hb0)) - (+(~^reg818)))) : reg483[(3'h7):(3'h5)]);
              reg1690 <= (reg889 != reg671);
              reg1691 = ((^(reg421 < reg602)) ?
                  $unsigned($unsigned(({reg698} >= reg1692))) : $unsigned(reg652[(3'h6):(2'h3)]));
            end
          for (forvar1693 = (1'h0); (forvar1693 < (3'h4)); forvar1693 = (forvar1693 + (1'h1)))
            begin
              reg1694 <= {$unsigned(reg1559[(1'h1):(1'h1)])};
              reg1695 <= (8'ha4);
              reg1696 <= $unsigned((({(reg607 - reg846), reg1580} ?
                      {$signed(reg218),
                          {reg1678, (7'h57), reg1525},
                          $unsigned(reg879)} : $signed(reg796[(3'h7):(1'h1)])) ?
                  $unsigned((~&(reg627 == reg371))) : (+$signed($signed(reg238)))));
            end
        end
    end
  assign wire1697 = $signed($signed(reg639[(4'h8):(3'h6)]));
  always
    @(posedge clk) begin
      for (forvar1698 = (1'h0); (forvar1698 < (3'h5)); forvar1698 = (forvar1698 + (1'h1)))
        begin
          if (reg1576)
            begin
              reg1699 = (~^(8'hbd));
              reg1700 <= $unsigned($signed((($signed(reg399) ?
                      $signed(reg705) : $signed(reg324)) ?
                  ({reg884, (8'hb2)} * (reg507 ?
                      reg360 : reg1617)) : $unsigned(reg1533[(1'h0):(1'h0)]))));
              reg1701 = $unsigned({reg728,
                  reg287[(4'hb):(4'h8)],
                  ((~&(reg832 ? (8'ha5) : wire191)) != reg635)});
            end
          else
            begin
              reg1699 = (reg741 <<< $signed((^~$signed(reg832))));
              reg1700 <= wire195;
              reg1701 = {reg1680};
              reg1702 = ((&((&(reg707 ?
                      (8'hbc) : reg484)) < $unsigned(reg470))) ?
                  {(reg429[(2'h3):(2'h3)] ?
                          reg1594[(4'hf):(3'h5)] : $signed((reg327 >> reg216))),
                      ({(reg880 != reg650),
                          (reg313 ~^ reg373)} <<< $signed($signed(reg1497)))} : (8'haf));
            end
          for (forvar1703 = (1'h0); (forvar1703 < (2'h3)); forvar1703 = (forvar1703 + (1'h1)))
            begin
              reg1704 = (({reg496[(5'h14):(1'h1)],
                          $unsigned($signed(reg1598)),
                          reg283} ?
                      (~|{(~&reg468)}) : (($unsigned((7'h41)) ?
                              (reg1584 ? reg440 : reg324) : $unsigned(reg702)) ?
                          (-reg1548) : ((wire194 ?
                              reg1532 : reg434) != $unsigned(reg1501)))) ?
                  (reg236[(3'h7):(1'h1)] * ((-reg863[(4'hc):(4'ha)]) ?
                      ($signed(reg745) | (reg370 ?
                          reg810 : reg206)) : (+(~^reg321)))) : $signed(reg1683[(3'h4):(1'h1)]));
              reg1705 <= $signed($unsigned(reg483));
              reg1706 = {reg742,
                  ($unsigned((reg299[(4'hb):(3'h5)] ^ (reg210 ?
                      (8'hbe) : reg763))) - $unsigned(reg871[(3'h6):(3'h4)]))};
              reg1707 = {(^reg762),
                  reg312,
                  ($unsigned((+((7'h49) + (7'h51)))) ?
                      ((^(reg421 ?
                          reg210 : reg1657)) <= $unsigned((~reg269))) : $unsigned(((reg1558 ?
                              reg1514 : reg708) ?
                          (8'hb9) : $unsigned((8'ha1)))))};
              reg1708 <= $unsigned(($signed(reg470[(4'h9):(2'h3)]) ?
                  (~&$signed((reg699 ?
                      reg494 : reg850))) : ({$unsigned(reg1705),
                          reg1554[(4'hb):(4'hb)],
                          reg492[(1'h1):(1'h1)]} ?
                      $signed((!(8'h9d))) : reg1562[(4'ha):(1'h1)])));
            end
          for (forvar1709 = (1'h0); (forvar1709 < (1'h1)); forvar1709 = (forvar1709 + (1'h1)))
            begin
              reg1710 = $signed(({reg283[(1'h0):(1'h0)],
                  (^(wire350 ? reg745 : reg475)),
                  {reg313, $signed(reg259)}} <= (8'hae)));
            end
          for (forvar1711 = (1'h0); (forvar1711 < (3'h4)); forvar1711 = (forvar1711 + (1'h1)))
            begin
              reg1712 <= reg742[(2'h3):(2'h2)];
              reg1713 = (+(({$unsigned((8'ha1)),
                          ((8'ha1) ? reg300 : reg1572),
                          (wire351 ? reg388 : reg1591)} ?
                      $unsigned(((7'h43) ?
                          (7'h48) : reg210)) : reg287[(4'he):(4'h9)]) ?
                  $unsigned((!$unsigned(reg741))) : (((reg1670 ?
                          reg462 : (8'hac)) ?
                      {reg696,
                          reg778,
                          reg775} : (~|reg493)) << reg853[(4'he):(1'h1)])));
              reg1714 <= $unsigned(reg484[(1'h0):(1'h0)]);
              reg1715 = reg589;
              reg1716 = reg389[(2'h2):(2'h2)];
            end
        end
      if (((7'h44) ?
          (7'h56) : {(-$signed(reg276)),
              (~|($signed(reg592) + (~reg878))),
              (^((reg1587 >> reg593) ? (reg415 - reg1713) : {(8'hb7)}))}))
        begin
          if (({$unsigned($signed((reg834 ? reg1600 : reg1552)))} ?
              (|(~reg671[(2'h2):(1'h0)])) : $unsigned(reg652)))
            begin
              reg1717 <= $signed((^~(8'hb2)));
              reg1718 = {$unsigned($signed((&reg597[(1'h1):(1'h1)])))};
              reg1719 <= $unsigned(reg483[(2'h2):(1'h1)]);
              reg1720 = ((!reg364[(2'h2):(1'h0)]) ~^ {$signed(reg362[(5'h13):(4'ha)])});
              reg1721 <= (($unsigned((reg638[(5'h10):(4'h9)] ?
                  (reg773 <<< reg841) : wire754[(1'h0):(1'h0)])) <= (^reg218[(4'hd):(1'h0)])) & (8'hb3));
              reg1722 <= ($signed((reg589[(5'h13):(1'h1)] == (reg393 ?
                  reg781 : $signed((8'haf))))) & $signed(({$unsigned((8'hbb)),
                  {reg1696, reg1524},
                  reg1694} < $signed($signed(reg1670)))));
            end
          else
            begin
              reg1718 = $signed((&{((reg674 ? reg1554 : (8'hab)) ?
                      (+reg879) : reg1665),
                  $signed($signed(reg362))}));
              reg1719 <= (wire584[(2'h2):(1'h0)] ?
                  reg880 : $signed(reg371[(3'h4):(1'h0)]));
              reg1721 <= $signed((&reg827));
              reg1723 = $unsigned(reg828);
              reg1724 <= reg1525;
              reg1725 <= reg345;
              reg1726 <= $signed((!$unsigned(reg462)));
            end
          reg1727 = ({reg1712, $signed((~(8'hbd))), reg839[(2'h3):(2'h3)]} ?
              $unsigned(reg507) : $unsigned((reg389 * ($unsigned((8'hb2)) ?
                  $unsigned(reg258) : (reg205 ? (8'hb5) : reg728)))));
          for (forvar1728 = (1'h0); (forvar1728 < (3'h5)); forvar1728 = (forvar1728 + (1'h1)))
            begin
              reg1729 = {reg773[(2'h2):(1'h1)],
                  ($unsigned((reg1664 ^ $signed(reg846))) || (^~((reg206 ?
                      (8'h9d) : reg307) + (reg627 * reg1560))))};
              reg1730 = $unsigned(({$signed(reg1702[(1'h0):(1'h0)])} ?
                  (reg1720[(3'h5):(2'h2)] >> (+reg1644[(2'h3):(2'h2)])) : $unsigned(((&reg1651) < reg602))));
              reg1731 <= (^~({(7'h4c),
                  $unsigned(reg1594)} >>> reg698[(5'h17):(5'h11)]));
              reg1732 <= {reg805[(4'h8):(3'h5)], reg1665[(5'h10):(1'h0)]};
              reg1733 <= ($unsigned($signed(reg1614)) ?
                  reg1688[(5'h17):(4'h9)] : reg429[(3'h6):(3'h6)]);
              reg1734 <= ((reg252 >= (-(reg444[(5'h13):(4'ha)] >>> {reg201,
                  reg1701,
                  reg359}))) & ((8'ha3) ? reg638[(4'hd):(1'h0)] : reg1688));
            end
        end
      else
        begin
          reg1718 = reg1675;
          for (forvar1719 = (1'h0); (forvar1719 < (2'h2)); forvar1719 = (forvar1719 + (1'h1)))
            begin
              reg1721 <= $unsigned(($unsigned(reg436[(3'h4):(1'h0)]) != ((~{reg287,
                      reg1600,
                      (7'h56)}) ?
                  $signed((~|(7'h48))) : $unsigned((reg324 ?
                      wire194 : reg345)))));
              reg1723 = $signed((-reg1603));
              reg1727 = (reg225 >>> reg587);
              reg1728 <= reg1718[(2'h2):(1'h1)];
            end
        end
      for (forvar1735 = (1'h0); (forvar1735 < (3'h6)); forvar1735 = (forvar1735 + (1'h1)))
        begin
          reg1736 = (-$unsigned($signed(((^reg1527) ?
              wire1613[(4'hf):(2'h2)] : (reg648 >> reg402)))));
          reg1737 = (&$unsigned(((reg1733 ?
              (reg704 & reg833) : {reg641}) >> (~^reg268[(3'h5):(1'h1)]))));
        end
      reg1738 <= {wire192};
    end
  assign wire1739 = (8'hb3);
  always
    @(posedge clk) begin
      if ((reg424 ?
          ((reg252 * $unsigned((reg782 ?
              reg1615 : reg664))) ^ $unsigned((+(reg494 ?
              reg1670 : reg853)))) : reg696))
        begin
          reg1740 <= ((reg228[(3'h6):(3'h6)] ?
                  {{{reg1552}, (wire1739 == reg744), reg767},
                      $signed((reg1694 ? reg503 : reg435)),
                      reg389[(1'h1):(1'h0)]} : (((&reg278) ?
                      {reg1614,
                          reg805} : reg871[(3'h4):(1'h1)]) != $signed((~^reg507)))) ?
              (~&(|reg1550)) : (~reg456[(1'h0):(1'h0)]));
          reg1741 <= reg307[(4'hc):(4'ha)];
          if ({$signed({(((7'h4c) ?
                      reg491 : reg1632) != reg1566[(5'h1b):(4'hf)])})})
            begin
              reg1742 <= ((~$unsigned(((^reg1696) && $signed((7'h48))))) ?
                  ((reg1670[(3'h6):(2'h3)] ?
                          ((reg249 ? reg208 : (7'h50)) ?
                              {reg1508} : (reg872 || reg515)) : ($signed(reg604) ?
                              $signed(reg393) : $signed(reg1532))) ?
                      ($signed($signed(reg399)) ?
                          reg664 : (!reg652)) : $signed(reg832[(1'h0):(1'h0)])) : {$unsigned((~&reg300))});
              reg1743 = $signed($unsigned((8'ha2)));
              reg1744 <= $signed(reg346[(1'h1):(1'h1)]);
              reg1745 = (reg773 && (&$signed(reg203[(5'h10):(4'ha)])));
              reg1746 = reg1725;
            end
          else
            begin
              reg1743 = {reg1591,
                  ($signed(((~&reg657) ?
                      reg1594[(4'hc):(3'h4)] : $signed(wire350))) && $unsigned(reg278)),
                  ((reg480 << (reg319 ?
                      {reg1598,
                          reg1705} : (+reg365))) >>> (((reg783 <= reg1594) ?
                          $unsigned(wire718) : (reg589 ? reg1695 : reg864)) ?
                      (reg316 == {reg1500, reg779, reg330}) : ({reg474,
                          reg403,
                          reg1686} | (+reg280))))};
              reg1745 = {((reg1580[(1'h0):(1'h0)] ?
                      reg335 : (8'hb1)) << reg1717),
                  $signed($signed(({reg341, reg703} ?
                      $signed(reg734) : $unsigned((7'h4a))))),
                  ({(^~reg511),
                      $signed(reg648)} ~^ (+$signed($signed(reg808))))};
            end
          for (forvar1747 = (1'h0); (forvar1747 < (3'h5)); forvar1747 = (forvar1747 + (1'h1)))
            begin
              reg1748 = (((~^$unsigned($unsigned(reg287))) >> {$unsigned((&reg1673))}) <<< (8'hbc));
            end
        end
      else
        begin
          for (forvar1740 = (1'h0); (forvar1740 < (1'h1)); forvar1740 = (forvar1740 + (1'h1)))
            begin
              reg1741 <= {(8'ha2),
                  reg589[(3'h7):(3'h5)],
                  $signed(reg1548[(5'h18):(3'h5)])};
              reg1743 = wire1697;
              reg1744 <= {(reg1514 ?
                      (reg793[(1'h1):(1'h0)] | (+(reg892 > reg837))) : reg850[(3'h4):(2'h3)]),
                  (reg424[(5'h11):(4'he)] & ($unsigned(reg386) ?
                      (&(reg881 <= (7'h56))) : ((+reg1683) ?
                          reg713 : $unsigned(reg453)))),
                  (~$unsigned(((reg793 ?
                      (7'h40) : reg503) * $signed(reg345))))};
              reg1745 = ($signed((~|$signed((reg813 > reg341)))) - ($unsigned($unsigned($signed((8'ha4)))) ?
                  ({$unsigned(reg1532),
                      (wire1494 < reg1596)} & reg872) : {reg818,
                      (((8'ha3) * (8'had)) ? (+(7'h53)) : reg654)}));
              reg1747 <= (reg501 >>> $unsigned((&(+$unsigned(reg653)))));
              reg1748 = $unsigned($signed($unsigned(reg653)));
            end
          reg1749 = $unsigned((reg364[(2'h3):(1'h0)] ?
              (8'hb3) : $unsigned($unsigned($unsigned(reg491)))));
          if ({reg330})
            begin
              reg1750 = reg844[(4'hf):(4'he)];
              reg1751 = {(reg512 ? (~&(7'h4c)) : wire193),
                  {$signed(reg635)},
                  ($unsigned((~^$signed(reg1527))) ^ $signed((!$unsigned(reg1632))))};
              reg1752 <= ((^~($signed(reg225[(3'h5):(1'h1)]) ^~ ({reg1537,
                      reg617,
                      reg345} ?
                  reg258 : (8'ha3)))) <<< ((~&(8'ha0)) << $unsigned($unsigned((reg1738 > reg509)))));
              reg1753 <= reg436[(3'h7):(3'h4)];
              reg1754 = reg795;
            end
          else
            begin
              reg1752 <= {(~^reg707),
                  ($unsigned(reg881[(4'hd):(1'h0)]) == $unsigned((-reg892[(5'h18):(5'h12)])))};
              reg1754 = $unsigned((({{reg1554},
                      reg1523,
                      {reg1500, reg1594, reg1603}} ?
                  (^reg727[(1'h0):(1'h0)]) : (~&(reg265 << reg881))) ~^ $signed(reg370[(2'h2):(1'h0)])));
              reg1755 <= $unsigned(reg842);
            end
          reg1756 = (!$unsigned($unsigned((&$unsigned(reg317)))));
          if ((7'h42))
            begin
              reg1757 <= forvar1740;
            end
          else
            begin
              reg1758 = (((~$unsigned((|reg669))) > $signed($unsigned((~&reg462)))) ?
                  reg1621[(1'h0):(1'h0)] : ({$unsigned(reg678[(3'h7):(3'h6)]),
                          $signed((^~reg757)),
                          $unsigned((~|reg364))} ?
                      ($unsigned((reg776 ?
                          reg672 : reg787)) ^ reg436[(2'h2):(1'h1)]) : (~^reg1578)));
              reg1759 = {(7'h56),
                  (~|(({(7'h4d), (8'ha8), reg252} ?
                      $signed(reg1514) : (~reg1738)) | ($signed((8'haa)) ?
                      (8'hbc) : reg1529))),
                  reg360[(5'h12):(4'he)]};
              reg1760 = ($signed($signed($signed((~^reg663)))) ^ (($unsigned($unsigned(reg643)) >>> ({(7'h42),
                      wire1697} ?
                  wire351 : (!reg435))) > {reg403,
                  reg446[(2'h3):(2'h2)],
                  {reg436[(3'h4):(2'h3)]}}));
              reg1761 <= reg727[(3'h5):(2'h2)];
              reg1762 <= $signed($unsigned((~|reg1632)));
              reg1763 = {(((reg199 ?
                      reg480 : (reg736 < reg1746)) >> $unsigned($unsigned(reg1600))) <= (&({reg1717,
                          reg502,
                          reg827} ?
                      (reg1679 ? reg589 : reg592) : (reg507 >>> reg1537)))),
                  {(($unsigned(reg801) ?
                          reg1527 : $unsigned(wire516)) - (|reg231)),
                      reg811[(5'h1b):(4'hc)]},
                  reg1627};
            end
          reg1764 = $unsigned((|reg424[(2'h3):(2'h2)]));
          reg1765 = (-$signed(reg324[(3'h4):(3'h4)]));
        end
      for (forvar1766 = (1'h0); (forvar1766 < (3'h6)); forvar1766 = (forvar1766 + (1'h1)))
        begin
          for (forvar1767 = (1'h0); (forvar1767 < (3'h5)); forvar1767 = (forvar1767 + (1'h1)))
            begin
              reg1768 = reg815;
              reg1769 = ($signed(($unsigned((reg1758 ? reg280 : reg505)) ?
                      ({(7'h44), reg587, reg1528} ?
                          ((7'h4c) >= (7'h4e)) : $signed(reg805)) : ((~^reg362) || {(8'ha3)}))) ?
                  ((~^reg702) < $unsigned(reg287)) : wire192[(2'h2):(1'h1)]);
            end
          reg1770 <= ($signed((reg359[(2'h2):(1'h0)] <= ((|reg327) >= reg813))) ?
              reg210[(2'h3):(2'h3)] : reg773[(4'h8):(3'h5)]);
          reg1771 = (~^(-(+(reg206 && (8'hbf)))));
        end
    end
  assign wire1772 = (7'h56);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module896
#(parameter param1491 = (((~(((8'hb7) - (8'hb0)) ? ((8'hba) ^~ (8'hb5)) : ((8'hb1) <<< (7'h4a)))) >> ((((8'hbf) > (8'hb5)) <<< ((8'h9e) ? (8'h9f) : (7'h56))) ^ (((8'h9d) ? (7'h54) : (7'h53)) && ((8'h9c) ? (8'ha2) : (8'hb4))))) ? (((|((8'hb4) << (8'hb8))) * (+((8'hb5) ? (7'h4c) : (7'h45)))) ? ((((8'hb2) & (8'hb8)) ^ ((7'h48) << (7'h41))) ? ((^~(7'h52)) ? {(8'h9f), (8'ha0)} : (^(8'ha0))) : {(&(8'hae))}) : (((+(8'ha7)) > ((7'h4d) ? (8'h9d) : (7'h53))) ? ((~&(7'h4e)) ^ {(8'hb4), (8'hb6)}) : ({(8'hba)} <= (&(7'h56))))) : (((~&(+(7'h55))) == (((7'h42) ? (8'h9d) : (8'ha9)) <<< {(8'h9c), (8'hb4), (7'h45)})) + (^~(~&((8'hb3) ? (8'hbf) : (8'hae)))))), 
parameter param1492 = (~(!(^({param1491} ? (8'hb5) : (param1491 + param1491))))), 
parameter param1493 = {param1491, (!(&{(8'hbd)})), ((&(((8'h9e) ? param1492 : param1492) ~^ param1491)) ^ param1492)})
(y, clk, wire897, wire898, wire899, wire900);
  output wire [(32'hd40):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire897;
  input wire signed [(5'h15):(1'h0)] wire898;
  input wire [(5'h12):(1'h0)] wire899;
  input wire signed [(4'hc):(1'h0)] wire900;
  wire signed [(5'h19):(1'h0)] wire1407;
  wire [(5'h10):(1'h0)] wire901;
  wire signed [(2'h3):(1'h0)] wire957;
  wire [(4'he):(1'h0)] wire976;
  wire [(5'h15):(1'h0)] wire977;
  wire signed [(4'hc):(1'h0)] wire978;
  wire [(5'h17):(1'h0)] wire1405;
  reg signed [(4'ha):(1'h0)] reg1490 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1489 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1486 = (1'h0);
  reg [(5'h14):(1'h0)] reg1484 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1483 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1482 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1480 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1479 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1477 = (1'h0);
  reg [(2'h3):(1'h0)] reg1476 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1475 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1472 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1468 = (1'h0);
  reg [(3'h5):(1'h0)] reg1467 = (1'h0);
  reg [(5'h10):(1'h0)] reg1466 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1465 = (1'h0);
  reg [(5'h16):(1'h0)] reg1463 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1456 = (1'h0);
  reg [(3'h5):(1'h0)] reg1455 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1450 = (1'h0);
  reg [(3'h6):(1'h0)] reg1449 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1446 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1445 = (1'h0);
  reg [(5'h19):(1'h0)] reg1443 = (1'h0);
  reg [(5'h14):(1'h0)] reg1442 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1441 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1440 = (1'h0);
  reg [(3'h6):(1'h0)] reg1439 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1436 = (1'h0);
  reg [(4'h8):(1'h0)] reg1434 = (1'h0);
  reg [(3'h5):(1'h0)] reg1433 = (1'h0);
  reg [(5'h13):(1'h0)] reg1427 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1422 = (1'h0);
  reg [(5'h11):(1'h0)] reg1420 = (1'h0);
  reg [(4'hc):(1'h0)] reg1418 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1417 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1415 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1414 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1412 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1411 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1409 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1408 = (1'h0);
  reg [(4'h9):(1'h0)] reg1004 = (1'h0);
  reg [(4'he):(1'h0)] reg1002 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1000 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg998 = (1'h0);
  reg [(5'h18):(1'h0)] reg997 = (1'h0);
  reg [(3'h6):(1'h0)] reg995 = (1'h0);
  reg [(3'h7):(1'h0)] reg994 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg993 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg992 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg991 = (1'h0);
  reg [(4'h8):(1'h0)] reg989 = (1'h0);
  reg [(5'h18):(1'h0)] reg988 = (1'h0);
  reg [(5'h15):(1'h0)] reg986 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg984 = (1'h0);
  reg [(5'h10):(1'h0)] reg983 = (1'h0);
  reg [(2'h2):(1'h0)] reg980 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg975 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg973 = (1'h0);
  reg [(5'h17):(1'h0)] reg972 = (1'h0);
  reg [(5'h1b):(1'h0)] reg971 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg968 = (1'h0);
  reg [(4'he):(1'h0)] reg966 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg965 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg963 = (1'h0);
  reg [(5'h14):(1'h0)] reg962 = (1'h0);
  reg [(5'h1f):(1'h0)] reg960 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg954 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg952 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg951 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg949 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg946 = (1'h0);
  reg [(5'h13):(1'h0)] reg944 = (1'h0);
  reg [(5'h1d):(1'h0)] reg943 = (1'h0);
  reg [(5'h15):(1'h0)] reg940 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg937 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg936 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg932 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg931 = (1'h0);
  reg [(2'h2):(1'h0)] reg930 = (1'h0);
  reg [(5'h1f):(1'h0)] reg928 = (1'h0);
  reg [(5'h16):(1'h0)] reg927 = (1'h0);
  reg [(3'h6):(1'h0)] reg923 = (1'h0);
  reg [(5'h1d):(1'h0)] reg921 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg920 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg918 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg915 = (1'h0);
  reg [(4'hc):(1'h0)] reg913 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg912 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg911 = (1'h0);
  reg [(5'h1d):(1'h0)] reg905 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg904 = (1'h0);
  reg [(4'hd):(1'h0)] reg902 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1482 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1488 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1487 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1485 = (1'h0);
  reg [(5'h10):(1'h0)] reg1481 = (1'h0);
  reg [(5'h18):(1'h0)] reg1478 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1474 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1473 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1471 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1470 = (1'h0);
  reg [(4'ha):(1'h0)] reg1464 = (1'h0);
  reg [(4'he):(1'h0)] reg1462 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1461 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1460 = (1'h0);
  reg [(4'he):(1'h0)] forvar1459 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1458 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1457 = (1'h0);
  reg [(4'h9):(1'h0)] reg1454 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1453 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1452 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1451 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1448 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar1447 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1444 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1429 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1438 = (1'h0);
  reg [(5'h10):(1'h0)] reg1437 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1435 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1432 = (1'h0);
  reg [(5'h15):(1'h0)] reg1431 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1430 = (1'h0);
  reg [(2'h3):(1'h0)] reg1429 = (1'h0);
  reg [(5'h15):(1'h0)] reg1428 = (1'h0);
  reg [(5'h10):(1'h0)] reg1426 = (1'h0);
  reg [(5'h11):(1'h0)] reg1425 = (1'h0);
  reg [(5'h17):(1'h0)] reg1424 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1423 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1421 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1419 = (1'h0);
  reg [(3'h7):(1'h0)] reg1416 = (1'h0);
  reg [(5'h12):(1'h0)] reg1413 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar1410 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1003 = (1'h0);
  reg [(3'h6):(1'h0)] reg1001 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar999 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar996 = (1'h0);
  reg [(4'hc):(1'h0)] reg981 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar979 = (1'h0);
  reg [(4'hb):(1'h0)] reg990 = (1'h0);
  reg [(4'h9):(1'h0)] reg987 = (1'h0);
  reg [(2'h3):(1'h0)] reg985 = (1'h0);
  reg [(5'h16):(1'h0)] reg982 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar981 = (1'h0);
  reg [(5'h16):(1'h0)] reg979 = (1'h0);
  reg [(3'h7):(1'h0)] reg974 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg970 = (1'h0);
  reg [(5'h19):(1'h0)] forvar969 = (1'h0);
  reg [(4'hf):(1'h0)] reg967 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg964 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar961 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg959 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg958 = (1'h0);
  reg [(4'h9):(1'h0)] reg956 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar941 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg955 = (1'h0);
  reg [(5'h13):(1'h0)] reg953 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg950 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg948 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg947 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg945 = (1'h0);
  reg [(5'h15):(1'h0)] reg942 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg941 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar910 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg939 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg938 = (1'h0);
  reg [(3'h7):(1'h0)] reg935 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg934 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg933 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar929 = (1'h0);
  reg [(5'h1c):(1'h0)] reg926 = (1'h0);
  reg [(5'h1a):(1'h0)] reg925 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg924 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg922 = (1'h0);
  reg [(5'h1f):(1'h0)] reg919 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg917 = (1'h0);
  reg [(5'h14):(1'h0)] reg916 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg914 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg910 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg909 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg908 = (1'h0);
  reg [(5'h19):(1'h0)] forvar907 = (1'h0);
  reg [(3'h6):(1'h0)] reg906 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar903 = (1'h0);
  assign y = {wire1407,
                 wire901,
                 wire957,
                 wire976,
                 wire977,
                 wire978,
                 wire1405,
                 reg1490,
                 reg1489,
                 reg1486,
                 reg1484,
                 reg1483,
                 reg1482,
                 reg1480,
                 reg1479,
                 reg1477,
                 reg1476,
                 reg1475,
                 reg1472,
                 reg1469,
                 reg1468,
                 reg1467,
                 reg1466,
                 reg1465,
                 reg1463,
                 reg1456,
                 reg1455,
                 reg1450,
                 reg1449,
                 reg1446,
                 reg1445,
                 reg1443,
                 reg1442,
                 reg1441,
                 reg1440,
                 reg1439,
                 reg1436,
                 reg1434,
                 reg1433,
                 reg1427,
                 reg1422,
                 reg1420,
                 reg1418,
                 reg1417,
                 reg1415,
                 reg1414,
                 reg1412,
                 reg1411,
                 reg1409,
                 reg1408,
                 reg1004,
                 reg1002,
                 reg1000,
                 reg998,
                 reg997,
                 reg995,
                 reg994,
                 reg993,
                 reg992,
                 reg991,
                 reg989,
                 reg988,
                 reg986,
                 reg984,
                 reg983,
                 reg980,
                 reg975,
                 reg973,
                 reg972,
                 reg971,
                 reg968,
                 reg966,
                 reg965,
                 reg963,
                 reg962,
                 reg960,
                 reg954,
                 reg952,
                 reg951,
                 reg949,
                 reg946,
                 reg944,
                 reg943,
                 reg940,
                 reg937,
                 reg936,
                 reg932,
                 reg931,
                 reg930,
                 reg928,
                 reg927,
                 reg923,
                 reg921,
                 reg920,
                 reg918,
                 reg915,
                 reg913,
                 reg912,
                 reg911,
                 reg905,
                 reg904,
                 reg902,
                 forvar1482,
                 reg1488,
                 reg1487,
                 reg1485,
                 reg1481,
                 reg1478,
                 reg1474,
                 reg1473,
                 reg1471,
                 reg1470,
                 reg1464,
                 reg1462,
                 reg1461,
                 reg1460,
                 forvar1459,
                 reg1458,
                 reg1457,
                 reg1454,
                 forvar1453,
                 reg1452,
                 reg1451,
                 reg1448,
                 forvar1447,
                 forvar1444,
                 forvar1429,
                 reg1438,
                 reg1437,
                 reg1435,
                 reg1432,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1426,
                 reg1425,
                 reg1424,
                 forvar1423,
                 reg1421,
                 forvar1419,
                 reg1416,
                 reg1413,
                 forvar1410,
                 reg1003,
                 reg1001,
                 forvar999,
                 forvar996,
                 reg981,
                 forvar979,
                 reg990,
                 reg987,
                 reg985,
                 reg982,
                 forvar981,
                 reg979,
                 reg974,
                 reg970,
                 forvar969,
                 reg967,
                 reg964,
                 forvar961,
                 reg959,
                 reg958,
                 reg956,
                 forvar941,
                 reg955,
                 reg953,
                 reg950,
                 reg948,
                 reg947,
                 reg945,
                 reg942,
                 reg941,
                 forvar910,
                 reg939,
                 reg938,
                 reg935,
                 reg934,
                 reg933,
                 forvar929,
                 reg926,
                 reg925,
                 reg924,
                 reg922,
                 reg919,
                 reg917,
                 reg916,
                 reg914,
                 reg910,
                 reg909,
                 reg908,
                 forvar907,
                 reg906,
                 forvar903,
                 (1'h0)};
  assign wire901 = (7'h4c);
  always
    @(posedge clk) begin
      reg902 <= $unsigned((wire899[(2'h3):(1'h1)] ?
          (((~^wire898) - (wire900 ?
              wire900 : wire897)) + $unsigned(wire897)) : (wire898 ~^ $unsigned(wire901))));
      for (forvar903 = (1'h0); (forvar903 < (3'h4)); forvar903 = (forvar903 + (1'h1)))
        begin
          reg904 <= $signed((wire897 ^ forvar903));
          reg905 <= $unsigned((~(-$unsigned($unsigned(wire897)))));
          reg906 = forvar903;
          for (forvar907 = (1'h0); (forvar907 < (3'h4)); forvar907 = (forvar907 + (1'h1)))
            begin
              reg908 = ($signed(($signed((wire900 ~^ wire901)) & ((^wire900) && reg906))) ^~ ((+({reg904,
                          wire898} ?
                      reg905 : {reg904, wire900, reg902})) ?
                  wire897[(4'h8):(3'h7)] : reg902[(3'h5):(2'h3)]));
              reg909 = (($unsigned(reg908) > wire900[(1'h0):(1'h0)]) <= (reg905 ?
                  (~|wire898[(4'hd):(3'h7)]) : ((&(~|wire899)) ^ ({reg905,
                      reg906,
                      reg904} & wire897[(4'ha):(2'h3)]))));
            end
        end
    end
  always
    @(posedge clk) begin
      if ((($signed((~&(reg905 ? reg902 : reg904))) > wire899[(3'h4):(3'h4)]) ?
          ((((reg904 > wire899) >> wire897[(5'h10):(5'h10)]) - ($unsigned(reg904) >>> (wire901 >= wire897))) > wire901) : (+{(|$signed(wire901)),
              ($unsigned(wire898) - $unsigned(wire899)),
              ((wire898 << wire900) ~^ $unsigned(wire897))})))
        begin
          reg910 = $unsigned({(^~wire899[(3'h5):(1'h0)])});
          if (wire901[(3'h6):(1'h0)])
            begin
              reg911 <= $signed({{(reg905 >>> $signed((8'hb9))),
                      (wire899 ? $unsigned(wire900) : reg905),
                      reg910[(5'h14):(5'h14)]},
                  reg904[(1'h1):(1'h0)],
                  wire901});
              reg912 <= wire898[(1'h0):(1'h0)];
              reg913 <= (~$unsigned((8'hbc)));
              reg914 = wire897;
            end
          else
            begin
              reg914 = {$signed(((~|(reg905 ?
                      reg905 : reg904)) * (reg910[(5'h1a):(5'h16)] && $unsigned(wire897)))),
                  wire900[(2'h2):(1'h1)],
                  ($signed((^{reg913, (7'h4b), wire899})) ?
                      (^(8'ha7)) : (((^wire898) ^ wire897) ?
                          (reg912 + $unsigned(reg911)) : wire899))};
              reg915 <= reg905;
              reg916 = (reg910[(5'h15):(4'h8)] << ({$unsigned((reg912 < reg910)),
                      ((wire901 ^ (8'hb1)) ? (8'hb7) : {(8'ha8), reg910})} ?
                  $signed(reg913[(3'h6):(3'h5)]) : ($unsigned((reg911 ?
                          reg902 : reg904)) ?
                      $unsigned($unsigned(wire899)) : wire899)));
              reg917 = $signed(reg904[(1'h0):(1'h0)]);
              reg918 <= wire900;
              reg919 = $unsigned($signed((reg917 < reg914)));
            end
          if (($unsigned(wire898) ?
              (7'h43) : ($unsigned($signed((-wire900))) >>> reg914[(1'h1):(1'h0)])))
            begin
              reg920 <= (($unsigned({$unsigned(reg902), $unsigned(reg911)}) ?
                      (|$signed(wire899)) : $unsigned((^(reg910 * reg914)))) ?
                  wire901 : reg912[(5'h16):(4'ha)]);
              reg921 <= ((~(($unsigned(wire898) ?
                      (wire900 ? (8'hb2) : reg902) : $signed(wire900)) ?
                  $unsigned($signed(reg920)) : $signed($unsigned(wire899)))) && (!$signed(wire899[(4'h9):(3'h5)])));
              reg922 = (reg911 ?
                  {$signed((|{reg902,
                          reg912,
                          (7'h53)}))} : ((^~$signed((reg916 | wire898))) ?
                      $unsigned($signed($signed(reg921))) : reg905[(5'h12):(2'h3)]));
              reg923 <= $signed(((|$signed({reg904,
                  reg914,
                  reg912})) ~^ {$unsigned({(8'ha7)}),
                  (reg918 ? (reg917 || reg917) : $signed(reg917)),
                  $signed((^(8'h9c)))}));
              reg924 = (&$signed(((7'h57) >> $unsigned(reg919))));
            end
          else
            begin
              reg922 = (reg905[(5'h1b):(5'h18)] ?
                  (~^$signed(reg924)) : (wire898[(3'h4):(2'h2)] ^~ ((reg911 != ((7'h45) ?
                          reg916 : wire899)) ?
                      $unsigned((&(8'h9d))) : reg912[(5'h17):(4'h8)])));
              reg924 = $signed(((!$unsigned((^~wire900))) + reg913[(2'h2):(1'h0)]));
              reg925 = wire897[(3'h7):(1'h0)];
              reg926 = reg919;
              reg927 <= reg922;
              reg928 <= reg918[(5'h11):(3'h6)];
            end
          for (forvar929 = (1'h0); (forvar929 < (1'h1)); forvar929 = (forvar929 + (1'h1)))
            begin
              reg930 <= (~$unsigned(((~^(-reg922)) >= ((wire901 == wire899) ?
                  $unsigned(reg915) : (wire898 - reg911)))));
              reg931 <= ($signed($unsigned((reg910[(4'he):(1'h0)] << (|forvar929)))) ?
                  $unsigned(reg912[(5'h17):(2'h2)]) : ($signed((reg928[(4'hc):(4'hb)] ?
                          $unsigned(reg904) : wire900[(3'h7):(1'h1)])) ?
                      $signed(reg921[(5'h1c):(5'h16)]) : ((reg930[(1'h1):(1'h0)] >= (reg913 ?
                          reg926 : forvar929)) || $unsigned(((7'h48) ?
                          (8'hbd) : reg926)))));
              reg932 <= ((8'ha8) ^ reg926[(3'h4):(2'h2)]);
              reg933 = {(wire900 ? (^(!(reg913 ? reg919 : reg921))) : reg912),
                  reg925,
                  ({($unsigned(reg925) ?
                          (reg919 ? (8'ha4) : reg932) : {reg925, wire899}),
                      $signed($signed(reg919)),
                      ((reg911 ~^ reg912) && $signed(reg926))} <= ((^~(reg914 ?
                          reg926 : reg910)) ?
                      $signed(reg910[(1'h0):(1'h0)]) : $unsigned((reg912 ?
                          reg911 : reg927))))};
              reg934 = ((^reg933) ? (~&reg913) : $signed(reg925));
              reg935 = reg912[(4'he):(2'h2)];
            end
          if ({$signed(($unsigned(wire897) ?
                  ((7'h4e) ? (!reg914) : $signed(reg916)) : wire901))})
            begin
              reg936 <= (reg933 ?
                  $unsigned($signed(((reg927 << wire899) ?
                      reg926[(3'h5):(1'h1)] : $unsigned(reg918)))) : $signed((8'ha1)));
              reg937 <= ($unsigned({((^reg932) << wire897),
                  reg925[(4'h8):(3'h6)],
                  (!reg910[(5'h16):(5'h11)])}) + reg925[(5'h13):(5'h13)]);
              reg938 = reg918;
            end
          else
            begin
              reg938 = reg925;
              reg939 = reg931[(4'hc):(4'h9)];
              reg940 <= ((reg914 >> (-((forvar929 | reg920) ?
                  reg933 : ((7'h52) ^ (8'had))))) >>> wire901[(4'hd):(4'hd)]);
            end
        end
      else
        begin
          for (forvar910 = (1'h0); (forvar910 < (3'h4)); forvar910 = (forvar910 + (1'h1)))
            begin
              reg914 = reg940[(5'h10):(4'h8)];
              reg915 <= $unsigned(({{forvar929, reg922, $unsigned(reg902)},
                  (reg905[(5'h1c):(4'h9)] >= (reg932 * reg934))} + reg932));
            end
          if (((!reg923[(3'h4):(1'h0)]) - $unsigned($unsigned((7'h57)))))
            begin
              reg918 <= reg912;
              reg920 <= reg933;
              reg922 = reg902[(2'h3):(1'h1)];
              reg924 = reg920[(2'h2):(1'h0)];
              reg925 = reg910[(4'hb):(2'h2)];
              reg927 <= reg915[(1'h0):(1'h0)];
            end
          else
            begin
              reg916 = ($unsigned((({reg930, reg911} ^ $signed(reg923)) ?
                      $signed((reg933 ? (7'h44) : reg912)) : {{reg940,
                              reg936,
                              reg902}})) ?
                  (|reg928) : (&reg912[(4'h9):(3'h4)]));
              reg917 = (+((8'ha8) ?
                  {$signed(reg922[(5'h13):(4'ha)]),
                      ((reg904 ^ wire898) <<< reg911[(5'h16):(4'he)])} : (^~{(reg911 ?
                          reg919 : reg921)})));
            end
        end
      if ((reg923 ? reg918[(5'h14):(5'h11)] : (!reg915[(3'h5):(1'h0)])))
        begin
          if (reg921[(1'h1):(1'h0)])
            begin
              reg941 = (~^reg918[(4'he):(4'ha)]);
              reg942 = (8'hbc);
              reg943 <= {(reg924 ?
                      (^reg910[(5'h1b):(5'h13)]) : {($unsigned(reg924) ?
                              (reg902 ? reg923 : wire899) : (&reg919))}),
                  wire899,
                  (^~(|(~|(reg912 >>> forvar910))))};
              reg944 <= (reg910 ?
                  $signed({(reg913[(1'h1):(1'h1)] <<< $unsigned(forvar929))}) : $unsigned((^(~|(reg930 ?
                      reg924 : reg910)))));
              reg945 = $signed((^(({reg922, reg935, reg919} ?
                      reg916[(5'h10):(4'hd)] : wire897) ?
                  $signed($unsigned(wire898)) : wire897)));
              reg946 <= {((+wire898[(3'h7):(3'h6)]) ?
                      reg915 : (|(reg914 ? (8'h9f) : wire898[(4'hf):(4'h9)]))),
                  $unsigned((~&$signed($unsigned(wire899))))};
              reg947 = (reg913 > (reg913[(3'h5):(1'h0)] >> {reg938}));
            end
          else
            begin
              reg943 <= $signed(reg946[(3'h7):(3'h4)]);
              reg945 = ($signed((-(~|(~&reg941)))) ?
                  $signed(reg937[(4'ha):(3'h4)]) : $unsigned(reg919));
              reg947 = reg905;
              reg948 = ((^wire897) == (+($signed(((7'h4a) + reg934)) ?
                  reg912 : ((forvar910 >>> reg945) ?
                      {reg940, reg938} : $signed(reg934)))));
              reg949 <= ($signed((reg937[(5'h13):(5'h13)] ?
                  ((reg915 << reg931) ?
                      (reg930 ?
                          reg917 : reg942) : (~^reg943)) : wire900)) && (!$signed($unsigned((forvar910 >> reg927)))));
            end
          if (($unsigned($signed({((7'h40) == reg916), {reg944}})) ?
              {((reg945 + (7'h50)) > (reg925 ?
                      (8'ha3) : $signed(reg946)))} : (-reg920[(2'h2):(1'h1)])))
            begin
              reg950 = $unsigned(((forvar929 > ((-reg923) <<< (reg949 ?
                  (8'hb4) : (7'h55)))) <= (8'h9d)));
            end
          else
            begin
              reg951 <= $signed(reg950[(3'h4):(2'h3)]);
              reg952 <= (8'hbc);
              reg953 = {((((^reg915) ?
                      reg913[(3'h4):(2'h2)] : (reg933 >> reg905)) <= ($unsigned(reg936) ?
                      $unsigned(reg941) : $unsigned(reg923))) | reg928)};
              reg954 <= $signed((($unsigned((reg942 >>> reg951)) & {((8'had) ?
                          reg953 : reg952),
                      (reg915 > reg919)}) ?
                  ((^reg914[(3'h6):(3'h4)]) ?
                      $signed($unsigned((8'hb9))) : reg944) : $signed(reg949[(5'h10):(4'hf)])));
              reg955 = reg935;
            end
        end
      else
        begin
          for (forvar941 = (1'h0); (forvar941 < (1'h0)); forvar941 = (forvar941 + (1'h1)))
            begin
              reg942 = (~|$signed($unsigned($unsigned($signed(wire899)))));
              reg945 = $signed(reg917);
            end
          reg946 <= reg905[(1'h0):(1'h0)];
        end
      reg956 = reg923[(1'h0):(1'h0)];
    end
  assign wire957 = reg940;
  always
    @(posedge clk) begin
      reg958 = $unsigned($signed($signed(({reg911, reg902, reg927} ?
          (wire897 - reg923) : $signed(reg946)))));
      reg959 = $unsigned(reg949[(4'he):(4'hb)]);
      reg960 <= wire901;
      for (forvar961 = (1'h0); (forvar961 < (2'h3)); forvar961 = (forvar961 + (1'h1)))
        begin
          if ({$signed(wire901)})
            begin
              reg962 <= reg904;
              reg963 <= (7'h46);
            end
          else
            begin
              reg962 <= $unsigned({({$unsigned(reg949)} ?
                      reg928 : (|((7'h4e) == (7'h43)))),
                  reg949[(3'h7):(1'h1)]});
              reg963 <= (reg931[(5'h19):(5'h17)] < (^~($unsigned((-reg915)) >>> {(reg944 ?
                      wire900 : wire957),
                  (reg960 ^ (8'hab)),
                  (reg912 ? reg963 : reg960)})));
            end
          if ($unsigned(((&{(reg958 >= reg962), (reg921 != reg937)}) ?
              (7'h4c) : reg920[(2'h2):(2'h2)])))
            begin
              reg964 = wire897;
            end
          else
            begin
              reg965 <= {reg931[(5'h18):(5'h14)],
                  $signed($signed(reg913)),
                  (!(^(~(reg913 ~^ reg918))))};
              reg966 <= (^reg965);
            end
          reg967 = (~^reg965[(1'h0):(1'h0)]);
          reg968 <= $unsigned(reg930);
          for (forvar969 = (1'h0); (forvar969 < (3'h5)); forvar969 = (forvar969 + (1'h1)))
            begin
              reg970 = reg920;
              reg971 <= (({$unsigned((^reg902))} ?
                  reg968 : (!$unsigned(reg927[(3'h6):(3'h6)]))) && $unsigned(($unsigned($unsigned(forvar969)) ?
                  {(reg959 - reg954),
                      $signed((7'h4a)),
                      $unsigned((7'h4d))} : wire900[(4'hb):(3'h6)])));
              reg972 <= {reg932, forvar969};
              reg973 <= $signed($unsigned({(~$signed(reg932)),
                  ($unsigned(wire957) | reg964)}));
              reg974 = ((reg943 ?
                      ((^$unsigned(reg971)) == {(forvar961 >>> forvar969)}) : (~^reg920[(1'h1):(1'h0)])) ?
                  {reg973} : (&{reg959}));
            end
          reg975 <= (+reg959[(5'h12):(4'hb)]);
        end
    end
  assign wire976 = $signed((&($unsigned((reg937 < reg920)) ~^ reg966)));
  assign wire977 = $unsigned(wire900);
  assign wire978 = reg951;
  always
    @(posedge clk) begin
      if (reg972[(3'h4):(2'h3)])
        begin
          reg979 = (reg936[(2'h3):(1'h0)] ?
              $unsigned(reg915) : (reg911[(1'h0):(1'h0)] ?
                  reg918[(4'hc):(2'h2)] : $unsigned((^(&reg951)))));
          reg980 <= (&($signed({(^~reg920),
              $signed(reg944)}) >> (($signed(reg965) ^~ wire901) * reg972)));
          for (forvar981 = (1'h0); (forvar981 < (1'h1)); forvar981 = (forvar981 + (1'h1)))
            begin
              reg982 = $signed((+$signed({reg927[(5'h15):(1'h1)],
                  reg936[(4'hc):(1'h0)],
                  reg944[(4'h8):(2'h2)]})));
              reg983 <= ((~^reg930) <= ($unsigned($signed((reg944 != (7'h44)))) ?
                  ((reg936[(4'hc):(4'h9)] >>> reg965) ~^ wire977) : $unsigned({reg960})));
              reg984 <= $signed(((~&{$signed(reg973), (wire977 && reg960)}) ?
                  $unsigned((~&(reg930 ? (7'h43) : reg962))) : (^~((reg940 ?
                          reg943 : reg982) ?
                      $signed(reg971) : (reg975 && reg946)))));
              reg985 = ($unsigned((reg975[(3'h5):(3'h5)] - (reg951[(1'h1):(1'h1)] ?
                      (7'h44) : {wire977}))) ?
                  {wire899,
                      $signed((~&(+forvar981))),
                      reg923} : (~|($unsigned($signed(reg968)) >> $signed(reg920[(1'h1):(1'h1)]))));
              reg986 <= {reg940[(4'h8):(2'h3)], $unsigned($signed(reg905))};
            end
          if (($unsigned(wire899) + reg949))
            begin
              reg987 = (^reg946);
              reg988 <= ({(((|forvar981) ?
                          $unsigned(reg949) : reg954[(5'h15):(5'h10)]) | (!{reg944,
                          reg944})),
                      {$signed($unsigned(reg962))}} ?
                  {{(reg971 ? $unsigned((7'h4d)) : (^~reg972)),
                          reg937,
                          $unsigned(reg962[(4'he):(1'h0)])}} : $signed($unsigned({(reg984 ?
                          reg962 : reg962),
                      {reg936, reg963, (8'ha9)},
                      ((7'h4a) <= reg973)})));
              reg989 <= (~^$signed(reg983));
            end
          else
            begin
              reg988 <= (&$signed(reg930[(2'h2):(2'h2)]));
              reg990 = reg973[(3'h5):(1'h0)];
              reg991 <= reg987[(3'h5):(3'h5)];
              reg992 <= {reg927,
                  $signed($unsigned((reg973[(1'h0):(1'h0)] ?
                      (wire900 ? (7'h55) : reg985) : $unsigned((7'h4f)))))};
              reg993 <= reg940;
            end
          reg994 <= reg915[(1'h1):(1'h1)];
          reg995 <= reg927;
        end
      else
        begin
          for (forvar979 = (1'h0); (forvar979 < (1'h1)); forvar979 = (forvar979 + (1'h1)))
            begin
              reg981 = (({$unsigned(wire976),
                      $signed({reg949, forvar979, reg986}),
                      (-{reg988})} < (((reg944 >= reg937) << {(8'hbf),
                          reg989,
                          reg980}) ?
                      {reg972, reg979} : ($unsigned(reg912) * reg968))) ?
                  {(7'h50),
                      {$signed((reg991 >> wire901))},
                      $unsigned(($signed((7'h4a)) ?
                          ((8'ha3) ?
                              wire897 : (8'ha4)) : $signed(reg990)))} : wire978[(1'h0):(1'h0)]);
              reg982 = $unsigned({$unsigned(wire899[(3'h5):(1'h1)]),
                  reg944,
                  reg983});
            end
        end
      for (forvar996 = (1'h0); (forvar996 < (3'h6)); forvar996 = (forvar996 + (1'h1)))
        begin
          reg997 <= reg918[(4'ha):(2'h2)];
          reg998 <= wire897[(4'h9):(2'h3)];
          for (forvar999 = (1'h0); (forvar999 < (2'h3)); forvar999 = (forvar999 + (1'h1)))
            begin
              reg1000 <= $signed((8'ha6));
              reg1001 = $signed((~|(^~$unsigned(wire898))));
              reg1002 <= (forvar996 ?
                  (wire898[(4'ha):(3'h7)] >> reg932[(4'hd):(3'h4)]) : ((8'hbc) ?
                      $unsigned(($signed(reg991) & $signed(reg951))) : reg985[(2'h2):(1'h1)]));
              reg1003 = reg936;
            end
          reg1004 <= (-($unsigned($unsigned((reg931 ?
              reg993 : reg944))) >> (~^(-(~^(7'h48))))));
        end
    end
  module1005 #() modinst1406 (wire1405, clk, wire978, reg1004, reg928, reg946, reg915);
  assign wire1407 = ({(!{{reg944}}),
                        $signed(reg992),
                        reg937[(4'hf):(3'h7)]} > ((reg988 < (reg989 ?
                        reg973 : reg988)) << ((((8'hb7) * reg940) ?
                            reg937[(4'ha):(1'h0)] : ((8'hbc) ?
                                reg920 : reg954)) ?
                        {$unsigned(reg963)} : ($unsigned(reg986) ?
                            (reg936 ^ reg905) : reg965[(4'h8):(3'h6)]))));
  always
    @(posedge clk) begin
      reg1408 <= ((&$signed((8'hb4))) ?
          wire901[(1'h1):(1'h1)] : (~^reg902[(2'h3):(2'h3)]));
      reg1409 <= ($signed(reg972) ?
          ($signed($signed(reg989[(2'h2):(2'h2)])) ?
              reg960 : {(reg991[(4'hf):(4'hb)] * (reg928 ? (7'h54) : reg995)),
                  reg983,
                  (((7'h46) ? reg968 : (7'h55)) ?
                      $signed(reg963) : $unsigned(wire977))}) : $signed($signed((^reg915[(4'hb):(3'h4)]))));
      for (forvar1410 = (1'h0); (forvar1410 < (1'h0)); forvar1410 = (forvar1410 + (1'h1)))
        begin
          if ((($unsigned({reg949, $unsigned((8'hb4)), (reg965 <<< reg913)}) ?
              ($signed($unsigned((8'hb0))) <<< ((reg1004 > (8'hbf)) ?
                  {reg1004, (8'hb1)} : {reg931,
                      reg1409})) : (+(reg915 * ((7'h57) ?
                  reg937 : wire1407)))) >> ($signed(reg966) ?
              (reg966[(3'h6):(1'h1)] ?
                  {((8'ha1) * wire1407)} : $signed($signed(reg1004))) : $unsigned(reg989))))
            begin
              reg1411 <= ((forvar1410 ?
                      ({(reg1004 + reg960), {wire897}} ?
                          $unsigned(reg940) : (!wire901[(4'hc):(1'h0)])) : $signed((reg905[(4'h8):(1'h1)] ?
                          $unsigned(reg965) : $unsigned(reg915)))) ?
                  ($unsigned(reg972) >>> ((reg988 >>> {reg972}) >> (7'h43))) : $unsigned(reg920[(1'h0):(1'h0)]));
              reg1412 <= (~|(($signed(reg931[(3'h7):(3'h7)]) || (((8'h9e) >= reg997) >>> (reg954 ?
                      reg918 : reg975))) ?
                  reg966[(4'hb):(3'h6)] : $unsigned(((|reg1004) * reg920))));
              reg1413 = {$unsigned(((&{reg998, reg963, reg972}) ?
                      {(forvar1410 ? reg904 : reg937),
                          (reg988 ^~ reg918)} : $signed((reg943 >= wire957)))),
                  ($unsigned((~|reg913)) ?
                      $unsigned({$signed(reg998),
                          (reg931 ?
                              (8'hbb) : reg993)}) : $unsigned(($unsigned((7'h45)) ?
                          (reg943 - reg952) : (~reg983)))),
                  {(~^($signed(reg989) ? reg980[(1'h1):(1'h1)] : (^~(7'h42)))),
                      (^~$signed($unsigned(wire899))),
                      (($unsigned(reg920) ?
                          (!(8'ha8)) : ((7'h53) ?
                              reg968 : forvar1410)) || reg963[(5'h16):(5'h15)])}};
              reg1414 <= (7'h4d);
              reg1415 <= reg904;
              reg1416 = {({$unsigned((&(7'h43)))} && $signed((~(wire1405 ?
                      wire1405 : reg995))))};
            end
          else
            begin
              reg1413 = $unsigned((~^(reg991 ?
                  reg992[(3'h5):(1'h0)] : (reg1414 * reg915))));
              reg1416 = $unsigned($unsigned(reg983));
              reg1417 <= (^~(&$unsigned(reg921)));
              reg1418 <= reg972[(5'h14):(3'h4)];
            end
          for (forvar1419 = (1'h0); (forvar1419 < (2'h3)); forvar1419 = (forvar1419 + (1'h1)))
            begin
              reg1420 <= (wire1407[(4'ha):(4'h9)] ?
                  ($unsigned({wire1405,
                      $signed(reg1411),
                      reg975[(4'h9):(3'h6)]}) << $signed(($unsigned(wire901) << (8'hb2)))) : reg972);
              reg1421 = (($signed((&reg944)) >> (8'h9e)) <= $unsigned(($unsigned(reg980[(1'h0):(1'h0)]) >> $unsigned($signed(reg963)))));
            end
          reg1422 <= $signed(reg952[(4'hf):(4'hc)]);
          for (forvar1423 = (1'h0); (forvar1423 < (1'h0)); forvar1423 = (forvar1423 + (1'h1)))
            begin
              reg1424 = (reg989[(3'h6):(1'h1)] >>> (~|reg984[(5'h10):(4'hc)]));
              reg1425 = $signed({{reg986[(5'h12):(4'hf)]},
                  reg904[(3'h6):(3'h4)],
                  {($unsigned((7'h57)) ? $unsigned(wire977) : (|reg1417))}});
              reg1426 = {(reg988 ?
                      (!{(reg954 ? (7'h47) : reg1002),
                          reg904,
                          reg994}) : (~|reg992)),
                  reg927[(4'hc):(1'h1)],
                  {(wire978[(4'hb):(2'h2)] ?
                          ((reg984 != wire957) ?
                              {reg1416} : $unsigned(reg1422)) : $signed({wire897,
                              reg998,
                              (7'h41)})),
                      (($signed((8'ha1)) >> $signed(reg943)) ?
                          $signed(reg1412[(3'h5):(3'h4)]) : $signed($signed(reg968)))}};
              reg1427 <= {{{(reg997[(3'h7):(3'h5)] ?
                              forvar1423 : $signed(reg994)),
                          ($signed(reg991) ^~ $signed(reg971))},
                      (($unsigned(forvar1410) * reg936[(4'h8):(1'h0)]) ?
                          (8'hb0) : reg1004[(2'h2):(2'h2)])}};
            end
        end
      reg1428 = reg918[(5'h18):(5'h18)];
      if (reg991[(5'h17):(5'h10)])
        begin
          reg1429 = wire976[(3'h4):(1'h0)];
          if ((((reg1409 | reg1411[(3'h7):(1'h0)]) ?
              ((^~(^~reg1413)) ?
                  reg905[(4'hd):(2'h3)] : ($unsigned(forvar1423) != $unsigned(forvar1423))) : $signed(reg1408[(1'h0):(1'h0)])) >>> ({wire977} >> reg1429)))
            begin
              reg1430 = {($signed((reg928[(5'h10):(4'ha)] ?
                          (wire1407 ? reg1408 : reg973) : $signed(reg1413))) ?
                      (~|$signed($signed(reg980))) : (reg943[(5'h15):(5'h14)] ?
                          (reg920[(1'h0):(1'h0)] ?
                              (wire898 | reg913) : (reg940 ?
                                  wire899 : (8'hb6))) : {reg915,
                              reg1004[(2'h2):(1'h0)]}))};
              reg1431 = ({reg1002,
                      reg968[(1'h1):(1'h1)],
                      (reg931 & $unsigned($signed(reg994)))} ?
                  (($unsigned(reg1420[(4'hf):(4'hd)]) ?
                          wire1407[(4'he):(3'h5)] : {(reg905 ?
                                  reg975 : reg937)}) ?
                      reg920 : (8'ha1)) : reg983[(4'hf):(4'ha)]);
              reg1432 = (^~($signed(reg965) ?
                  ((^$unsigned(reg1428)) ^ forvar1423[(5'h11):(4'ha)]) : (~&((7'h56) ^~ (reg986 ?
                      reg973 : reg944)))));
              reg1433 <= reg988;
              reg1434 <= {((|(^(|reg913))) ?
                      $signed(reg1421[(2'h3):(2'h2)]) : reg971),
                  (~^(($unsigned(reg1002) ? reg940 : (&(8'had))) ?
                      (~^$unsigned(reg998)) : (7'h55)))};
            end
          else
            begin
              reg1433 <= $unsigned(wire977[(4'hb):(3'h5)]);
              reg1434 <= wire900[(4'h8):(2'h3)];
              reg1435 = (+(|(|reg962)));
              reg1436 <= reg972;
            end
          if (($signed(reg993[(4'ha):(4'ha)]) ?
              reg960[(5'h1a):(5'h1a)] : reg923[(1'h1):(1'h1)]))
            begin
              reg1437 = (reg904 ? $unsigned($signed((-(~|reg913)))) : reg989);
              reg1438 = (-(reg973[(4'h9):(3'h6)] ?
                  $signed(($signed(reg913) ~^ $unsigned(reg972))) : ($unsigned(((8'had) ?
                      reg960 : wire976)) | (reg1421 ?
                      reg1427 : ((8'hb9) >> reg995)))));
            end
          else
            begin
              reg1439 <= $signed((~|({(reg998 ? reg1424 : reg918)} ?
                  $signed((reg928 & reg1411)) : {reg993[(2'h3):(2'h2)],
                      forvar1423[(1'h1):(1'h1)],
                      (~^reg965)})));
            end
          reg1440 <= $signed(reg998);
        end
      else
        begin
          for (forvar1429 = (1'h0); (forvar1429 < (3'h4)); forvar1429 = (forvar1429 + (1'h1)))
            begin
              reg1433 <= reg1424;
              reg1435 = reg1411;
              reg1436 <= reg936[(4'hb):(1'h0)];
              reg1439 <= (reg921 ?
                  $unsigned({$signed((reg1002 || reg937)),
                      reg928[(4'hd):(4'hc)],
                      reg913}) : reg936[(4'hb):(4'h8)]);
              reg1440 <= ($unsigned((7'h44)) ?
                  (-reg1418) : (-{$signed({reg904, reg1429}),
                      reg915[(2'h3):(2'h3)]}));
              reg1441 <= ($unsigned(((~((8'ha4) ?
                      reg1429 : (7'h55))) * ($unsigned(reg943) || $signed(reg983)))) ?
                  (!$signed((reg943[(5'h11):(3'h5)] ^ reg1429[(1'h0):(1'h0)]))) : reg968);
              reg1442 <= reg1431[(5'h15):(4'hf)];
            end
          reg1443 <= (+((reg943[(5'h15):(5'h15)] >= reg1413[(3'h7):(2'h3)]) <<< reg1427[(1'h1):(1'h0)]));
          for (forvar1444 = (1'h0); (forvar1444 < (1'h1)); forvar1444 = (forvar1444 + (1'h1)))
            begin
              reg1445 <= reg1422[(4'he):(4'h8)];
              reg1446 <= (wire976 ?
                  (($unsigned(reg965[(2'h2):(1'h0)]) >= {reg997,
                          $signed(reg973)}) ?
                      $signed($signed(reg1441)) : reg1432[(5'h10):(3'h5)]) : {$unsigned($unsigned((reg921 | reg984))),
                      {((reg1428 ? reg931 : wire976) ?
                              $unsigned(reg940) : (reg931 ?
                                  forvar1410 : (7'h4d))),
                          ((reg988 && reg980) ?
                              $unsigned((8'hb1)) : (reg944 - reg975)),
                          {(|reg911), reg951[(4'hc):(3'h7)]}}});
            end
          for (forvar1447 = (1'h0); (forvar1447 < (3'h4)); forvar1447 = (forvar1447 + (1'h1)))
            begin
              reg1448 = (reg1413[(5'h11):(4'hd)] ? reg1434 : (|reg1439));
              reg1449 <= $signed((~^($signed(reg920[(1'h0):(1'h0)]) ?
                  reg927[(1'h0):(1'h0)] : reg1414[(2'h3):(1'h0)])));
              reg1450 <= ($unsigned(reg991[(3'h6):(1'h1)]) >= $signed({reg918[(4'h8):(2'h2)],
                  $signed((reg911 <<< (8'hb9))),
                  $unsigned((+reg944))}));
              reg1451 = reg995[(3'h5):(1'h1)];
              reg1452 = ((wire978[(3'h4):(2'h3)] ?
                  (|((8'hac) << (reg971 ?
                      reg1442 : reg1424))) : {(reg997 >= ((7'h41) ?
                          reg951 : reg962))}) >= (((~$unsigned(reg962)) ?
                  ((reg966 ? forvar1423 : reg991) & (8'hbf)) : {reg940,
                      $unsigned(reg1415),
                      reg944}) << $signed($unsigned(reg995))));
            end
          for (forvar1453 = (1'h0); (forvar1453 < (1'h1)); forvar1453 = (forvar1453 + (1'h1)))
            begin
              reg1454 = reg911[(4'he):(4'hb)];
              reg1455 <= ((~|({(~reg1417),
                      {reg1409, reg1413},
                      (~&reg1449)} << reg968)) ?
                  reg1414[(4'hc):(4'h8)] : wire957);
              reg1456 <= {(reg940[(3'h4):(1'h0)] ?
                      forvar1453 : $unsigned((forvar1444 ?
                          {reg1431, reg1432} : (+reg1426)))),
                  $unsigned(reg1448),
                  reg986[(5'h12):(3'h4)]};
              reg1457 = (($signed({$unsigned(reg913),
                  (8'ha6)}) ^~ reg1426[(2'h3):(1'h1)]) <= (|reg1426));
              reg1458 = (({(reg1002[(4'hc):(4'h8)] << (reg1450 >> wire900)),
                      (-(reg1455 < reg1450))} ?
                  (8'hbe) : ({(reg1457 ? reg962 : reg1456)} ?
                      ((reg1438 ? reg1449 : reg931) >> (reg975 ?
                          reg1427 : (7'h4f))) : reg1409)) << reg983[(4'ha):(4'h9)]);
            end
          for (forvar1459 = (1'h0); (forvar1459 < (1'h1)); forvar1459 = (forvar1459 + (1'h1)))
            begin
              reg1460 = ($signed($signed($signed((&forvar1453)))) != $signed($signed(((~^reg936) ?
                  reg1455 : {reg1421, reg1436}))));
              reg1461 = (-$signed(($unsigned(reg1445[(2'h3):(2'h3)]) ?
                  reg1451[(1'h1):(1'h0)] : reg1433[(3'h5):(2'h3)])));
              reg1462 = reg992[(4'h8):(2'h2)];
              reg1463 <= $unsigned(wire899);
              reg1464 = forvar1459;
            end
          if ($signed((^~{(+(~^reg1463))})))
            begin
              reg1465 <= {reg994, reg943[(3'h7):(1'h0)]};
              reg1466 <= $unsigned(reg923[(2'h2):(1'h1)]);
              reg1467 <= reg984;
              reg1468 <= ((reg991[(4'hd):(1'h1)] == {($signed((8'ha2)) ?
                      (~^reg905) : $unsigned(reg1450)),
                  {{reg1451, reg1438},
                      reg1409[(4'h8):(2'h2)],
                      (wire978 ?
                          reg920 : reg911)}}) >> $signed(wire976[(3'h6):(2'h3)]));
              reg1469 <= reg1415;
              reg1470 = reg1456[(2'h2):(2'h2)];
              reg1471 = ((reg944 ?
                  ((!reg1469[(4'hb):(2'h2)]) ?
                      (reg1417[(4'h8):(1'h0)] <= forvar1453[(4'he):(4'h8)]) : $signed(((8'ha3) <<< (8'ha8)))) : (~^(!(^reg902)))) & reg1442);
            end
          else
            begin
              reg1470 = reg918;
              reg1472 <= ((!reg954[(3'h7):(3'h5)]) ?
                  (!$unsigned(reg1461)) : {$unsigned(reg965)});
              reg1473 = ($unsigned((((reg1461 ? wire978 : reg921) ?
                          $signed((8'hb3)) : (forvar1429 ? reg1463 : reg928)) ?
                      (^(forvar1410 <= forvar1410)) : $signed(reg932[(3'h6):(1'h0)]))) ?
                  $signed(forvar1447[(5'h10):(1'h0)]) : (reg975[(4'h9):(3'h6)] ?
                      {(+(reg1418 ?
                              reg946 : reg1431))} : $unsigned(((reg1439 ~^ reg1408) || $signed(reg1004)))));
              reg1474 = $unsigned({reg1466[(3'h7):(2'h2)]});
            end
        end
      reg1475 <= (reg1442 ? forvar1410[(5'h15):(5'h10)] : wire897);
      if (({$unsigned((~|(~|reg944))),
          (^$unsigned($unsigned((7'h43))))} ^ forvar1447[(5'h10):(5'h10)]))
        begin
          reg1476 <= reg1467;
          reg1477 <= {reg1430,
              {forvar1429[(4'h8):(4'h8)],
                  ({$signed(reg1411),
                      (reg1421 <= wire977),
                      (forvar1423 >> forvar1419)} * reg1467[(1'h0):(1'h0)]),
                  forvar1423},
              $signed(({(8'hae)} ?
                  (reg1472 ?
                      $unsigned(reg1435) : ((7'h4b) + wire900)) : forvar1429[(1'h0):(1'h0)]))};
          if ($signed(reg991))
            begin
              reg1478 = $signed(((-$unsigned($signed(forvar1410))) && reg960));
            end
          else
            begin
              reg1479 <= (+reg1472[(3'h6):(1'h0)]);
              reg1480 <= $signed(({$unsigned((7'h51))} == (!reg1470)));
            end
          reg1481 = ({$unsigned(reg904[(4'h8):(3'h6)])} ?
              ($unsigned(reg986[(5'h10):(4'h9)]) & reg1461[(1'h1):(1'h1)]) : ((8'hbe) + reg1417));
          reg1482 <= {$unsigned($unsigned((reg1433 ?
                  (reg1470 ? reg1422 : (8'hbe)) : (|wire898)))),
              $signed((~^$signed($unsigned(wire900)))),
              $unsigned((wire900[(3'h4):(2'h2)] ?
                  $signed(reg995[(3'h5):(3'h5)]) : {$signed(wire901)}))};
          reg1483 <= $signed(((forvar1447[(5'h18):(3'h6)] ?
              (+(~&reg1432)) : reg1439) <<< (reg930[(2'h2):(1'h0)] ?
              reg1463[(4'h9):(3'h6)] : ((~|reg1413) ?
                  (forvar1423 ? reg962 : reg1440) : $signed(reg927)))));
          if ((reg932[(1'h0):(1'h0)] ?
              $signed((~reg932[(4'ha):(3'h4)])) : wire977[(4'hf):(4'hd)]))
            begin
              reg1484 <= (reg997 ?
                  {$unsigned(reg1475[(3'h7):(3'h4)]),
                      ((&(~reg1448)) + ($signed(reg1440) != $signed((8'ha4)))),
                      reg989[(3'h5):(1'h0)]} : $unsigned($unsigned(reg998)));
              reg1485 = forvar1459[(3'h4):(1'h0)];
              reg1486 <= ((~|{forvar1423,
                      (reg989 == $signed(reg1440)),
                      (~&$signed(reg1434))}) ?
                  reg1481 : (reg1477 > $signed($unsigned((reg984 != reg1450)))));
            end
          else
            begin
              reg1485 = reg1416;
              reg1487 = ((-forvar1419) ?
                  $unsigned(($unsigned(reg1417) ?
                      reg1430[(5'h10):(5'h10)] : ((reg1443 ? (8'ha7) : reg936) ?
                          (8'ha4) : $signed((7'h47))))) : $unsigned(reg988));
              reg1488 = (forvar1447 ?
                  (~|reg1479[(1'h1):(1'h1)]) : reg1485[(3'h5):(2'h3)]);
            end
        end
      else
        begin
          if ({(-reg1433[(2'h3):(1'h1)]),
              forvar1444[(2'h3):(2'h2)],
              (reg1424[(1'h1):(1'h1)] ?
                  reg1441[(1'h1):(1'h1)] : (|((reg940 ? reg1002 : reg1427) ?
                      {wire900, reg1434, forvar1459} : (reg1004 ^~ (8'ha5)))))})
            begin
              reg1476 <= reg946;
              reg1477 <= {$signed({reg992, $unsigned(reg1428)}),
                  $signed($signed((&$signed(forvar1453)))),
                  {reg905}};
              reg1478 = $signed((($unsigned((reg913 <<< reg962)) ?
                      (reg1461 ?
                          $signed(reg968) : $unsigned(wire957)) : $unsigned((8'hac))) ?
                  (forvar1423[(3'h6):(2'h2)] >= (-(reg904 >= reg1470))) : $signed(reg1428[(5'h15):(5'h14)])));
            end
          else
            begin
              reg1476 <= $unsigned((~|(^~$signed((&(7'h52))))));
              reg1478 = reg937[(1'h0):(1'h0)];
              reg1479 <= $signed(((reg952 ?
                  $signed($signed(reg1464)) : ({reg937,
                      forvar1447} != $signed(reg1429))) & (reg1471[(4'hb):(4'h8)] ?
                  (8'ha1) : (reg1463[(2'h2):(1'h0)] ?
                      (reg918 == (7'h4a)) : (reg973 != wire977)))));
              reg1481 = {(reg1442 >= $signed((((7'h4f) != (7'h45)) & reg980))),
                  (^~reg1441),
                  $signed($signed(reg1477[(4'he):(3'h4)]))};
            end
          for (forvar1482 = (1'h0); (forvar1482 < (2'h3)); forvar1482 = (forvar1482 + (1'h1)))
            begin
              reg1485 = $unsigned((!($signed({reg989,
                  reg918}) >>> $unsigned((+reg936)))));
              reg1487 = reg968;
              reg1489 <= (reg1483 >= ($unsigned((!$unsigned(reg927))) ?
                  $signed((~|$signed((8'hb2)))) : ((reg1455 ?
                          {forvar1410} : (forvar1419 ? reg1477 : (8'hb9))) ?
                      reg1440 : reg1457[(3'h6):(3'h5)])));
              reg1490 <= $signed((~^reg963));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module517
#(parameter param582 = {(((-((8'hac) ? (8'hbc) : (7'h45))) || {((7'h49) + (7'h52)), {(7'h49), (8'hb3), (8'ha6)}}) * ((&(~(8'had))) <= (|((7'h58) & (7'h4b))))), ((!(((8'hba) - (7'h50)) && {(8'hb9), (8'h9e)})) ^ (~|((~|(8'hb9)) <<< (+(8'hb3)))))}, 
parameter param583 = (param582 <<< (param582 ? param582 : (((^param582) ? (param582 | param582) : param582) ? ((param582 ~^ param582) << (param582 << param582)) : (((7'h54) ^ param582) ? (~^param582) : (-param582))))))
(y, clk, wire521, wire520, wire519, wire518);
  output wire [(32'h341):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire521;
  input wire [(5'h18):(1'h0)] wire520;
  input wire [(5'h1a):(1'h0)] wire519;
  input wire [(4'hd):(1'h0)] wire518;
  wire [(3'h5):(1'h0)] wire581;
  wire [(4'ha):(1'h0)] wire580;
  wire [(5'h11):(1'h0)] wire523;
  reg signed [(4'h8):(1'h0)] reg579 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg578 = (1'h0);
  reg [(4'h8):(1'h0)] reg577 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg575 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg574 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg572 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg571 = (1'h0);
  reg [(5'h13):(1'h0)] reg567 = (1'h0);
  reg [(5'h10):(1'h0)] reg564 = (1'h0);
  reg [(5'h1a):(1'h0)] reg556 = (1'h0);
  reg [(5'h11):(1'h0)] reg551 = (1'h0);
  reg [(4'he):(1'h0)] reg550 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg548 = (1'h0);
  reg [(5'h1e):(1'h0)] reg547 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg545 = (1'h0);
  reg [(4'hc):(1'h0)] reg543 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg538 = (1'h0);
  reg [(5'h18):(1'h0)] reg533 = (1'h0);
  reg [(5'h1c):(1'h0)] reg531 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg530 = (1'h0);
  reg [(5'h1e):(1'h0)] reg529 = (1'h0);
  reg [(4'hd):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg526 = (1'h0);
  reg [(5'h1c):(1'h0)] reg524 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg576 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar573 = (1'h0);
  reg [(3'h5):(1'h0)] reg570 = (1'h0);
  reg [(5'h13):(1'h0)] reg569 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg568 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg566 = (1'h0);
  reg [(5'h15):(1'h0)] reg565 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg561 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg562 = (1'h0);
  reg [(3'h5):(1'h0)] forvar561 = (1'h0);
  reg [(4'he):(1'h0)] reg560 = (1'h0);
  reg [(5'h16):(1'h0)] reg559 = (1'h0);
  reg [(3'h4):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg557 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg555 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg554 = (1'h0);
  reg [(4'ha):(1'h0)] reg553 = (1'h0);
  reg [(2'h2):(1'h0)] reg552 = (1'h0);
  reg [(4'ha):(1'h0)] reg549 = (1'h0);
  reg [(2'h3):(1'h0)] reg546 = (1'h0);
  reg [(4'h9):(1'h0)] reg544 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar542 = (1'h0);
  reg [(5'h1b):(1'h0)] reg541 = (1'h0);
  reg [(5'h1a):(1'h0)] reg540 = (1'h0);
  reg [(4'h8):(1'h0)] forvar539 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg537 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg536 = (1'h0);
  reg [(2'h3):(1'h0)] reg535 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar534 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg527 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg525 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg522 = (1'h0);
  assign y = {wire581,
                 wire580,
                 wire523,
                 reg579,
                 reg578,
                 reg577,
                 reg575,
                 reg574,
                 reg572,
                 reg571,
                 reg567,
                 reg564,
                 reg556,
                 reg551,
                 reg550,
                 reg548,
                 reg547,
                 reg545,
                 reg543,
                 reg538,
                 reg533,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg526,
                 reg524,
                 reg576,
                 forvar573,
                 reg570,
                 reg569,
                 reg568,
                 reg566,
                 reg565,
                 reg561,
                 reg563,
                 reg562,
                 forvar561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg549,
                 reg546,
                 reg544,
                 forvar542,
                 reg541,
                 reg540,
                 forvar539,
                 reg537,
                 reg536,
                 reg535,
                 forvar534,
                 reg532,
                 reg527,
                 reg525,
                 reg522,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg522 = ($unsigned(($signed(wire519[(5'h13):(4'hf)]) ?
          (~^$signed(wire520)) : ((~wire518) >>> $unsigned(wire521)))) << (wire520[(5'h18):(4'hb)] >> wire519[(5'h14):(2'h2)]));
    end
  assign wire523 = $signed((wire520[(1'h1):(1'h1)] ?
                       $unsigned($signed($unsigned(wire520))) : $signed($unsigned(wire519))));
  always
    @(posedge clk) begin
      if ((!$unsigned(wire519)))
        begin
          reg524 <= wire523[(4'hb):(4'h8)];
        end
      else
        begin
          reg525 = (wire520 ?
              ($signed(({wire523, wire519} ?
                  {(7'h4e),
                      reg524} : (7'h45))) >> (($signed(wire521) | wire520) <= (7'h41))) : wire518);
          reg526 <= wire523;
          reg527 = wire520;
          reg528 <= (~^($unsigned(($unsigned((8'hba)) << reg526)) - ((^(wire519 ?
                  wire520 : (7'h4a))) ?
              ($signed(wire518) ?
                  reg525 : wire518[(3'h4):(2'h2)]) : $signed({wire523,
                  (8'hb8),
                  wire523}))));
          if (wire521[(5'h13):(4'hb)])
            begin
              reg529 <= (reg528 ?
                  reg524[(3'h4):(1'h1)] : $signed({($unsigned(reg525) + (reg526 ?
                          reg526 : reg526))}));
              reg530 <= ($signed($unsigned(((reg529 ^~ wire521) ?
                  (|wire521) : reg527))) | (wire521 ?
                  {$signed((7'h49)), reg527[(4'hf):(2'h3)]} : (((reg527 ?
                      reg527 : reg526) << (wire521 ^ wire523)) <= (reg526[(3'h4):(2'h3)] ?
                      reg529[(5'h17):(1'h1)] : (wire521 >= wire519)))));
              reg531 <= wire523;
              reg532 = reg531;
              reg533 <= $unsigned($signed(reg532[(1'h0):(1'h0)]));
            end
          else
            begin
              reg532 = (-wire519);
            end
          for (forvar534 = (1'h0); (forvar534 < (3'h4)); forvar534 = (forvar534 + (1'h1)))
            begin
              reg535 = (7'h43);
              reg536 = {(($unsigned((reg533 ? (7'h54) : reg524)) << (^(reg527 ?
                          reg524 : reg529))) ?
                      reg526[(4'ha):(2'h2)] : ($signed({reg527,
                          (8'hb7)}) - $signed((8'h9d))))};
              reg537 = (-({$signed(((8'haf) ? reg527 : reg530)),
                  ({wire520, reg524, forvar534} ?
                      $signed((7'h4d)) : (wire518 ?
                          reg526 : (7'h4c)))} <= {$unsigned(reg530),
                  reg531,
                  $signed($unsigned(reg532))}));
            end
        end
      reg538 <= forvar534;
      for (forvar539 = (1'h0); (forvar539 < (3'h6)); forvar539 = (forvar539 + (1'h1)))
        begin
          reg540 = ($signed((!$signed((8'h9f)))) ?
              $signed((8'hb7)) : (reg527[(5'h16):(4'he)] ?
                  reg530[(1'h1):(1'h0)] : ((reg525[(3'h6):(1'h0)] << (wire521 ?
                          wire518 : reg537)) ?
                      {reg532[(2'h3):(1'h0)],
                          wire519[(2'h2):(2'h2)]} : ($unsigned(reg524) ?
                          $signed(reg524) : $signed(reg530)))));
          reg541 = $signed((8'hae));
          for (forvar542 = (1'h0); (forvar542 < (3'h5)); forvar542 = (forvar542 + (1'h1)))
            begin
              reg543 <= $unsigned($signed($unsigned($signed((-reg532)))));
              reg544 = $unsigned(((+$signed((wire520 ? reg525 : reg541))) ?
                  ((!$unsigned(reg535)) >>> (~&reg538[(2'h3):(1'h1)])) : reg538[(1'h0):(1'h0)]));
              reg545 <= (~$unsigned((&($unsigned(forvar539) < (reg524 ?
                  reg541 : (8'haf))))));
              reg546 = $signed($unsigned(({((8'h9e) ? forvar539 : reg533),
                  reg525,
                  (8'hb0)} * (~$unsigned((7'h53))))));
              reg547 <= (7'h57);
              reg548 <= $unsigned(((7'h52) ?
                  reg529[(5'h12):(4'h8)] : $signed($unsigned((forvar542 <= forvar539)))));
            end
          reg549 = reg530[(2'h3):(1'h1)];
          reg550 <= $unsigned((7'h53));
          reg551 <= ((&$unsigned(({reg543} ^~ {(7'h47)}))) <<< reg532[(1'h0):(1'h0)]);
          if ((-(reg529[(5'h14):(3'h6)] ?
              (|reg524[(4'hc):(1'h0)]) : $signed(reg546[(2'h3):(1'h0)]))))
            begin
              reg552 = wire519;
              reg553 = (&($signed(({reg540, forvar534, forvar542} <= ((7'h55) ?
                  reg529 : reg536))) >> reg543));
              reg554 = $unsigned(($unsigned($signed({reg528, reg529})) ?
                  {((reg544 && reg535) ?
                          (reg528 ?
                              (7'h45) : reg525) : $signed(reg546))} : (~^(reg533[(3'h4):(2'h3)] > (+(8'ha0))))));
              reg555 = ($unsigned($unsigned($unsigned(forvar542))) != ((reg543[(4'hb):(3'h4)] == (+(8'hb4))) <<< (&(^$unsigned(reg554)))));
            end
          else
            begin
              reg552 = (~&($signed(((~wire523) ?
                  (reg546 >> wire519) : $signed((7'h48)))) == (($unsigned((7'h43)) ?
                  (reg526 || reg541) : {wire519,
                      reg533}) >= $signed($signed(reg540)))));
              reg556 <= $unsigned(reg541[(5'h17):(3'h6)]);
              reg557 = ($signed((&((!forvar542) > wire518))) ?
                  (forvar542[(4'ha):(2'h3)] ?
                      (reg525 ?
                          $signed((reg546 ? reg531 : (8'ha6))) : ((reg555 ?
                              reg550 : reg535) <= $signed((8'hb1)))) : reg528) : $signed(($signed($unsigned(reg545)) - reg544[(3'h6):(3'h5)])));
              reg558 = ((-$signed({(wire518 ? reg525 : reg531),
                  $signed(reg556)})) < {$unsigned((~&{reg544,
                      reg556,
                      reg527}))});
            end
        end
      if ({reg528[(4'ha):(4'h9)], forvar534[(3'h5):(2'h2)], $unsigned((7'h51))})
        begin
          reg559 = (^~(forvar534 ?
              {$unsigned((reg554 ?
                      reg524 : reg549))} : {(wire520[(4'hd):(2'h2)] ?
                      {wire523, reg526} : ((7'h54) >>> reg546)),
                  (^~$unsigned((8'hbe)))}));
          reg560 = reg543[(3'h7):(3'h4)];
          for (forvar561 = (1'h0); (forvar561 < (2'h3)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 = {$unsigned((({reg545, wire523, reg552} ?
                      $unsigned(wire518) : reg547[(5'h1a):(5'h13)]) == $unsigned(reg535))),
                  reg535};
            end
          reg563 = (^reg524[(1'h0):(1'h0)]);
        end
      else
        begin
          reg559 = reg525[(1'h0):(1'h0)];
          if ((&{$unsigned((~(&reg559)))}))
            begin
              reg560 = $unsigned(((reg548[(1'h0):(1'h0)] ?
                  ($unsigned(reg552) ?
                      ((8'hbe) && reg553) : forvar542[(3'h4):(1'h1)]) : ($unsigned(reg551) <= (!wire520))) || (reg531 ?
                  forvar534 : wire521)));
              reg561 = (^$signed($unsigned(reg528)));
              reg564 <= $unsigned($unsigned(reg526[(4'hb):(2'h2)]));
              reg565 = wire523;
              reg566 = ((-(|(!reg556))) ?
                  (~^$signed((+$signed(reg560)))) : reg553);
              reg567 <= reg545[(5'h1b):(3'h4)];
            end
          else
            begin
              reg564 <= (((reg525[(2'h2):(2'h2)] ?
                      reg524[(3'h7):(3'h7)] : {(^reg547),
                          forvar561}) ^~ (!((reg533 ?
                      reg566 : (8'ha4)) < reg545))) ?
                  $signed($signed(reg564)) : $unsigned(((^~reg560) ~^ reg558[(3'h4):(2'h3)])));
              reg565 = reg544;
              reg566 = {({$signed((&reg551)),
                          $signed(((8'h9c) ? reg541 : reg546))} ?
                      $signed((reg550 > $unsigned(reg558))) : reg555),
                  {($unsigned((reg532 ?
                          reg540 : (7'h56))) ^ (~|$unsigned((8'haa)))),
                      (reg547 <<< reg537[(3'h4):(1'h0)])}};
              reg568 = $signed(reg531);
              reg569 = (~&reg528[(4'hb):(2'h3)]);
              reg570 = $signed(($signed((reg524 ?
                      $signed(reg567) : $unsigned(reg552))) ?
                  ($unsigned($unsigned(reg565)) >>> wire523) : $unsigned(forvar561)));
              reg571 <= reg535;
            end
          reg572 <= $unsigned(($signed($unsigned({(7'h40),
              (8'hb9)})) * ($signed($unsigned(reg546)) ?
              $signed({wire518}) : ((reg535 >>> (7'h47)) > (reg567 ?
                  reg553 : wire518)))));
          for (forvar573 = (1'h0); (forvar573 < (3'h4)); forvar573 = (forvar573 + (1'h1)))
            begin
              reg574 <= (7'h4d);
              reg575 <= reg553;
              reg576 = wire518[(2'h2):(1'h1)];
            end
          reg577 <= (^~{reg538});
          reg578 <= reg576;
        end
      reg579 <= ((wire520 ?
              (((reg578 ? wire518 : reg552) == (reg557 ^~ (8'ha9))) ?
                  {reg558,
                      wire521[(4'h9):(4'h9)],
                      $unsigned(reg558)} : ((reg574 << (8'h9d)) ?
                      $signed(reg559) : reg544[(3'h7):(1'h1)])) : reg556[(4'he):(4'hd)]) ?
          ($signed({{reg553, reg557}}) ?
              (~((reg554 ? reg533 : reg545) ?
                  wire520[(4'h8):(3'h4)] : $unsigned(reg526))) : reg531[(3'h7):(2'h3)]) : reg544[(4'h8):(1'h1)]);
    end
  assign wire580 = {((~|$signed($unsigned(reg529))) | ($unsigned(reg538) ?
                           (-{reg543,
                               reg524,
                               wire520}) : $signed(reg526[(5'h12):(4'hc)]))),
                       (^$unsigned(reg547[(3'h5):(1'h0)]))};
  assign wire581 = (wire521[(5'h10):(4'hb)] | $unsigned($unsigned($signed($unsigned(reg575)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1005
#(parameter param1403 = {{(~^(((8'ha5) ? (7'h56) : (7'h43)) ? ((8'h9d) ? (8'hb3) : (7'h4e)) : {(7'h4c), (8'hb3)})), ((+(&(8'hb1))) <<< ((~&(7'h45)) ? (-(8'haf)) : ((8'hb9) ? (8'ha7) : (8'ha4))))}}, 
parameter param1404 = {((&((^~(8'hbf)) <<< (param1403 & param1403))) || (((^param1403) - (param1403 ? param1403 : param1403)) && param1403))})
(y, clk, wire1010, wire1009, wire1008, wire1007, wire1006);
  output wire [(32'h199b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire1010;
  input wire [(4'h9):(1'h0)] wire1009;
  input wire [(5'h1f):(1'h0)] wire1008;
  input wire [(2'h2):(1'h0)] wire1007;
  input wire signed [(5'h1a):(1'h0)] wire1006;
  wire signed [(3'h5):(1'h0)] wire1364;
  wire signed [(5'h12):(1'h0)] wire1231;
  wire [(5'h17):(1'h0)] wire1230;
  wire [(4'h9):(1'h0)] wire1229;
  wire [(5'h1d):(1'h0)] wire1228;
  wire signed [(5'h1a):(1'h0)] wire1226;
  wire [(5'h10):(1'h0)] wire1082;
  reg [(5'h15):(1'h0)] reg1402 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1401 = (1'h0);
  reg [(4'hc):(1'h0)] reg1400 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1395 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1365 = (1'h0);
  reg [(4'he):(1'h0)] reg1390 = (1'h0);
  reg [(5'h15):(1'h0)] reg1388 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1386 = (1'h0);
  reg [(2'h2):(1'h0)] reg1382 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1381 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1380 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1375 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1373 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1372 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1370 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1368 = (1'h0);
  reg [(5'h14):(1'h0)] reg1367 = (1'h0);
  reg [(4'hc):(1'h0)] reg1366 = (1'h0);
  reg [(5'h10):(1'h0)] reg1363 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1352 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1361 = (1'h0);
  reg [(2'h2):(1'h0)] reg1360 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1359 = (1'h0);
  reg [(5'h10):(1'h0)] reg1358 = (1'h0);
  reg [(4'h9):(1'h0)] reg1357 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1355 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1344 = (1'h0);
  reg [(4'ha):(1'h0)] reg1342 = (1'h0);
  reg [(4'hc):(1'h0)] reg1339 = (1'h0);
  reg [(5'h11):(1'h0)] reg1338 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1336 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1335 = (1'h0);
  reg [(5'h14):(1'h0)] reg1334 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1332 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1324 = (1'h0);
  reg [(3'h7):(1'h0)] reg1323 = (1'h0);
  reg [(5'h18):(1'h0)] reg1322 = (1'h0);
  reg [(4'hb):(1'h0)] reg1321 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1318 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1315 = (1'h0);
  reg [(5'h16):(1'h0)] reg1314 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1313 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1309 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1308 = (1'h0);
  reg [(5'h17):(1'h0)] reg1307 = (1'h0);
  reg [(4'hf):(1'h0)] reg1302 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1301 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1298 = (1'h0);
  reg [(4'ha):(1'h0)] reg1293 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1292 = (1'h0);
  reg [(4'h9):(1'h0)] reg1291 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1289 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1286 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1281 = (1'h0);
  reg [(5'h15):(1'h0)] reg1280 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1279 = (1'h0);
  reg [(5'h16):(1'h0)] reg1277 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1276 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1272 = (1'h0);
  reg [(5'h18):(1'h0)] reg1269 = (1'h0);
  reg [(5'h13):(1'h0)] reg1268 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1267 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1266 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1263 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1262 = (1'h0);
  reg [(2'h3):(1'h0)] reg1259 = (1'h0);
  reg [(5'h10):(1'h0)] reg1258 = (1'h0);
  reg [(4'ha):(1'h0)] reg1254 = (1'h0);
  reg [(4'h8):(1'h0)] reg1251 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1246 = (1'h0);
  reg [(3'h5):(1'h0)] reg1245 = (1'h0);
  reg [(5'h18):(1'h0)] reg1241 = (1'h0);
  reg [(3'h6):(1'h0)] reg1238 = (1'h0);
  reg [(4'ha):(1'h0)] reg1237 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1236 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1235 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1227 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1225 = (1'h0);
  reg [(5'h13):(1'h0)] reg1204 = (1'h0);
  reg [(5'h15):(1'h0)] reg1196 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1222 = (1'h0);
  reg [(3'h6):(1'h0)] reg1221 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1219 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1218 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1216 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1208 = (1'h0);
  reg [(4'h8):(1'h0)] reg1207 = (1'h0);
  reg [(5'h18):(1'h0)] reg1206 = (1'h0);
  reg [(2'h3):(1'h0)] reg1203 = (1'h0);
  reg [(4'hd):(1'h0)] reg1198 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1197 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1194 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1193 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1192 = (1'h0);
  reg [(5'h13):(1'h0)] reg1191 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1189 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1188 = (1'h0);
  reg [(4'hf):(1'h0)] reg1187 = (1'h0);
  reg [(4'he):(1'h0)] reg1175 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1184 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1183 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1179 = (1'h0);
  reg [(5'h15):(1'h0)] reg1177 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1172 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1170 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1167 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1165 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1161 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1159 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1158 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1156 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1155 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1152 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1151 = (1'h0);
  reg [(5'h15):(1'h0)] reg1149 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1148 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1146 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1145 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1144 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1142 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1139 = (1'h0);
  reg [(5'h12):(1'h0)] reg1138 = (1'h0);
  reg [(4'hb):(1'h0)] reg1136 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1133 = (1'h0);
  reg [(4'hb):(1'h0)] reg1132 = (1'h0);
  reg [(4'h8):(1'h0)] reg1130 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1127 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1126 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1124 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1122 = (1'h0);
  reg [(4'h8):(1'h0)] reg1121 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1118 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1117 = (1'h0);
  reg [(2'h3):(1'h0)] reg1112 = (1'h0);
  reg [(5'h14):(1'h0)] reg1106 = (1'h0);
  reg [(2'h3):(1'h0)] reg1102 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1101 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1100 = (1'h0);
  reg [(3'h7):(1'h0)] reg1099 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1094 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1093 = (1'h0);
  reg [(4'he):(1'h0)] reg1092 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1089 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1088 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1087 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1086 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1085 = (1'h0);
  reg [(4'h9):(1'h0)] reg1078 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1077 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1076 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1074 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1071 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1070 = (1'h0);
  reg [(4'ha):(1'h0)] reg1066 = (1'h0);
  reg [(5'h12):(1'h0)] reg1056 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1055 = (1'h0);
  reg [(4'hc):(1'h0)] reg1053 = (1'h0);
  reg [(4'h8):(1'h0)] reg1052 = (1'h0);
  reg [(4'hb):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1049 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1048 = (1'h0);
  reg [(5'h16):(1'h0)] reg1041 = (1'h0);
  reg [(3'h7):(1'h0)] reg1038 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1043 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1042 = (1'h0);
  reg [(2'h2):(1'h0)] reg1030 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1035 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1034 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1033 = (1'h0);
  reg [(5'h17):(1'h0)] reg1032 = (1'h0);
  reg [(4'h9):(1'h0)] reg1027 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1025 = (1'h0);
  reg [(5'h11):(1'h0)] reg1024 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1016 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1015 = (1'h0);
  reg [(5'h11):(1'h0)] reg1013 = (1'h0);
  reg [(5'h11):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1011 = (1'h0);
  reg [(5'h16):(1'h0)] reg1399 = (1'h0);
  reg [(5'h11):(1'h0)] reg1398 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1397 = (1'h0);
  reg [(2'h2):(1'h0)] reg1396 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1394 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1393 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1366 = (1'h0);
  reg [(3'h6):(1'h0)] reg1392 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1391 = (1'h0);
  reg [(5'h15):(1'h0)] reg1389 = (1'h0);
  reg [(2'h3):(1'h0)] reg1387 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1385 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1383 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1379 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1378 = (1'h0);
  reg [(5'h14):(1'h0)] reg1377 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1376 = (1'h0);
  reg [(3'h5):(1'h0)] reg1374 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1371 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1369 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1365 = (1'h0);
  reg [(4'hb):(1'h0)] reg1362 = (1'h0);
  reg [(3'h7):(1'h0)] reg1354 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1343 = (1'h0);
  reg [(2'h3):(1'h0)] reg1356 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1354 = (1'h0);
  reg [(3'h4):(1'h0)] reg1353 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1352 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1351 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1350 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1349 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1348 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1347 = (1'h0);
  reg [(4'h9):(1'h0)] reg1346 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1345 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar1343 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1341 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1340 = (1'h0);
  reg [(4'h8):(1'h0)] reg1337 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1333 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1331 = (1'h0);
  reg [(4'he):(1'h0)] reg1330 = (1'h0);
  reg [(5'h16):(1'h0)] reg1329 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1328 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1327 = (1'h0);
  reg [(5'h18):(1'h0)] reg1326 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1325 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1320 = (1'h0);
  reg [(4'h8):(1'h0)] reg1319 = (1'h0);
  reg [(4'ha):(1'h0)] reg1317 = (1'h0);
  reg [(3'h7):(1'h0)] reg1316 = (1'h0);
  reg [(4'hb):(1'h0)] reg1312 = (1'h0);
  reg [(4'hb):(1'h0)] reg1311 = (1'h0);
  reg [(4'h8):(1'h0)] reg1310 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1306 = (1'h0);
  reg [(3'h4):(1'h0)] reg1305 = (1'h0);
  reg [(3'h6):(1'h0)] reg1304 = (1'h0);
  reg [(3'h5):(1'h0)] reg1303 = (1'h0);
  reg [(5'h10):(1'h0)] reg1300 = (1'h0);
  reg [(3'h7):(1'h0)] reg1299 = (1'h0);
  reg [(5'h18):(1'h0)] reg1297 = (1'h0);
  reg [(4'hb):(1'h0)] reg1296 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1295 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1294 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1290 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1288 = (1'h0);
  reg [(4'hc):(1'h0)] reg1287 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1285 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1284 = (1'h0);
  reg [(5'h10):(1'h0)] reg1283 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1282 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1278 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1275 = (1'h0);
  reg [(4'he):(1'h0)] reg1274 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1273 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1271 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1270 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1265 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1264 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1261 = (1'h0);
  reg [(3'h6):(1'h0)] reg1260 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1257 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar1256 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1255 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1253 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1252 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1250 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1249 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1248 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1247 = (1'h0);
  reg [(4'hb):(1'h0)] reg1244 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1243 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1242 = (1'h0);
  reg [(5'h10):(1'h0)] reg1240 = (1'h0);
  reg [(5'h16):(1'h0)] reg1239 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1234 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1233 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1232 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1224 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1200 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1190 = (1'h0);
  reg [(5'h15):(1'h0)] reg1223 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1220 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1217 = (1'h0);
  reg [(2'h2):(1'h0)] reg1215 = (1'h0);
  reg [(4'hb):(1'h0)] reg1214 = (1'h0);
  reg [(3'h5):(1'h0)] reg1213 = (1'h0);
  reg [(3'h7):(1'h0)] reg1212 = (1'h0);
  reg [(5'h13):(1'h0)] reg1211 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1210 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1209 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1205 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1204 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1202 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1201 = (1'h0);
  reg [(4'hf):(1'h0)] reg1200 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1199 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1196 = (1'h0);
  reg [(4'h8):(1'h0)] reg1195 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1190 = (1'h0);
  reg [(5'h12):(1'h0)] reg1186 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1185 = (1'h0);
  reg [(4'hf):(1'h0)] reg1182 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1181 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1180 = (1'h0);
  reg [(5'h12):(1'h0)] reg1178 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1175 = (1'h0);
  reg [(4'h9):(1'h0)] reg1174 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1173 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1171 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1169 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1168 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1166 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1164 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1163 = (1'h0);
  reg [(4'hd):(1'h0)] reg1162 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1160 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1157 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1154 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1148 = (1'h0);
  reg [(5'h12):(1'h0)] reg1153 = (1'h0);
  reg [(5'h17):(1'h0)] reg1150 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1147 = (1'h0);
  reg [(5'h17):(1'h0)] reg1143 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1125 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1122 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1115 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1141 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1140 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1137 = (1'h0);
  reg [(3'h6):(1'h0)] reg1135 = (1'h0);
  reg [(5'h17):(1'h0)] reg1134 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1131 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1129 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1128 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar1125 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1123 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1120 = (1'h0);
  reg [(5'h18):(1'h0)] reg1119 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1116 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1115 = (1'h0);
  reg [(5'h15):(1'h0)] reg1114 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1113 = (1'h0);
  reg [(5'h11):(1'h0)] reg1111 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1110 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1109 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1108 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1107 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1105 = (1'h0);
  reg [(5'h14):(1'h0)] reg1104 = (1'h0);
  reg [(4'hb):(1'h0)] reg1103 = (1'h0);
  reg [(5'h12):(1'h0)] reg1098 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1097 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1095 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1091 = (1'h0);
  reg [(5'h11):(1'h0)] reg1090 = (1'h0);
  reg [(4'hd):(1'h0)] reg1084 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1083 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1081 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1080 = (1'h0);
  reg [(5'h15):(1'h0)] reg1079 = (1'h0);
  reg [(4'h8):(1'h0)] reg1075 = (1'h0);
  reg [(4'hf):(1'h0)] reg1073 = (1'h0);
  reg [(4'ha):(1'h0)] reg1072 = (1'h0);
  reg [(5'h11):(1'h0)] reg1069 = (1'h0);
  reg [(3'h6):(1'h0)] reg1068 = (1'h0);
  reg [(2'h2):(1'h0)] reg1067 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1065 = (1'h0);
  reg [(3'h7):(1'h0)] reg1064 = (1'h0);
  reg [(2'h3):(1'h0)] reg1063 = (1'h0);
  reg [(5'h19):(1'h0)] reg1062 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1061 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1060 = (1'h0);
  reg [(2'h2):(1'h0)] reg1059 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1058 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1057 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1054 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1051 = (1'h0);
  reg [(3'h6):(1'h0)] reg1047 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1046 = (1'h0);
  reg [(2'h3):(1'h0)] reg1045 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1044 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1039 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1041 = (1'h0);
  reg [(5'h14):(1'h0)] reg1040 = (1'h0);
  reg [(4'hc):(1'h0)] reg1039 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1038 = (1'h0);
  reg [(5'h14):(1'h0)] reg1037 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1036 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar1029 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1026 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1012 = (1'h0);
  reg [(2'h3):(1'h0)] reg1031 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1030 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1029 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1028 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1026 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1023 = (1'h0);
  reg [(2'h3):(1'h0)] reg1022 = (1'h0);
  reg [(5'h19):(1'h0)] reg1021 = (1'h0);
  reg [(5'h15):(1'h0)] reg1020 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1019 = (1'h0);
  reg [(5'h12):(1'h0)] reg1018 = (1'h0);
  reg [(5'h13):(1'h0)] reg1017 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1014 = (1'h0);
  assign y = {wire1364,
                 wire1231,
                 wire1230,
                 wire1229,
                 wire1228,
                 wire1226,
                 wire1082,
                 reg1402,
                 reg1401,
                 reg1400,
                 reg1395,
                 reg1365,
                 reg1390,
                 reg1388,
                 reg1386,
                 reg1382,
                 reg1381,
                 reg1380,
                 reg1375,
                 reg1373,
                 reg1372,
                 reg1370,
                 reg1368,
                 reg1367,
                 reg1366,
                 reg1363,
                 reg1352,
                 reg1361,
                 reg1360,
                 reg1359,
                 reg1358,
                 reg1357,
                 reg1355,
                 reg1344,
                 reg1342,
                 reg1339,
                 reg1338,
                 reg1336,
                 reg1335,
                 reg1334,
                 reg1332,
                 reg1324,
                 reg1323,
                 reg1322,
                 reg1321,
                 reg1318,
                 reg1315,
                 reg1314,
                 reg1313,
                 reg1309,
                 reg1308,
                 reg1307,
                 reg1302,
                 reg1301,
                 reg1298,
                 reg1293,
                 reg1292,
                 reg1291,
                 reg1289,
                 reg1286,
                 reg1281,
                 reg1280,
                 reg1279,
                 reg1277,
                 reg1276,
                 reg1272,
                 reg1269,
                 reg1268,
                 reg1267,
                 reg1266,
                 reg1263,
                 reg1262,
                 reg1259,
                 reg1258,
                 reg1254,
                 reg1251,
                 reg1246,
                 reg1245,
                 reg1241,
                 reg1238,
                 reg1237,
                 reg1236,
                 reg1235,
                 reg1227,
                 reg1225,
                 reg1204,
                 reg1196,
                 reg1222,
                 reg1221,
                 reg1219,
                 reg1218,
                 reg1216,
                 reg1208,
                 reg1207,
                 reg1206,
                 reg1203,
                 reg1198,
                 reg1197,
                 reg1194,
                 reg1193,
                 reg1192,
                 reg1191,
                 reg1189,
                 reg1188,
                 reg1187,
                 reg1175,
                 reg1184,
                 reg1183,
                 reg1179,
                 reg1177,
                 reg1172,
                 reg1170,
                 reg1167,
                 reg1165,
                 reg1161,
                 reg1159,
                 reg1158,
                 reg1156,
                 reg1155,
                 reg1152,
                 reg1151,
                 reg1149,
                 reg1148,
                 reg1146,
                 reg1145,
                 reg1144,
                 reg1142,
                 reg1139,
                 reg1138,
                 reg1136,
                 reg1133,
                 reg1132,
                 reg1130,
                 reg1127,
                 reg1126,
                 reg1124,
                 reg1122,
                 reg1121,
                 reg1118,
                 reg1117,
                 reg1112,
                 reg1106,
                 reg1102,
                 reg1101,
                 reg1100,
                 reg1099,
                 reg1096,
                 reg1094,
                 reg1093,
                 reg1092,
                 reg1089,
                 reg1088,
                 reg1087,
                 reg1086,
                 reg1085,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1074,
                 reg1071,
                 reg1070,
                 reg1066,
                 reg1056,
                 reg1055,
                 reg1053,
                 reg1052,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1041,
                 reg1038,
                 reg1043,
                 reg1042,
                 reg1030,
                 reg1035,
                 reg1034,
                 reg1033,
                 reg1032,
                 reg1027,
                 reg1025,
                 reg1024,
                 reg1016,
                 reg1015,
                 reg1013,
                 reg1012,
                 reg1011,
                 reg1399,
                 reg1398,
                 forvar1397,
                 reg1396,
                 forvar1394,
                 forvar1393,
                 forvar1366,
                 reg1392,
                 reg1391,
                 reg1389,
                 reg1387,
                 reg1385,
                 forvar1384,
                 reg1383,
                 reg1379,
                 reg1378,
                 reg1377,
                 reg1376,
                 reg1374,
                 reg1371,
                 reg1369,
                 forvar1365,
                 reg1362,
                 reg1354,
                 reg1343,
                 reg1356,
                 forvar1354,
                 reg1353,
                 forvar1352,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1348,
                 reg1347,
                 reg1346,
                 reg1345,
                 forvar1343,
                 reg1341,
                 reg1340,
                 reg1337,
                 reg1333,
                 reg1331,
                 reg1330,
                 reg1329,
                 reg1328,
                 reg1327,
                 reg1326,
                 reg1325,
                 reg1320,
                 reg1319,
                 reg1317,
                 reg1316,
                 reg1312,
                 reg1311,
                 reg1310,
                 reg1306,
                 reg1305,
                 reg1304,
                 reg1303,
                 reg1300,
                 reg1299,
                 reg1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 reg1290,
                 reg1288,
                 reg1287,
                 reg1285,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1278,
                 reg1275,
                 reg1274,
                 reg1273,
                 forvar1271,
                 forvar1270,
                 forvar1265,
                 reg1264,
                 reg1261,
                 reg1260,
                 forvar1257,
                 forvar1256,
                 reg1255,
                 reg1253,
                 forvar1252,
                 reg1250,
                 reg1249,
                 reg1248,
                 reg1247,
                 reg1244,
                 forvar1243,
                 reg1242,
                 reg1240,
                 reg1239,
                 reg1234,
                 reg1233,
                 forvar1232,
                 reg1224,
                 forvar1200,
                 forvar1190,
                 reg1223,
                 reg1220,
                 reg1217,
                 reg1215,
                 reg1214,
                 reg1213,
                 reg1212,
                 reg1211,
                 reg1210,
                 reg1209,
                 reg1205,
                 forvar1204,
                 reg1202,
                 reg1201,
                 reg1200,
                 reg1199,
                 forvar1196,
                 reg1195,
                 reg1190,
                 reg1186,
                 reg1185,
                 reg1182,
                 reg1181,
                 reg1180,
                 reg1178,
                 reg1176,
                 forvar1175,
                 reg1174,
                 reg1173,
                 reg1171,
                 forvar1169,
                 reg1168,
                 reg1166,
                 reg1164,
                 reg1163,
                 reg1162,
                 reg1160,
                 reg1157,
                 reg1154,
                 forvar1148,
                 reg1153,
                 reg1150,
                 reg1147,
                 reg1143,
                 reg1125,
                 forvar1122,
                 forvar1115,
                 forvar1141,
                 reg1140,
                 reg1137,
                 reg1135,
                 reg1134,
                 forvar1131,
                 reg1129,
                 reg1128,
                 forvar1125,
                 reg1123,
                 reg1120,
                 reg1119,
                 reg1116,
                 reg1115,
                 reg1114,
                 reg1113,
                 reg1111,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1107,
                 reg1105,
                 reg1104,
                 reg1103,
                 reg1098,
                 reg1097,
                 reg1095,
                 reg1091,
                 reg1090,
                 reg1084,
                 forvar1083,
                 reg1081,
                 reg1080,
                 reg1079,
                 reg1075,
                 reg1073,
                 reg1072,
                 reg1069,
                 reg1068,
                 reg1067,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 reg1057,
                 reg1054,
                 reg1051,
                 reg1047,
                 reg1046,
                 reg1045,
                 reg1044,
                 forvar1039,
                 forvar1041,
                 reg1040,
                 reg1039,
                 forvar1038,
                 reg1037,
                 reg1036,
                 forvar1029,
                 reg1026,
                 forvar1012,
                 reg1031,
                 forvar1030,
                 reg1029,
                 reg1028,
                 forvar1026,
                 reg1023,
                 reg1022,
                 reg1021,
                 reg1020,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1014,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1011 <= $signed((wire1007 ?
          wire1008 : (!($unsigned(wire1008) ?
              wire1006 : (wire1008 >>> wire1007)))));
      if ($signed(wire1010))
        begin
          if (wire1010[(1'h0):(1'h0)])
            begin
              reg1012 <= $signed(wire1008[(4'h9):(1'h0)]);
              reg1013 <= $signed(($unsigned(reg1011) >= {$signed($signed(wire1006)),
                  wire1010[(2'h3):(1'h1)],
                  (^$signed(wire1009))}));
            end
          else
            begin
              reg1012 <= ($unsigned($signed(((wire1009 ? reg1012 : wire1008) ?
                  wire1007 : wire1006))) && (&wire1006));
              reg1013 <= (^~reg1011[(5'h11):(4'h9)]);
              reg1014 = wire1010[(4'ha):(3'h4)];
            end
          if (wire1007[(1'h1):(1'h0)])
            begin
              reg1015 <= (((wire1007[(1'h1):(1'h0)] ?
                  (+$signed(wire1009)) : ($unsigned(reg1011) ?
                      (~|reg1014) : wire1010[(3'h4):(2'h3)])) > {(~^(~|reg1014)),
                  $signed($unsigned(wire1007))}) >= $signed((reg1013 ?
                  (((8'hae) ? wire1007 : wire1008) ?
                      wire1010[(4'h9):(1'h0)] : (^~wire1007)) : reg1011[(5'h11):(4'ha)])));
              reg1016 <= (|(wire1007[(1'h0):(1'h0)] ?
                  $signed($signed(wire1009)) : (-{$unsigned(reg1012)})));
              reg1017 = ($unsigned(($signed(reg1013) ?
                      (8'hac) : {{wire1006, reg1016}, $signed(reg1015)})) ?
                  $signed(((reg1013[(4'hb):(3'h7)] ?
                      (!(7'h52)) : $unsigned(reg1013)) ^~ (+reg1015))) : $unsigned(((~|$unsigned(wire1010)) ?
                      $signed((^~wire1007)) : reg1012)));
              reg1018 = $signed(wire1009[(3'h6):(3'h5)]);
              reg1019 = $unsigned($signed(($unsigned(reg1014) ?
                  ($signed(reg1018) ?
                      reg1017 : {wire1009, reg1011, reg1016}) : ((reg1011 ?
                          wire1010 : wire1009) ?
                      (reg1016 ?
                          wire1007 : reg1017) : reg1012[(3'h6):(3'h6)]))));
              reg1020 = $signed((~(($unsigned(wire1006) * (reg1011 != reg1014)) ^ wire1009[(3'h4):(1'h0)])));
              reg1021 = (!reg1012[(4'h9):(1'h1)]);
            end
          else
            begin
              reg1017 = $unsigned($signed({reg1019[(4'hc):(2'h2)]}));
              reg1018 = $unsigned(({$unsigned(reg1017)} ?
                  wire1010[(3'h4):(3'h4)] : (wire1010 ?
                      (reg1020 ?
                          $signed((7'h47)) : wire1007) : reg1019[(5'h10):(4'he)])));
            end
          reg1022 = {(&(-(|(wire1006 ? reg1015 : (8'hb4))))),
              $unsigned(reg1011[(5'h11):(3'h4)]),
              {((reg1011[(4'hc):(3'h7)] > $signed(wire1007)) ?
                      ($unsigned((8'h9f)) <<< ((8'haa) <= (8'ha5))) : wire1007[(1'h1):(1'h1)])}};
          if ((reg1018[(4'hf):(3'h4)] ?
              $unsigned($unsigned(reg1020)) : $unsigned(reg1014[(5'h10):(4'ha)])))
            begin
              reg1023 = {(($unsigned(((7'h46) + reg1021)) ?
                          ($signed(wire1006) >>> (8'had)) : reg1018) ?
                      ($unsigned($unsigned(reg1013)) ?
                          reg1017 : {reg1022,
                              {reg1020, reg1018}}) : wire1010[(4'h8):(3'h4)]),
                  (~reg1021[(3'h6):(2'h3)])};
            end
          else
            begin
              reg1024 <= $unsigned(((~&$unsigned((reg1016 != reg1020))) <<< $unsigned(reg1019)));
              reg1025 <= $signed($unsigned(reg1020));
            end
          for (forvar1026 = (1'h0); (forvar1026 < (2'h2)); forvar1026 = (forvar1026 + (1'h1)))
            begin
              reg1027 <= reg1018[(3'h4):(2'h2)];
              reg1028 = reg1013[(3'h6):(1'h0)];
              reg1029 = (wire1007[(1'h1):(1'h1)] ?
                  reg1027[(3'h6):(3'h6)] : (($unsigned($signed(reg1020)) <<< (((7'h41) || reg1012) ?
                          $unsigned(wire1010) : ((7'h46) >> reg1013))) ?
                      (((reg1015 ? wire1010 : (8'hbe)) ?
                          reg1011[(4'he):(4'h9)] : wire1006) | $signed($signed(reg1020))) : wire1008));
            end
          for (forvar1030 = (1'h0); (forvar1030 < (1'h1)); forvar1030 = (forvar1030 + (1'h1)))
            begin
              reg1031 = forvar1030;
              reg1032 <= $signed(reg1027[(3'h6):(2'h3)]);
              reg1033 <= $signed({$signed($signed(reg1013[(2'h3):(1'h0)])),
                  ((7'h44) ^~ reg1018)});
              reg1034 <= {$signed(reg1018), $signed(wire1010), reg1020};
            end
          reg1035 <= forvar1026[(2'h2):(2'h2)];
        end
      else
        begin
          for (forvar1012 = (1'h0); (forvar1012 < (1'h1)); forvar1012 = (forvar1012 + (1'h1)))
            begin
              reg1013 <= $unsigned((forvar1012 & reg1011[(4'hb):(3'h7)]));
              reg1014 = (|$signed($unsigned($signed(reg1020[(5'h12):(4'ha)]))));
              reg1015 <= $unsigned($unsigned($unsigned({$signed(reg1019),
                  {(7'h44)},
                  {reg1035, (8'hac)}})));
              reg1017 = reg1021;
              reg1024 <= ({(((wire1009 ? reg1028 : wire1009) ?
                          $signed((7'h4b)) : reg1020[(4'h8):(3'h6)]) ^~ $unsigned($unsigned((8'ha3)))),
                      (^~(reg1027 ? reg1017[(1'h0):(1'h0)] : (+(7'h53)))),
                      $signed($unsigned($signed(wire1006)))} ?
                  (8'hb7) : ($unsigned(reg1024) ?
                      $signed(reg1031) : ((7'h51) ?
                          reg1012[(4'he):(1'h1)] : reg1032[(5'h10):(4'hf)])));
              reg1026 = ($unsigned(wire1009) + {$signed((~^reg1014[(4'h8):(3'h4)])),
                  $unsigned(((reg1031 ? reg1022 : reg1015) ?
                      (7'h55) : $signed(reg1022)))});
              reg1028 = (reg1015 ?
                  (!(((reg1013 ^~ reg1012) ? reg1018 : (8'ha0)) ?
                      ((forvar1012 ^ reg1034) ?
                          reg1013[(3'h4):(2'h3)] : (reg1019 ?
                              reg1013 : forvar1012)) : ({reg1033,
                              wire1008,
                              wire1010} ?
                          (+reg1021) : (reg1027 && reg1017)))) : reg1012[(4'hb):(4'h9)]);
            end
          for (forvar1029 = (1'h0); (forvar1029 < (3'h5)); forvar1029 = (forvar1029 + (1'h1)))
            begin
              reg1030 <= reg1029;
            end
        end
      if (($unsigned($unsigned($signed(reg1032[(1'h1):(1'h0)]))) ?
          reg1019 : $unsigned({reg1014[(5'h12):(5'h11)]})))
        begin
          reg1036 = (|($unsigned(wire1008[(5'h1c):(5'h12)]) ?
              reg1012 : reg1028[(4'hd):(3'h7)]));
          reg1037 = ((reg1025[(3'h6):(1'h1)] ?
              $signed($unsigned({(7'h48)})) : $signed(({(8'hb2)} ?
                  (~|forvar1026) : (reg1014 >= reg1012)))) * reg1023);
          for (forvar1038 = (1'h0); (forvar1038 < (1'h0)); forvar1038 = (forvar1038 + (1'h1)))
            begin
              reg1039 = ($signed(reg1031[(2'h2):(1'h1)]) || wire1006[(5'h11):(1'h0)]);
              reg1040 = {(~&(^~$signed($signed(forvar1030))))};
            end
          for (forvar1041 = (1'h0); (forvar1041 < (3'h6)); forvar1041 = (forvar1041 + (1'h1)))
            begin
              reg1042 <= forvar1038;
              reg1043 <= $unsigned(wire1010[(2'h2):(1'h1)]);
            end
        end
      else
        begin
          reg1038 <= $unsigned(reg1022);
          for (forvar1039 = (1'h0); (forvar1039 < (3'h6)); forvar1039 = (forvar1039 + (1'h1)))
            begin
              reg1041 <= (^~(|(7'h44)));
              reg1044 = (((~reg1040[(4'h9):(3'h4)]) ?
                  (wire1007 ?
                      {(^~reg1030), $signed(reg1019)} : {(forvar1012 ?
                              wire1007 : reg1027),
                          reg1038}) : reg1042[(2'h2):(2'h2)]) <<< (^reg1041));
              reg1045 = (+$signed($signed($signed((reg1030 ?
                  reg1020 : wire1007)))));
              reg1046 = {(~&($signed($unsigned(reg1027)) ?
                      (!(reg1033 ? reg1018 : forvar1012)) : (+reg1029)))};
            end
          if ((8'hb6))
            begin
              reg1047 = $unsigned(reg1028[(3'h6):(1'h1)]);
              reg1048 <= reg1030[(1'h0):(1'h0)];
              reg1049 <= reg1018;
              reg1050 <= $signed({$signed($signed($unsigned(reg1048)))});
              reg1051 = (~^$unsigned((8'hb9)));
              reg1052 <= wire1007[(1'h1):(1'h0)];
            end
          else
            begin
              reg1048 <= {(7'h4a)};
              reg1049 <= (forvar1030[(4'h9):(1'h1)] ?
                  ($unsigned({(reg1028 * reg1032)}) ?
                      $unsigned((|$signed((7'h58)))) : reg1026) : (8'hbb));
              reg1051 = (forvar1038[(2'h3):(1'h0)] ?
                  reg1034[(3'h4):(2'h3)] : (~&(~{$signed(reg1051),
                      $unsigned(forvar1041),
                      (reg1028 ? reg1020 : reg1046)})));
              reg1052 <= reg1052;
              reg1053 <= reg1048[(1'h1):(1'h1)];
              reg1054 = {reg1028,
                  (reg1013 ?
                      (~&((|reg1013) ?
                          (forvar1041 ^ (8'hb6)) : $unsigned(reg1030))) : ((~&$unsigned(forvar1026)) ?
                          $signed(reg1017[(2'h2):(1'h1)]) : $unsigned(reg1034))),
                  reg1053[(4'hc):(3'h4)]};
              reg1055 <= ($signed((~&reg1034[(3'h5):(2'h2)])) << ((&$signed(reg1035)) ?
                  ($signed($signed(reg1037)) ?
                      reg1023[(5'h10):(4'hc)] : ($unsigned(reg1042) < $signed(reg1027))) : (~&$unsigned($signed((7'h4a))))));
            end
        end
      reg1056 <= $unsigned(($signed((8'h9d)) && $unsigned((reg1015[(5'h18):(5'h18)] ?
          (+reg1045) : $signed((8'hbc))))));
      if ((reg1020[(4'hf):(1'h1)] ? reg1021 : $unsigned(reg1023)))
        begin
          reg1057 = ({({$unsigned(forvar1026)} ?
                  (reg1012[(4'ha):(3'h7)] >> (reg1011 ?
                      reg1045 : reg1041)) : (^~(7'h4a))),
              (~&$unsigned((&reg1052)))} * {$signed(reg1053),
              {reg1026[(5'h14):(3'h5)], $unsigned({(8'hb4)})}});
          if (($signed(($unsigned((reg1053 && reg1033)) >> reg1019[(4'hd):(3'h4)])) ?
              (~&(~^reg1039[(4'hb):(2'h3)])) : {$signed(reg1021),
                  $unsigned({$signed(reg1012), (reg1014 ^ reg1012)})}))
            begin
              reg1058 = $unsigned(reg1047);
            end
          else
            begin
              reg1058 = ($unsigned(reg1018) ^~ $signed(($signed(forvar1026) ?
                  $unsigned(((8'ha5) ?
                      (7'h41) : reg1012)) : $signed($signed(reg1036)))));
              reg1059 = (|$unsigned(($unsigned((reg1024 - reg1051)) <= reg1036[(2'h2):(2'h2)])));
              reg1060 = reg1026[(5'h10):(2'h3)];
              reg1061 = reg1039[(3'h4):(1'h0)];
              reg1062 = {wire1010, reg1037[(5'h11):(4'hf)]};
              reg1063 = forvar1030;
            end
          reg1064 = $unsigned(reg1046);
          reg1065 = reg1022;
          reg1066 <= reg1054[(1'h1):(1'h0)];
          if ({wire1010[(2'h3):(2'h3)],
              reg1056[(3'h4):(1'h0)],
              $signed((reg1019[(4'hc):(2'h3)] == reg1063))})
            begin
              reg1067 = $signed(($signed((^(&reg1042))) >>> (reg1064 > $unsigned(forvar1041[(1'h0):(1'h0)]))));
              reg1068 = reg1029[(3'h7):(3'h5)];
              reg1069 = ($unsigned({((~&reg1041) ?
                      (reg1039 + wire1006) : (reg1056 ?
                          reg1057 : (7'h41)))}) << $signed((reg1019[(2'h2):(1'h0)] - reg1038)));
              reg1070 <= $signed((^{((reg1031 ? reg1068 : reg1058) & (wire1006 ?
                      reg1065 : (7'h47))),
                  $unsigned($unsigned((7'h54)))}));
              reg1071 <= ((!(reg1011 >>> {(reg1055 > (8'ha4)),
                      $signed(reg1051)})) ?
                  (-(reg1022 * reg1048)) : (reg1049 != $signed($signed(reg1027))));
            end
          else
            begin
              reg1067 = $unsigned(forvar1026[(2'h2):(1'h0)]);
              reg1070 <= reg1032;
            end
          if ((|((|(7'h4b)) ?
              $signed(($unsigned(reg1043) + wire1009[(3'h7):(3'h6)])) : (reg1027[(4'h9):(3'h6)] ~^ $unsigned((reg1027 ^~ forvar1041))))))
            begin
              reg1072 = (~|reg1024);
              reg1073 = ((($signed((reg1044 ? reg1062 : reg1038)) ?
                          reg1031[(1'h0):(1'h0)] : ((reg1012 ~^ reg1050) | (reg1028 > wire1009))) ?
                      reg1038[(1'h1):(1'h0)] : ($unsigned($signed(forvar1039)) ^ (reg1027[(4'h9):(4'h8)] ?
                          {(8'ha0), reg1021} : (^reg1060)))) ?
                  (-(~^(~|(reg1032 ? reg1050 : reg1072)))) : (+(reg1031 ?
                      $signed((&reg1070)) : wire1008)));
            end
          else
            begin
              reg1074 <= $unsigned($signed((reg1015[(5'h1f):(5'h1e)] ?
                  (~&(~&reg1031)) : reg1062[(1'h1):(1'h0)])));
              reg1075 = (7'h55);
              reg1076 <= $unsigned($unsigned((reg1055 >= (reg1072 ^ $unsigned(reg1038)))));
              reg1077 <= (^($signed(reg1031) ^ reg1012[(4'hc):(3'h5)]));
              reg1078 <= wire1010[(3'h4):(3'h4)];
            end
        end
      else
        begin
          reg1066 <= ((^~($signed(((8'ha4) ? forvar1026 : reg1026)) ?
              (~reg1048) : $signed($signed(forvar1041)))) >= $unsigned((((&reg1023) > $signed((8'ha7))) > $signed(reg1051[(1'h0):(1'h0)]))));
          if ($unsigned(reg1020[(5'h10):(4'h9)]))
            begin
              reg1070 <= (($unsigned($signed((~forvar1038))) <= (~&($signed((7'h56)) & ((8'hb9) ?
                  (8'ha4) : reg1047)))) ^ $unsigned((((8'hb0) >= $signed(reg1061)) ?
                  $signed(wire1008[(1'h0):(1'h0)]) : $signed(reg1023))));
              reg1071 <= $unsigned(reg1042);
              reg1074 <= $signed($unsigned((reg1034 ?
                  (((8'hb6) || reg1071) >= $signed(forvar1041)) : ((7'h42) ?
                      forvar1012 : ((8'hb9) ? reg1021 : reg1036)))));
              reg1076 <= $unsigned($unsigned(reg1048));
              reg1079 = $unsigned($signed((&(reg1016 ~^ (reg1076 <= reg1068)))));
            end
          else
            begin
              reg1070 <= {$unsigned(reg1057)};
              reg1072 = $signed((reg1050[(4'hb):(2'h3)] ~^ reg1066));
              reg1073 = ($unsigned($unsigned(reg1011[(3'h5):(2'h2)])) ?
                  {reg1053[(3'h7):(3'h4)]} : $signed((^($signed(reg1012) || (reg1029 <<< reg1070)))));
              reg1074 <= (|($signed(reg1069[(5'h10):(4'hf)]) ?
                  reg1075 : reg1052));
              reg1076 <= (~$signed(((~&reg1053) ? (~^(~reg1016)) : (7'h55))));
            end
          reg1080 = {(7'h51),
              reg1059[(1'h1):(1'h0)],
              $signed({$unsigned(reg1023), reg1032[(5'h14):(4'ha)]})};
          reg1081 = (8'hbf);
        end
    end
  assign wire1082 = reg1042[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar1083 = (1'h0); (forvar1083 < (1'h1)); forvar1083 = (forvar1083 + (1'h1)))
        begin
          reg1084 = ({$signed((|(reg1042 ? wire1009 : (7'h42))))} ?
              reg1052 : $signed((!$signed({reg1011, reg1070, reg1012}))));
          reg1085 <= {(+$signed(((~^(8'hbe)) ?
                  reg1084[(3'h7):(1'h1)] : $signed(reg1084)))),
              reg1070[(4'hc):(3'h7)],
              (~reg1071[(3'h6):(1'h0)])};
          reg1086 <= reg1049[(2'h2):(1'h0)];
          reg1087 <= (~(($unsigned((reg1016 ? reg1086 : (7'h57))) << reg1049) ?
              reg1032[(4'hf):(3'h4)] : reg1086[(5'h10):(1'h0)]));
          if ($unsigned(reg1074))
            begin
              reg1088 <= reg1024[(1'h1):(1'h0)];
              reg1089 <= $signed($unsigned($unsigned((!forvar1083[(1'h1):(1'h0)]))));
              reg1090 = $signed(reg1038);
              reg1091 = reg1074;
            end
          else
            begin
              reg1090 = {(~|wire1007[(1'h0):(1'h0)])};
              reg1092 <= $signed($signed(((&(7'h4a)) ?
                  ($signed(wire1009) ?
                      $unsigned((7'h4b)) : reg1074[(5'h12):(4'hc)]) : reg1087[(4'h8):(1'h1)])));
              reg1093 <= (~^(~^reg1012));
              reg1094 <= $signed(($signed({$signed(reg1086)}) ?
                  $signed(reg1055[(1'h1):(1'h0)]) : $unsigned((((8'hbb) && (7'h54)) ?
                      $signed(wire1082) : (reg1071 == reg1015)))));
              reg1095 = {reg1091};
              reg1096 <= $unsigned(((|$signed(reg1012[(4'h8):(2'h2)])) ^~ (($signed(wire1010) < reg1087) ^ ($unsigned(reg1078) ?
                  $signed(reg1027) : (reg1043 ? reg1013 : reg1048)))));
              reg1097 = reg1074;
            end
        end
      reg1098 = (wire1008[(3'h7):(1'h0)] ?
          reg1053 : (~|$unsigned(wire1082[(3'h6):(3'h4)])));
      if (reg1094[(3'h7):(3'h7)])
        begin
          reg1099 <= ($unsigned($signed($unsigned($unsigned(reg1087)))) ?
              (~&reg1016) : reg1056);
          if ($signed($signed(((reg1048 == $unsigned(reg1013)) == {(reg1055 <<< reg1070),
              (reg1035 < reg1070)}))))
            begin
              reg1100 <= {wire1006};
              reg1101 <= reg1035;
              reg1102 <= $signed($unsigned((~&reg1078)));
            end
          else
            begin
              reg1103 = $unsigned((~&$signed(($signed(wire1008) < $unsigned((7'h47))))));
              reg1104 = ((~$signed((^~wire1082[(4'ha):(3'h6)]))) ?
                  (|(reg1074 * $signed((~^reg1102)))) : $unsigned(({(-reg1102),
                      (reg1074 <= (8'hb7)),
                      $signed(reg1033)} || (!(reg1032 ? reg1085 : wire1010)))));
            end
          if ((!{((reg1104 ?
                  $signed(reg1016) : $unsigned(reg1077)) >> ($unsigned(reg1095) < (7'h4d))),
              $unsigned(reg1093)}))
            begin
              reg1105 = $signed((8'hb3));
              reg1106 <= $signed(((|wire1010[(2'h2):(1'h0)]) ?
                  $signed(reg1049[(3'h6):(3'h6)]) : ($signed($unsigned(reg1076)) <<< reg1093[(3'h5):(1'h1)])));
              reg1107 = $unsigned(reg1056[(3'h4):(1'h1)]);
              reg1108 = (8'hb8);
              reg1109 = $signed({($signed(reg1055[(2'h3):(1'h1)]) ?
                      ($signed(reg1030) ^~ $signed(reg1042)) : reg1011),
                  $unsigned($unsigned($unsigned(reg1015)))});
              reg1110 = (((reg1089 ? (+$unsigned(reg1100)) : reg1030) ?
                      reg1105 : ($unsigned((^~(8'h9d))) <<< (~|(reg1056 ?
                          (7'h58) : reg1092)))) ?
                  (~^(~|$signed(reg1107))) : (~|{(~reg1050)}));
              reg1111 = (reg1071 ?
                  (~^reg1095[(1'h1):(1'h0)]) : $unsigned((~(wire1008 ?
                      (!reg1096) : reg1098))));
            end
          else
            begin
              reg1106 <= reg1087;
              reg1112 <= ($unsigned(wire1009[(3'h6):(3'h5)]) ~^ $signed(reg1013[(3'h6):(2'h3)]));
            end
          reg1113 = {((~&(7'h45)) ?
                  {$unsigned($signed(reg1104))} : reg1111[(4'hc):(3'h6)])};
          reg1114 = (reg1035 && $unsigned(reg1097[(3'h4):(2'h3)]));
        end
      else
        begin
          reg1103 = $unsigned(($unsigned(($unsigned(wire1006) ^ (reg1043 != (8'ha2)))) >= reg1011));
        end
      if (reg1105)
        begin
          reg1115 = $unsigned($signed($signed((~reg1113))));
          if ((~(reg1090 ^ reg1066)))
            begin
              reg1116 = reg1087[(4'hb):(2'h3)];
              reg1117 <= ({$signed(((wire1009 != reg1078) ?
                          reg1033[(4'he):(1'h1)] : (wire1082 >> reg1050))),
                      (+(reg1030 || reg1053[(4'hb):(3'h7)])),
                      (^~$signed({reg1087}))} ?
                  $signed(($signed((reg1011 ?
                      reg1114 : reg1077)) + ($signed(reg1104) ?
                      reg1035 : (reg1049 ?
                          reg1084 : reg1074)))) : ($unsigned((reg1043[(3'h5):(1'h1)] ?
                          (reg1096 & (8'hb2)) : {reg1085, reg1025, reg1115})) ?
                      (8'hac) : (~(^reg1090[(4'hf):(3'h6)]))));
              reg1118 <= $signed((^reg1089[(4'h9):(3'h4)]));
              reg1119 = ((^~(reg1090[(4'h8):(3'h4)] ?
                  reg1027[(4'h9):(2'h2)] : $unsigned($signed(reg1105)))) + (8'ha4));
              reg1120 = (7'h44);
              reg1121 <= ({reg1091,
                      (((|reg1110) == (reg1103 ? (7'h45) : forvar1083)) ?
                          (-(reg1098 ? reg1077 : (8'hb6))) : (8'hb3))} ?
                  reg1050[(2'h3):(1'h1)] : (7'h49));
              reg1122 <= reg1119[(4'hb):(4'h9)];
            end
          else
            begin
              reg1117 <= (reg1118 ?
                  $signed(((((7'h4e) ? (8'ha0) : (8'ha9)) == $signed((8'ha3))) ?
                      ((^~reg1097) >> ((8'had) ?
                          wire1009 : reg1035)) : ((!reg1030) < {reg1012}))) : (^(reg1119[(5'h10):(3'h7)] ?
                      (|reg1092[(1'h0):(1'h0)]) : reg1015)));
              reg1118 <= {reg1048[(2'h3):(1'h0)], reg1089};
              reg1119 = ($unsigned(reg1055[(3'h4):(3'h4)]) == $unsigned(reg1093));
              reg1120 = wire1010;
              reg1123 = {($unsigned({$unsigned(reg1034),
                      reg1011}) - {forvar1083,
                      (^~reg1033[(2'h3):(1'h1)]),
                      (8'ha9)})};
              reg1124 <= $unsigned($signed((7'h56)));
            end
          for (forvar1125 = (1'h0); (forvar1125 < (3'h5)); forvar1125 = (forvar1125 + (1'h1)))
            begin
              reg1126 <= reg1042;
              reg1127 <= {(reg1111[(2'h2):(1'h0)] ?
                      reg1024[(4'hb):(4'ha)] : reg1110),
                  $unsigned(($unsigned($signed((8'ha2))) ?
                      (7'h47) : reg1092[(1'h0):(1'h0)])),
                  {(~(reg1092 + reg1087))}};
              reg1128 = (^(^~reg1116));
              reg1129 = ((|$signed(((reg1119 - reg1086) | (reg1071 != reg1012)))) - reg1122);
              reg1130 <= reg1112[(2'h3):(2'h2)];
            end
          for (forvar1131 = (1'h0); (forvar1131 < (3'h4)); forvar1131 = (forvar1131 + (1'h1)))
            begin
              reg1132 <= reg1127;
            end
          if ($unsigned($signed((reg1048 < $unsigned($signed(reg1030))))))
            begin
              reg1133 <= ((!reg1024) ^~ reg1024[(5'h10):(3'h6)]);
              reg1134 = ($unsigned(((~&(reg1024 ? reg1130 : reg1093)) ?
                  (7'h4a) : $unsigned((reg1123 >> reg1124)))) * $signed((7'h49)));
              reg1135 = $unsigned(forvar1125);
            end
          else
            begin
              reg1133 <= (8'hb5);
              reg1136 <= (|($signed($unsigned(reg1088[(2'h3):(2'h2)])) ?
                  $unsigned((forvar1083[(1'h1):(1'h0)] <<< reg1133)) : $unsigned($signed((reg1050 ?
                      reg1053 : reg1133)))));
              reg1137 = wire1006[(5'h12):(4'hb)];
              reg1138 <= reg1013;
              reg1139 <= forvar1083[(1'h0):(1'h0)];
              reg1140 = reg1106;
            end
          for (forvar1141 = (1'h0); (forvar1141 < (2'h3)); forvar1141 = (forvar1141 + (1'h1)))
            begin
              reg1142 <= $signed((~^($signed($signed(reg1112)) ?
                  (reg1118 ?
                      $signed(reg1098) : {reg1091,
                          reg1121,
                          (7'h53)}) : ((~|wire1006) != (|reg1030)))));
            end
        end
      else
        begin
          for (forvar1115 = (1'h0); (forvar1115 < (3'h5)); forvar1115 = (forvar1115 + (1'h1)))
            begin
              reg1116 = reg1108[(3'h6):(2'h3)];
              reg1117 <= $signed($signed($signed($unsigned(reg1053[(3'h5):(3'h5)]))));
              reg1118 <= $signed((7'h4f));
            end
          reg1121 <= reg1025[(1'h0):(1'h0)];
          for (forvar1122 = (1'h0); (forvar1122 < (3'h5)); forvar1122 = (forvar1122 + (1'h1)))
            begin
              reg1123 = reg1035[(5'h1e):(3'h7)];
            end
          reg1125 = {$unsigned(reg1104),
              reg1030,
              (+$unsigned((~|reg1107[(4'he):(2'h3)])))};
          reg1126 <= forvar1115[(4'h9):(3'h6)];
          reg1127 <= $unsigned(($signed($signed((reg1093 == reg1090))) ?
              (7'h56) : reg1024));
        end
      reg1143 = {(~&(8'hb7)),
          ($unsigned((~&$signed(reg1056))) <<< reg1042),
          (reg1105[(4'hb):(4'h8)] ?
              {$unsigned({reg1113, (7'h46), reg1140}),
                  $unsigned((reg1120 ?
                      wire1010 : reg1033))} : $unsigned(reg1032))};
      if ($unsigned(($signed(((^reg1101) ?
          ((8'hbc) == reg1103) : $signed(reg1130))) != reg1102[(1'h1):(1'h0)])))
        begin
          if ($unsigned($signed(reg1084)))
            begin
              reg1144 <= (8'hac);
              reg1145 <= ((7'h54) == (($unsigned((~^reg1096)) ?
                      reg1116[(3'h4):(2'h3)] : ((reg1115 ? reg1076 : (7'h4c)) ?
                          reg1110 : (reg1122 ? reg1101 : reg1116))) ?
                  reg1034 : (reg1113[(1'h0):(1'h0)] ?
                      ($signed(reg1016) ?
                          (forvar1125 ?
                              (8'hba) : forvar1122) : forvar1115[(1'h1):(1'h1)]) : reg1144)));
              reg1146 <= (((^(~^$signed(reg1087))) ?
                  $unsigned($unsigned({reg1100})) : reg1109) ^ $unsigned((7'h40)));
              reg1147 = $unsigned($unsigned(reg1066[(2'h3):(2'h2)]));
            end
          else
            begin
              reg1147 = $unsigned($signed((|(reg1127 ^~ $signed(reg1097)))));
              reg1148 <= reg1089;
              reg1149 <= reg1070;
              reg1150 = $unsigned($unsigned(reg1095[(2'h2):(1'h1)]));
              reg1151 <= $unsigned($signed((reg1148 <<< {$unsigned(reg1066)})));
              reg1152 <= ((-(((!reg1136) >= (wire1010 ? reg1078 : forvar1122)) ?
                  reg1140[(3'h7):(3'h5)] : $signed($unsigned(reg1027)))) >> (&(((reg1089 ?
                          wire1010 : reg1146) ?
                      reg1077 : $unsigned(reg1016)) ?
                  reg1137[(5'h14):(4'hd)] : $unsigned(reg1151))));
              reg1153 = {$unsigned(((reg1041 ?
                      (~&(7'h42)) : $unsigned(reg1117)) + (-reg1076)))};
            end
        end
      else
        begin
          reg1147 = (!(reg1092 < (((^~reg1035) ^ {(8'had)}) ?
              $signed(reg1066) : $signed((reg1123 ? reg1103 : reg1138)))));
          for (forvar1148 = (1'h0); (forvar1148 < (2'h3)); forvar1148 = (forvar1148 + (1'h1)))
            begin
              reg1149 <= (^~reg1084[(4'h8):(4'h8)]);
              reg1151 <= ((~((((8'hb1) | reg1032) ~^ wire1006[(4'hc):(4'ha)]) ?
                      reg1070 : reg1106)) ?
                  reg1092[(2'h2):(1'h0)] : wire1082[(2'h2):(1'h1)]);
              reg1153 = $unsigned($unsigned($unsigned(((~^reg1121) ?
                  (^~reg1140) : forvar1125[(4'hc):(3'h6)]))));
              reg1154 = (reg1086[(4'ha):(3'h6)] ?
                  reg1109[(5'h14):(4'hd)] : ({($unsigned(reg1108) << (reg1153 ?
                              reg1016 : reg1097))} ?
                      ((((7'h43) - reg1032) ?
                          $unsigned(reg1092) : $unsigned(reg1135)) * $signed($unsigned(reg1099))) : (reg1050[(4'ha):(4'ha)] <<< (~^$unsigned(wire1008)))));
              reg1155 <= ($signed($unsigned((~&(-reg1011)))) <<< $signed(reg1116));
              reg1156 <= {$unsigned(reg1153[(3'h6):(3'h5)])};
              reg1157 = reg1050[(4'hb):(4'h8)];
            end
          if (reg1153)
            begin
              reg1158 <= ((|$unsigned(reg1113)) ?
                  reg1041 : (reg1090[(2'h3):(2'h2)] << reg1038[(3'h4):(2'h2)]));
              reg1159 <= (^~reg1093[(5'h12):(4'he)]);
            end
          else
            begin
              reg1158 <= $unsigned((7'h4e));
              reg1160 = {$signed(((|(~|reg1153)) << $signed((~&reg1077)))),
                  ($signed(reg1119[(4'ha):(3'h5)]) ?
                      $signed(((reg1119 ^ reg1102) >> reg1033)) : $signed((reg1155 <= reg1043))),
                  reg1090[(4'hc):(1'h0)]};
              reg1161 <= ($signed(reg1086[(3'h6):(3'h4)]) << (forvar1083[(1'h1):(1'h0)] & ($signed(reg1103) >= {$signed(reg1087),
                  (reg1155 ? reg1144 : reg1127)})));
              reg1162 = wire1010;
              reg1163 = (!$unsigned($signed($unsigned(reg1077))));
              reg1164 = (reg1107 ?
                  {reg1156[(2'h2):(1'h1)]} : ($signed(reg1162) * $signed((~{reg1012}))));
              reg1165 <= (($unsigned({(8'ha6)}) ?
                      forvar1122 : ($signed(reg1024) ?
                          $signed({reg1066}) : (^~{(7'h53),
                              reg1066,
                              reg1071}))) ?
                  reg1015 : (^{(((8'hb7) ?
                          reg1105 : (8'ha5)) + wire1006[(4'hb):(4'h9)]),
                      $signed(reg1164)}));
            end
          reg1166 = (^~forvar1115);
          reg1167 <= reg1102;
          reg1168 = ($unsigned(({$unsigned(wire1008)} ?
                  $unsigned(reg1160[(4'he):(1'h0)]) : reg1033)) ?
              (reg1085 <= reg1115) : ($unsigned(reg1077[(5'h17):(4'ha)]) ?
                  {(^reg1140[(4'ha):(3'h5)])} : reg1108[(4'ha):(2'h3)]));
          for (forvar1169 = (1'h0); (forvar1169 < (1'h0)); forvar1169 = (forvar1169 + (1'h1)))
            begin
              reg1170 <= $unsigned(reg1052[(2'h2):(1'h1)]);
            end
        end
      reg1171 = {(-wire1008)};
    end
  always
    @(posedge clk) begin
      reg1172 <= (($unsigned((&reg1132)) ?
          ($signed(reg1159) ?
              reg1145 : $signed((7'h57))) : $unsigned((reg1148 >>> $unsigned(reg1144)))) & reg1012);
      if ((reg1146[(3'h5):(3'h5)] || reg1117))
        begin
          reg1173 = (^~(reg1112 ?
              ((reg1071[(5'h17):(1'h1)] ?
                  wire1008 : {reg1112,
                      reg1132,
                      wire1010}) ^~ ($unsigned(reg1170) ?
                  (reg1066 <<< (7'h45)) : (|reg1076))) : $signed(((~&(7'h4c)) ?
                  reg1092[(4'hc):(3'h4)] : {reg1030, reg1124}))));
          reg1174 = reg1167[(3'h6):(2'h3)];
          for (forvar1175 = (1'h0); (forvar1175 < (3'h5)); forvar1175 = (forvar1175 + (1'h1)))
            begin
              reg1176 = (reg1145[(4'he):(1'h0)] & reg1048);
              reg1177 <= (reg1033[(4'h8):(2'h2)] * ({reg1148[(4'hb):(1'h1)]} * $unsigned(reg1145)));
            end
          reg1178 = $unsigned((~|$unsigned($unsigned($signed(reg1016)))));
          if (reg1174)
            begin
              reg1179 <= ((((reg1032[(4'h9):(1'h0)] ?
                      (reg1174 ? reg1099 : reg1136) : $signed((8'hbb))) ?
                  $signed(reg1149[(4'he):(2'h3)]) : $signed($signed((7'h57)))) > ((((8'hbe) ?
                          reg1092 : reg1118) ?
                      $unsigned(reg1027) : (reg1071 ? reg1173 : reg1078)) ?
                  reg1161 : $signed(reg1035[(5'h1f):(4'ha)]))) | $signed((+reg1117[(1'h1):(1'h0)])));
              reg1180 = ($signed((&reg1093)) <<< $signed((reg1055 | (+$signed(reg1145)))));
            end
          else
            begin
              reg1179 <= (|$unsigned(reg1092[(2'h2):(1'h0)]));
              reg1180 = $signed($signed(((8'had) ?
                  reg1170[(4'hf):(4'hc)] : (~&$unsigned((8'hb3))))));
              reg1181 = reg1130;
            end
          if ((&$signed((reg1170[(3'h6):(1'h1)] ?
              (reg1066 | (reg1013 ?
                  reg1142 : reg1074)) : ((reg1052 << reg1112) >>> reg1130[(3'h4):(2'h3)])))))
            begin
              reg1182 = ($signed(reg1050) ?
                  ($signed(reg1033) - $signed($signed(((8'hae) & reg1056)))) : {(reg1032[(4'hc):(2'h3)] ?
                          reg1012[(3'h6):(2'h3)] : ((reg1099 ?
                                  reg1070 : reg1048) ?
                              $unsigned((8'hbb)) : reg1180))});
            end
          else
            begin
              reg1183 <= (reg1043[(2'h3):(2'h2)] + ((reg1078[(3'h5):(2'h3)] && $unsigned($unsigned(reg1074))) & (&reg1126)));
            end
          reg1184 <= reg1070;
        end
      else
        begin
          reg1175 <= reg1086;
          reg1177 <= ($signed(reg1093) | reg1172);
          if (reg1138[(4'hf):(3'h7)])
            begin
              reg1179 <= (~|(reg1085 ?
                  (~$signed(reg1032[(5'h11):(3'h7)])) : $unsigned((!(reg1076 + reg1159)))));
              reg1180 = $unsigned((^{$signed(reg1099[(1'h0):(1'h0)]),
                  reg1052[(1'h1):(1'h1)]}));
              reg1183 <= wire1007;
              reg1184 <= (&$unsigned(reg1136[(4'ha):(4'ha)]));
            end
          else
            begin
              reg1179 <= ($signed((($signed(reg1152) + reg1078[(3'h5):(3'h4)]) ?
                      {((7'h41) & reg1043), (7'h4a), {(7'h57)}} : ((^~(8'hbf)) ?
                          (reg1133 != reg1092) : ((7'h43) ?
                              reg1132 : reg1136)))) ?
                  (|(+$unsigned($unsigned(reg1156)))) : ($unsigned((7'h46)) ?
                      (7'h4b) : ($signed($signed(reg1155)) || reg1148)));
              reg1180 = reg1182;
              reg1181 = wire1009[(3'h6):(3'h4)];
              reg1182 = $unsigned(($unsigned(reg1038) ?
                  $signed(reg1048[(2'h3):(1'h0)]) : {reg1139[(2'h3):(1'h1)]}));
              reg1185 = ($signed(reg1086) < $signed($signed(reg1184)));
              reg1186 = {((~(~^(reg1077 ?
                      reg1030 : reg1030))) >>> $signed(($signed(reg1035) == $unsigned(reg1122))))};
              reg1187 <= $signed(((7'h4a) ?
                  $signed(reg1181) : (reg1089 ?
                      reg1133[(2'h2):(1'h0)] : $signed((reg1127 * reg1033)))));
            end
          reg1188 <= $unsigned({($signed((8'had)) ?
                  (((7'h41) ? (7'h52) : reg1087) ~^ (-reg1138)) : (8'hbc)),
              (&$unsigned((+reg1035)))});
        end
      reg1189 <= (|(~|reg1012[(3'h4):(2'h2)]));
      if ($signed(($unsigned((reg1056[(3'h4):(1'h0)] >> $unsigned(reg1170))) == $unsigned({$signed(reg1041)}))))
        begin
          if ((&{$signed((&{reg1180}))}))
            begin
              reg1190 = (8'hab);
              reg1191 <= (!{(((reg1032 || (8'hac)) >>> (~|reg1066)) == ($signed((8'ha2)) <= ((8'hae) ?
                      (7'h51) : reg1027))),
                  reg1015,
                  (~|$signed((reg1024 >> reg1078)))});
              reg1192 <= $unsigned(reg1034[(4'ha):(3'h7)]);
              reg1193 <= reg1034;
              reg1194 <= (~|reg1158[(5'h13):(4'he)]);
              reg1195 = (((!(((8'hbe) | reg1025) < (reg1145 ?
                  reg1118 : reg1087))) || $signed($signed((reg1038 ?
                  reg1148 : (8'ha4))))) <<< reg1186[(5'h10):(1'h0)]);
            end
          else
            begin
              reg1190 = $signed(((|($unsigned(reg1034) ?
                  {reg1033, (7'h53)} : (7'h41))) < (reg1035[(5'h1c):(3'h4)] ?
                  {reg1056} : $unsigned(reg1024))));
              reg1191 <= ((~^$signed((reg1167 ?
                  ((8'hb4) | reg1148) : (reg1133 != reg1151)))) << (($unsigned((~&wire1082)) ^~ $signed(reg1112[(2'h3):(2'h3)])) ?
                  (+((reg1145 > (7'h4a)) ?
                      $unsigned((7'h40)) : ((8'hbf) ?
                          reg1013 : reg1158))) : (+reg1191)));
              reg1195 = (+wire1009[(1'h0):(1'h0)]);
            end
          for (forvar1196 = (1'h0); (forvar1196 < (1'h0)); forvar1196 = (forvar1196 + (1'h1)))
            begin
              reg1197 <= reg1170[(5'h12):(4'ha)];
              reg1198 <= (~|(reg1117[(3'h4):(3'h4)] ?
                  (^~reg1165[(2'h2):(1'h0)]) : (~reg1100)));
              reg1199 = $unsigned(reg1155[(3'h6):(1'h1)]);
              reg1200 = ((~^reg1088) <<< reg1146);
              reg1201 = reg1158[(5'h1c):(5'h1c)];
              reg1202 = (-$unsigned($signed($unsigned($unsigned((7'h47))))));
            end
          reg1203 <= $unsigned($signed((&(reg1013 & (reg1013 >= reg1042)))));
          for (forvar1204 = (1'h0); (forvar1204 < (2'h2)); forvar1204 = (forvar1204 + (1'h1)))
            begin
              reg1205 = (&$unsigned(((7'h4b) <= ({reg1043, (8'hba), (7'h57)} ?
                  {reg1148, reg1200} : $signed(reg1189)))));
            end
          if ((8'ha6))
            begin
              reg1206 <= (forvar1196 ?
                  ((7'h58) >>> reg1112[(2'h3):(2'h2)]) : (&reg1198));
              reg1207 <= {(~(reg1192[(5'h19):(5'h14)] ? wire1008 : (8'ha7))),
                  (~|reg1118[(5'h1a):(4'h9)]),
                  $signed($signed((^reg1089)))};
              reg1208 <= reg1056[(4'h8):(2'h2)];
              reg1209 = reg1027;
              reg1210 = ((reg1121 ?
                      (((reg1190 ? (8'hb9) : reg1096) ?
                              $signed(reg1013) : ((7'h46) + reg1191)) ?
                          ((reg1130 ?
                              reg1139 : reg1013) <<< (-(7'h53))) : $unsigned($signed((8'hb8)))) : $unsigned(reg1034[(2'h2):(2'h2)])) ?
                  {reg1112} : reg1138);
            end
          else
            begin
              reg1209 = (!$unsigned((|reg1093)));
              reg1210 = {reg1133[(2'h3):(2'h2)]};
            end
          if ($signed((7'h48)))
            begin
              reg1211 = $signed((~(((reg1144 ? (7'h55) : (7'h56)) ?
                      {reg1096} : $signed(reg1208)) ?
                  $signed(reg1158) : ((reg1184 != forvar1196) ?
                      $signed((7'h58)) : reg1193[(3'h4):(3'h4)]))));
              reg1212 = reg1177;
              reg1213 = $unsigned((reg1158 ?
                  ($signed((~|reg1174)) ^ reg1187[(4'h8):(3'h4)]) : $signed(reg1100)));
              reg1214 = reg1013;
              reg1215 = (~|{((reg1049[(1'h0):(1'h0)] ?
                          {reg1066} : $unsigned(reg1142)) ?
                      reg1016 : reg1172[(4'h8):(2'h3)])});
              reg1216 <= (8'ha8);
              reg1217 = (reg1179 ?
                  reg1208 : ($signed($unsigned(((7'h42) ? reg1071 : reg1085))) ?
                      ($unsigned((reg1032 & reg1071)) || $unsigned(reg1112[(1'h1):(1'h0)])) : reg1155));
            end
          else
            begin
              reg1216 <= {{($signed({(7'h40)}) - (&reg1053[(3'h7):(1'h0)])),
                      ((~$signed(reg1043)) ?
                          $unsigned((reg1187 ?
                              reg1130 : reg1041)) : $unsigned(reg1088[(1'h0):(1'h0)]))},
                  ((reg1100[(5'h14):(3'h7)] ?
                      reg1033[(3'h6):(1'h0)] : {(~|reg1106)}) ^ reg1173)};
              reg1218 <= (~|($signed({(reg1174 ? reg1074 : (8'haa)),
                  (7'h4f)}) < $unsigned($unsigned(reg1206))));
              reg1219 <= $signed((&{{(reg1074 ? reg1185 : (7'h40)),
                      $signed(reg1142),
                      reg1211[(5'h12):(4'h8)]}}));
              reg1220 = (^~reg1130[(3'h6):(3'h4)]);
              reg1221 <= reg1118[(5'h1a):(5'h13)];
              reg1222 <= reg1179[(3'h7):(2'h2)];
            end
          reg1223 = (^~$signed(reg1187[(3'h4):(2'h2)]));
        end
      else
        begin
          for (forvar1190 = (1'h0); (forvar1190 < (3'h4)); forvar1190 = (forvar1190 + (1'h1)))
            begin
              reg1191 <= reg1159[(3'h5):(3'h5)];
              reg1192 <= $unsigned((($unsigned((reg1032 ? reg1149 : reg1206)) ?
                      (^(reg1027 | reg1049)) : $unsigned(((8'hb8) ?
                          reg1027 : reg1038))) ?
                  forvar1175[(3'h6):(1'h0)] : ({reg1146[(2'h2):(2'h2)]} <= $unsigned(reg1087))));
              reg1195 = (($signed((~^((7'h49) ?
                      reg1152 : (8'had)))) - ((~|((8'hb2) ?
                          reg1094 : reg1042)) ?
                      {(reg1183 ? (8'ha8) : reg1180)} : ($signed(reg1176) ?
                          $unsigned(reg1094) : $unsigned(reg1152)))) ?
                  (^~$unsigned((reg1034 ?
                      reg1144 : (reg1145 ~^ (7'h50))))) : {reg1138[(4'he):(4'hb)]});
              reg1196 <= reg1172;
              reg1199 = reg1013[(3'h5):(3'h5)];
            end
          for (forvar1200 = (1'h0); (forvar1200 < (2'h2)); forvar1200 = (forvar1200 + (1'h1)))
            begin
              reg1203 <= {((7'h48) ?
                      reg1193 : ((|(reg1092 ~^ reg1077)) ?
                          $signed(reg1133) : reg1155[(2'h3):(1'h0)]))};
              reg1204 <= $unsigned(reg1208[(1'h1):(1'h1)]);
            end
          if ($unsigned($signed($unsigned($signed($signed(reg1096))))))
            begin
              reg1205 = {$unsigned($unsigned($unsigned($signed(reg1130))))};
              reg1206 <= ($unsigned(((|reg1130) & {$unsigned((8'hbd)),
                      ((7'h4e) != reg1213)})) ?
                  $unsigned((((reg1206 ?
                      reg1112 : reg1112) == reg1176[(3'h5):(1'h0)]) != (reg1016 ?
                      $signed(reg1078) : (reg1156 || reg1189)))) : $unsigned($signed($signed(((8'hb8) ?
                      reg1187 : reg1035)))));
              reg1207 <= (((($unsigned((8'hb6)) ?
                      (reg1015 ~^ reg1179) : reg1066) | reg1196[(4'h9):(2'h3)]) && reg1025[(3'h5):(2'h3)]) ?
                  (wire1082 | $signed($unsigned(reg1212))) : $signed($unsigned({(reg1100 ?
                          reg1112 : reg1016),
                      forvar1200,
                      ((7'h57) * reg1012)})));
              reg1209 = (^~({(+reg1127)} ~^ $unsigned(reg1159[(3'h6):(1'h1)])));
            end
          else
            begin
              reg1205 = reg1013[(4'he):(4'h8)];
              reg1209 = reg1011[(5'h14):(4'hc)];
              reg1216 <= (reg1217 & $signed(((+reg1126[(4'h8):(3'h5)]) && $unsigned({(8'hb6),
                  reg1175,
                  reg1190}))));
              reg1218 <= ((~&reg1118) ?
                  ({{(reg1148 ?
                              (7'h4e) : reg1127)}} ~^ $signed((8'ha2))) : (~^((~$unsigned(reg1155)) ?
                      {forvar1175, reg1086} : $signed(((8'hb3) ?
                          reg1185 : reg1218)))));
            end
          if ((-(&$unsigned(reg1156))))
            begin
              reg1219 <= (~|(reg1093 >= ((+$signed((8'ha7))) >= $signed(((7'h42) + reg1027)))));
              reg1221 <= forvar1175[(1'h1):(1'h1)];
              reg1222 <= reg1038[(1'h1):(1'h0)];
              reg1223 = reg1133;
              reg1224 = $unsigned(($signed((~(reg1087 ?
                  reg1206 : reg1175))) <= forvar1190));
            end
          else
            begin
              reg1220 = reg1099[(3'h5):(3'h4)];
              reg1221 <= {((~&$signed((reg1066 ? (8'hae) : reg1179))) ?
                      ($unsigned((forvar1200 ? reg1167 : reg1012)) ?
                          {(|reg1011),
                              {reg1205, reg1076},
                              $signed(reg1223)} : {(&reg1132),
                              (7'h51),
                              $signed(reg1186)}) : (7'h48)),
                  $signed($unsigned($signed((reg1174 ? reg1216 : reg1041)))),
                  $unsigned($signed(reg1155))};
              reg1223 = $signed((~^$signed(reg1146[(3'h5):(1'h1)])));
              reg1224 = ($signed(reg1156[(4'h8):(3'h4)]) ?
                  ($signed(reg1192) == (((reg1179 & reg1181) != {reg1156}) >>> (reg1042 ?
                      $unsigned(reg1088) : $signed(reg1172)))) : $unsigned(reg1186));
              reg1225 <= (^~($signed($signed((!reg1152))) << ({(^reg1042)} << (|reg1127))));
            end
        end
    end
  assign wire1226 = $unsigned($unsigned(reg1056));
  always
    @(posedge clk) begin
      reg1227 <= (((8'hab) ? reg1088 : reg1096) ?
          (-((((8'hb9) ? reg1121 : (8'ha8)) * (reg1192 ^ (8'hbb))) ?
              (~(reg1049 << reg1106)) : (reg1225[(2'h2):(1'h1)] + $unsigned(reg1102)))) : reg1148);
    end
  assign wire1228 = $signed(($unsigned((!reg1049[(3'h5):(3'h5)])) ?
                        reg1159[(3'h5):(2'h3)] : reg1106[(5'h12):(4'h8)]));
  assign wire1229 = reg1070[(5'h11):(4'h8)];
  assign wire1230 = (8'haa);
  assign wire1231 = reg1170;
  always
    @(posedge clk) begin
      for (forvar1232 = (1'h0); (forvar1232 < (3'h4)); forvar1232 = (forvar1232 + (1'h1)))
        begin
          if (reg1172)
            begin
              reg1233 = $unsigned((^~$signed(((reg1035 ?
                  reg1127 : reg1086) & (reg1225 ? reg1100 : reg1138)))));
              reg1234 = (reg1124[(5'h18):(3'h5)] & $signed(($unsigned((reg1184 ~^ reg1206)) < ((reg1148 == reg1049) <<< $signed(reg1159)))));
              reg1235 <= reg1196;
              reg1236 <= $signed($signed((&{$signed(reg1011)})));
              reg1237 <= reg1204;
              reg1238 <= $signed(reg1100[(5'h10):(2'h2)]);
              reg1239 = ($unsigned($signed(($signed(reg1187) ?
                      reg1179 : $unsigned(reg1148)))) ?
                  $signed(((^~$unsigned((8'h9f))) ?
                      (~(reg1221 && reg1102)) : (!reg1027[(2'h2):(1'h1)]))) : $unsigned((reg1170 ?
                      reg1074[(4'ha):(1'h0)] : (reg1076 ?
                          $unsigned((8'hb0)) : (reg1117 < reg1132)))));
            end
          else
            begin
              reg1235 <= $unsigned((|(reg1074 ?
                  ({reg1221, forvar1232} << {reg1034,
                      reg1034,
                      (8'hbb)}) : ((8'hb6) ? {reg1121} : $unsigned(reg1086)))));
            end
          reg1240 = {{reg1170[(3'h4):(2'h2)]}};
          reg1241 <= $signed((reg1240[(4'h8):(2'h3)] ?
              (~&(|{reg1035, reg1218, reg1027})) : ($signed($signed(reg1088)) ?
                  (reg1032[(4'he):(2'h3)] ?
                      (^wire1229) : (reg1206 < reg1151)) : (((7'h4e) ?
                          reg1234 : reg1077) ?
                      {(7'h44), reg1145} : {reg1218, reg1130}))));
          reg1242 = (({(wire1007 ? ((8'hb9) <= reg1235) : $unsigned(reg1145)),
                      $signed($signed(reg1235))} ?
                  (!(-$signed(reg1011))) : (+((reg1066 >> wire1082) & (^~reg1233)))) ?
              reg1102 : {reg1066[(2'h2):(1'h1)], reg1048});
          for (forvar1243 = (1'h0); (forvar1243 < (3'h4)); forvar1243 = (forvar1243 + (1'h1)))
            begin
              reg1244 = (($signed(((-reg1146) ?
                      reg1197[(5'h15):(5'h10)] : reg1239[(4'ha):(4'ha)])) == (reg1238 << $unsigned($signed(reg1043)))) ?
                  {(8'ha4),
                      (reg1013 ?
                          (~|(reg1038 ?
                              reg1024 : reg1070)) : reg1074[(5'h13):(4'h9)]),
                      (($signed(reg1208) >>> $signed(reg1175)) ?
                          (+(reg1076 ?
                              reg1207 : reg1076)) : (((7'h4f) ^~ reg1197) ?
                              reg1188[(2'h2):(1'h1)] : (reg1239 ^~ reg1024)))} : ((8'hae) ?
                      reg1138[(3'h4):(2'h2)] : wire1230[(5'h15):(3'h4)]));
            end
          if ($signed((((reg1024[(4'hb):(4'hb)] ?
                  (8'hb9) : (reg1092 ? reg1071 : reg1239)) == {{reg1133},
                  (&reg1225)}) ?
              reg1237 : reg1156)))
            begin
              reg1245 <= (^~(&(reg1066[(2'h2):(1'h0)] ?
                  ($unsigned(reg1094) ?
                      (7'h49) : $unsigned(reg1240)) : ($unsigned(reg1092) ?
                      (!forvar1243) : $signed(reg1038)))));
              reg1246 <= (-({(reg1094 < $signed((8'hbf))),
                  reg1049[(1'h1):(1'h0)],
                  ($signed(reg1130) * (reg1102 >>> (8'h9e)))} == reg1025));
              reg1247 = ((~|$signed($signed((reg1242 == wire1008)))) - ($signed({$unsigned(reg1122)}) ?
                  (!$unsigned(reg1124)) : (^~wire1006)));
              reg1248 = wire1230[(5'h14):(1'h0)];
              reg1249 = $unsigned({$unsigned((~&reg1099[(2'h2):(1'h0)])),
                  {reg1207[(2'h2):(1'h1)], $unsigned((!forvar1232))},
                  $signed($unsigned(((8'hb1) ? reg1050 : reg1112)))});
            end
          else
            begin
              reg1245 <= {reg1074};
            end
        end
      reg1250 = reg1233;
      reg1251 <= (reg1117[(4'h8):(3'h6)] ?
          ({$signed(((8'haa) ? reg1087 : reg1241)), (8'ha9)} ?
              reg1027 : (((~|reg1250) ? (^reg1078) : {reg1194}) ?
                  $signed($signed(reg1235)) : {$signed(reg1027),
                      reg1148,
                      reg1161[(3'h7):(2'h3)]})) : (($signed(reg1175) ?
              (reg1197[(5'h13):(4'hd)] ?
                  (reg1117 | reg1155) : wire1229) : (^~(reg1184 > reg1043))) && $unsigned(reg1066)));
      for (forvar1252 = (1'h0); (forvar1252 < (1'h1)); forvar1252 = (forvar1252 + (1'h1)))
        begin
          reg1253 = reg1239;
          reg1254 <= reg1152[(5'h17):(2'h3)];
          reg1255 = (^(wire1229 ^ wire1082));
        end
      for (forvar1256 = (1'h0); (forvar1256 < (3'h6)); forvar1256 = (forvar1256 + (1'h1)))
        begin
          for (forvar1257 = (1'h0); (forvar1257 < (1'h1)); forvar1257 = (forvar1257 + (1'h1)))
            begin
              reg1258 <= (($signed($signed((^~reg1055))) ?
                  $signed($unsigned((|reg1138))) : ((^~reg1175[(2'h3):(2'h3)]) ?
                      $signed((~&(8'ha4))) : (~&reg1175[(4'ha):(2'h2)]))) + (reg1070[(1'h1):(1'h1)] <= reg1179));
              reg1259 <= wire1229;
              reg1260 = ($signed((({reg1038, reg1258} ?
                      (forvar1257 ?
                          (7'h43) : reg1149) : {reg1011}) - reg1089[(4'ha):(3'h5)])) ?
                  ($signed(wire1231[(5'h11):(4'hd)]) != reg1197[(3'h7):(1'h0)]) : reg1117[(1'h1):(1'h1)]);
              reg1261 = $unsigned($unsigned(reg1244[(4'h8):(4'h8)]));
              reg1262 <= (8'ha1);
              reg1263 <= reg1076[(3'h4):(3'h4)];
              reg1264 = reg1236[(5'h14):(4'he)];
            end
          for (forvar1265 = (1'h0); (forvar1265 < (1'h1)); forvar1265 = (forvar1265 + (1'h1)))
            begin
              reg1266 <= ($signed((~^reg1221)) ?
                  (reg1089 ?
                      (((~|reg1183) <<< reg1225[(3'h6):(1'h0)]) ?
                          ({(8'h9c), forvar1257, reg1071} ?
                              {reg1053,
                                  reg1050,
                                  reg1227} : $signed(reg1094)) : reg1042) : {((reg1043 != reg1121) >> $signed(reg1093)),
                          reg1032}) : $signed((-reg1078)));
              reg1267 <= (~$signed($signed((~$signed(reg1066)))));
              reg1268 <= reg1012[(3'h4):(2'h2)];
              reg1269 <= ($signed(((&reg1152) ?
                      $unsigned(reg1149) : reg1245[(1'h1):(1'h1)])) ?
                  $unsigned(({(+reg1102),
                      (reg1106 && (8'hb1))} | ((reg1221 == reg1034) * reg1152))) : (!$signed((~&(wire1231 ?
                      wire1226 : reg1208)))));
            end
        end
      for (forvar1270 = (1'h0); (forvar1270 < (2'h3)); forvar1270 = (forvar1270 + (1'h1)))
        begin
          for (forvar1271 = (1'h0); (forvar1271 < (1'h1)); forvar1271 = (forvar1271 + (1'h1)))
            begin
              reg1272 <= (reg1053[(3'h6):(3'h5)] ?
                  reg1235 : {{reg1179, $unsigned(reg1244[(2'h3):(2'h2)])}});
              reg1273 = (!wire1007[(2'h2):(1'h1)]);
              reg1274 = $signed(((|{(reg1225 * (7'h43)),
                  (8'hb8),
                  {(8'ha6), (7'h52), forvar1232}}) || wire1010));
              reg1275 = reg1139[(4'hf):(4'hc)];
              reg1276 <= $unsigned($unsigned(forvar1257));
              reg1277 <= ({$signed(reg1155)} ?
                  {$signed(((~&reg1012) ? (reg1235 >>> (8'ha5)) : (^reg1170))),
                      ($signed(reg1088[(3'h6):(2'h2)]) ?
                          (+$signed((7'h54))) : $signed(reg1191))} : $signed(reg1219[(5'h1c):(5'h1a)]));
              reg1278 = reg1088;
            end
          reg1279 <= {({(^{(8'haf)})} ?
                  (((reg1273 > reg1055) ?
                          (reg1151 >> reg1155) : $unsigned(wire1231)) ?
                      $unsigned((reg1027 ^~ reg1070)) : (!(8'hbf))) : ((((7'h4a) ^ reg1118) + (|(8'h9f))) && wire1007)),
              (7'h47)};
          if ($unsigned(((!$signed((reg1027 ? reg1049 : reg1250))) ?
              $signed({(-reg1092)}) : (((wire1008 | reg1241) + (~|reg1102)) ?
                  reg1148 : $signed((8'ha3))))))
            begin
              reg1280 <= {$unsigned((reg1189 ^ $signed((~reg1219))))};
              reg1281 <= (8'hb2);
              reg1282 = (&$signed(reg1187[(4'h9):(1'h1)]));
              reg1283 = reg1106;
              reg1284 = ($signed((-wire1229[(4'h8):(3'h4)])) < $signed($unsigned(reg1167[(1'h1):(1'h1)])));
              reg1285 = ($signed({($unsigned(reg1266) | reg1112),
                      reg1284[(5'h15):(3'h4)],
                      {(reg1088 != reg1238), (~&reg1138)}}) ?
                  {$signed((!(~forvar1265))),
                      $unsigned((^reg1099[(1'h1):(1'h0)]))} : (&$unsigned((reg1234 >= reg1172))));
              reg1286 <= (reg1034 <= reg1193[(1'h1):(1'h1)]);
            end
          else
            begin
              reg1282 = (((~((reg1266 ? reg1089 : reg1207) ?
                  $signed(reg1208) : {reg1032})) || (reg1233[(4'hb):(1'h1)] ^ reg1124[(5'h15):(5'h15)])) > (((-reg1184) - reg1094[(3'h5):(2'h3)]) - $unsigned((8'hbf))));
              reg1286 <= (^($unsigned({reg1241}) ?
                  {reg1077[(5'h12):(5'h12)],
                      reg1278,
                      (reg1032 != reg1269)} : wire1229[(2'h3):(1'h1)]));
              reg1287 = reg1277[(4'h9):(3'h4)];
              reg1288 = (^~(reg1066[(1'h1):(1'h0)] ?
                  {reg1027[(1'h0):(1'h0)]} : {$unsigned($signed(reg1198)),
                      (forvar1243 ?
                          (reg1261 <<< reg1269) : (reg1136 ?
                              reg1027 : reg1283))}));
            end
          reg1289 <= reg1093[(5'h12):(4'ha)];
          if ((($signed({(reg1241 == reg1078),
                  ((8'haf) >= reg1255),
                  reg1165[(1'h1):(1'h0)]}) + $unsigned((8'hbe))) ?
              (^~(reg1161[(4'h8):(2'h3)] || (((8'hb3) ?
                  reg1087 : reg1188) > $signed(reg1219)))) : ((7'h56) ?
                  reg1088[(3'h4):(3'h4)] : (reg1016[(3'h5):(3'h4)] + (7'h4b)))))
            begin
              reg1290 = reg1183;
              reg1291 <= (~&reg1216);
              reg1292 <= (7'h57);
              reg1293 <= reg1282[(5'h13):(5'h12)];
            end
          else
            begin
              reg1290 = ($signed($signed((reg1025 + $signed(reg1148)))) ^ $unsigned($unsigned(reg1144[(5'h1e):(5'h1b)])));
              reg1291 <= ((^~($unsigned((8'hb8)) <<< $unsigned((wire1228 ?
                      (7'h47) : (8'ha9))))) ?
                  reg1194 : (^$signed((reg1032 | reg1118))));
              reg1292 <= {(~|({(wire1010 << reg1287), reg1175[(1'h1):(1'h0)]} ?
                      ($unsigned(reg1234) ?
                          ((7'h50) | (7'h41)) : $signed(reg1124)) : reg1159)),
                  $signed((+{{reg1283}}))};
              reg1294 = (7'h44);
              reg1295 = (8'hba);
              reg1296 = ((~&reg1249[(5'h15):(3'h7)]) <<< (reg1225[(3'h7):(3'h6)] * (-reg1285[(4'h9):(3'h7)])));
              reg1297 = (|reg1144[(4'h9):(4'h8)]);
            end
        end
      if (reg1204)
        begin
          reg1298 <= $signed(reg1269);
          reg1299 = $signed($unsigned(reg1191[(1'h0):(1'h0)]));
          reg1300 = (($unsigned($signed(reg1118[(5'h16):(4'hb)])) ~^ ((7'h4f) ^ $unsigned((7'h4a)))) & ($signed(((8'hb0) >= (reg1041 ?
                  reg1025 : reg1183))) ?
              reg1151[(3'h5):(2'h2)] : {reg1285[(1'h1):(1'h0)], reg1144}));
          reg1301 <= (((~^reg1187[(1'h0):(1'h0)]) ?
              reg1074[(3'h6):(2'h3)] : reg1293[(2'h2):(2'h2)]) << (reg1274 ?
              reg1155[(3'h6):(3'h4)] : {$unsigned(reg1207[(3'h6):(1'h1)]),
                  $unsigned($unsigned(reg1249))}));
          reg1302 <= reg1032;
          if ($signed((reg1193[(3'h4):(2'h3)] ?
              ($signed(reg1148) ?
                  $signed((&(7'h4a))) : ((reg1086 >> reg1236) ?
                      reg1183[(3'h5):(1'h0)] : wire1007[(1'h1):(1'h1)])) : $signed(reg1050))))
            begin
              reg1303 = reg1148[(4'ha):(4'ha)];
              reg1304 = (~^($unsigned(((^reg1124) ?
                  reg1077[(5'h19):(4'h8)] : $signed((7'h54)))) < reg1041[(2'h2):(1'h1)]));
              reg1305 = $unsigned($signed(($signed(reg1187) >>> wire1010)));
              reg1306 = ({reg1092[(4'he):(3'h6)],
                  $unsigned($signed(reg1198)),
                  $signed($signed((reg1289 ? reg1096 : reg1282)))} < {reg1236,
                  (reg1227[(1'h0):(1'h0)] == reg1139[(4'hd):(3'h6)])});
              reg1307 <= reg1303;
            end
          else
            begin
              reg1307 <= (~^(reg1298[(5'h18):(3'h6)] ?
                  $signed(((reg1011 <<< (8'hac)) ?
                      {reg1269, reg1055, reg1193} : {reg1161,
                          reg1077,
                          reg1258})) : $unsigned((((7'h52) - reg1267) ?
                      $unsigned(reg1238) : reg1094))));
              reg1308 <= reg1293[(3'h6):(3'h6)];
              reg1309 <= (($unsigned(($signed(reg1261) <<< (|reg1275))) ?
                  reg1093 : ({(&reg1050), $signed(reg1117)} ?
                      (reg1233[(3'h7):(3'h5)] <<< {reg1101}) : reg1127)) >> (reg1237[(4'h9):(2'h3)] ?
                  $unsigned(reg1136[(1'h1):(1'h0)]) : (+reg1086[(5'h10):(4'hf)])));
              reg1310 = reg1127[(3'h7):(3'h4)];
              reg1311 = $signed({(((reg1203 <= reg1158) & forvar1271[(3'h6):(2'h2)]) ?
                      (&(reg1077 && reg1025)) : $unsigned(reg1085[(5'h1a):(4'h8)])),
                  (|($unsigned(reg1206) ? $signed(reg1260) : (|(8'hba))))});
              reg1312 = $unsigned(reg1260[(1'h0):(1'h0)]);
            end
        end
      else
        begin
          reg1298 <= reg1172[(4'hc):(4'h9)];
          if ($unsigned(reg1294))
            begin
              reg1299 = {reg1284,
                  ((reg1225[(1'h0):(1'h0)] >> (!(reg1127 || reg1248))) ?
                      reg1130[(1'h0):(1'h0)] : $signed($signed($unsigned(reg1189))))};
            end
          else
            begin
              reg1301 <= ({reg1179[(4'hb):(1'h1)],
                  reg1260[(2'h3):(2'h2)],
                  $signed($signed($unsigned(reg1292)))} <= reg1145[(4'hd):(3'h4)]);
              reg1302 <= ($unsigned(reg1016[(5'h18):(3'h5)]) != reg1194);
              reg1303 = $signed({((-$signed(reg1277)) + $signed((reg1303 ?
                      (7'h47) : reg1167))),
                  ($unsigned(reg1296[(4'ha):(3'h5)]) ?
                      $signed((8'had)) : $unsigned($signed(reg1074))),
                  ((|reg1241) ?
                      $unsigned(reg1066) : ((reg1033 >>> reg1208) ?
                          (wire1009 ?
                              reg1198 : reg1015) : $unsigned(reg1038)))});
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg1236)
        begin
          if ((reg1241[(5'h10):(2'h3)] > reg1177))
            begin
              reg1313 <= {$unsigned($unsigned(((|reg1187) <= $unsigned(reg1246))))};
              reg1314 <= (^~$signed($unsigned(reg1313[(5'h12):(4'he)])));
              reg1315 <= $signed($signed(reg1133));
              reg1316 = (8'hae);
              reg1317 = (-reg1218[(4'hd):(1'h1)]);
            end
          else
            begin
              reg1316 = ({(((reg1048 ?
                      reg1238 : reg1289) >> $signed(reg1208)) ~^ (|(reg1197 ?
                      (8'hbb) : (7'h52)))),
                  {{(~|reg1259), (reg1308 ? reg1121 : (7'h45)), reg1272},
                      ((reg1152 <= reg1192) ?
                          {reg1198, (8'hbd), reg1138} : reg1033[(4'hf):(4'ha)]),
                      reg1267}} ~^ reg1096);
              reg1318 <= reg1101;
              reg1319 = (+$signed($signed(reg1011[(4'h8):(3'h4)])));
              reg1320 = $unsigned({reg1206[(5'h13):(4'hf)],
                  {(reg1307 * (reg1279 ^ (7'h57))),
                      reg1219[(5'h18):(4'hc)],
                      reg1096},
                  ($unsigned(reg1066) ?
                      $unsigned(((7'h49) ^ reg1187)) : $signed(((8'hb7) ?
                          reg1085 : (7'h4f))))});
              reg1321 <= reg1191;
              reg1322 <= $signed((~(7'h48)));
              reg1323 <= ((~((8'ha4) ^ {reg1142[(1'h0):(1'h0)]})) > (^~reg1236));
            end
          if (reg1320)
            begin
              reg1324 <= ((&(|reg1241)) ^ $unsigned(reg1013));
              reg1325 = $unsigned($unsigned({reg1124[(5'h1d):(5'h14)],
                  $unsigned((reg1318 ? reg1221 : reg1070))}));
              reg1326 = {(|(7'h53)),
                  $unsigned($signed(((reg1159 ? reg1276 : reg1042) ?
                      $unsigned(reg1136) : reg1179[(4'hb):(3'h7)])))};
            end
          else
            begin
              reg1325 = (7'h56);
              reg1326 = reg1124[(5'h13):(3'h5)];
            end
          if (wire1230[(5'h15):(4'hf)])
            begin
              reg1327 = (reg1074[(5'h16):(5'h10)] >> reg1025[(3'h5):(2'h3)]);
              reg1328 = reg1245[(3'h4):(2'h3)];
              reg1329 = {(~|(((+reg1030) ?
                      (reg1030 ?
                          reg1189 : wire1229) : reg1016[(5'h14):(4'h9)]) > $signed(reg1194)))};
              reg1330 = $signed((($signed((~&(8'haa))) <<< ((+reg1070) >> (reg1151 ?
                  reg1241 : reg1094))) * reg1193));
              reg1331 = $signed((($unsigned((~&reg1266)) <<< reg1324[(4'hb):(3'h7)]) ?
                  ($unsigned(reg1101) ?
                      ($signed(reg1208) ?
                          reg1309 : reg1152) : reg1118) : ((reg1052[(3'h5):(3'h5)] ?
                      (^(8'h9c)) : (reg1035 ?
                          reg1268 : reg1324)) * ($signed((8'h9c)) ?
                      $signed((8'ha2)) : $unsigned(reg1259)))));
            end
          else
            begin
              reg1327 = reg1314[(4'hd):(3'h5)];
            end
          reg1332 <= $signed(reg1025);
          reg1333 = ($unsigned($unsigned((~^reg1076[(1'h0):(1'h0)]))) ?
              (|$signed(reg1050)) : (~&reg1011));
          if (reg1093[(3'h5):(3'h5)])
            begin
              reg1334 <= ($unsigned({$unsigned($signed(reg1206))}) < $unsigned($signed(reg1279[(3'h5):(1'h1)])));
              reg1335 <= $signed($signed(wire1226));
              reg1336 <= (~|$unsigned({(~&$signed(reg1085)),
                  $signed((reg1096 ? reg1219 : reg1112))}));
            end
          else
            begin
              reg1334 <= $signed(((7'h54) - (-reg1146)));
            end
        end
      else
        begin
          if ($signed(reg1165))
            begin
              reg1313 <= (8'ha0);
              reg1314 <= reg1136[(3'h7):(2'h2)];
              reg1316 = (8'h9d);
            end
          else
            begin
              reg1313 <= reg1259[(2'h2):(2'h2)];
              reg1314 <= $signed(((-reg1121[(3'h7):(2'h3)]) ?
                  $signed(reg1038[(1'h1):(1'h1)]) : reg1237[(4'ha):(3'h5)]));
              reg1316 = ((reg1087 ?
                      ($unsigned(reg1170[(4'h9):(1'h1)]) | $unsigned(reg1258[(3'h7):(2'h3)])) : (+reg1087[(4'hb):(3'h7)])) ?
                  (((^(8'hbf)) ?
                          ((^~reg1218) ^ (7'h4f)) : reg1309[(3'h4):(2'h2)]) ?
                      $signed($unsigned(reg1314)) : ({(reg1015 ?
                              reg1099 : reg1219),
                          reg1066,
                          (reg1207 ?
                              (7'h48) : reg1188)} >= reg1331)) : (7'h41));
              reg1317 = ({$signed((~|$signed(reg1328)))} == reg1301[(2'h3):(1'h0)]);
              reg1318 <= {(reg1309 ?
                      reg1085 : ({$unsigned(reg1313),
                          reg1011} ~^ {(!(7'h42))})),
                  (reg1203 | ((-reg1245) ?
                      $signed({reg1049,
                          reg1237,
                          reg1025}) : ((reg1216 && reg1194) ^ reg1302[(4'hc):(3'h5)])))};
              reg1321 <= $unsigned($unsigned(reg1222[(5'h12):(4'hf)]));
            end
          if (($unsigned($unsigned(((reg1187 ^~ reg1277) << reg1099))) * $unsigned(($unsigned($signed(reg1133)) << reg1315[(2'h3):(1'h1)]))))
            begin
              reg1325 = (((reg1262[(5'h15):(5'h15)] ?
                  reg1207[(1'h0):(1'h0)] : $unsigned((~&reg1076))) << $signed(reg1281[(4'hd):(3'h7)])) & reg1126[(4'ha):(2'h2)]);
              reg1326 = reg1291[(4'h8):(3'h5)];
              reg1332 <= $signed(reg1262);
              reg1333 = $signed($signed($unsigned($signed((reg1301 ?
                  reg1117 : reg1316)))));
              reg1337 = reg1025;
              reg1338 <= reg1197;
              reg1339 <= {reg1262[(5'h11):(5'h10)]};
            end
          else
            begin
              reg1322 <= reg1126[(3'h7):(2'h2)];
              reg1325 = $unsigned(reg1237);
            end
          reg1340 = reg1151;
          reg1341 = (-(7'h4d));
          reg1342 <= $signed(reg1333);
        end
      if (((-$signed((!(reg1158 & reg1145)))) ?
          $unsigned((($unsigned(reg1280) ?
              (reg1188 ^ reg1331) : ((8'ha6) - reg1158)) && ($signed(reg1326) ?
              (7'h43) : (&reg1043)))) : {(reg1142[(1'h0):(1'h0)] ?
                  reg1030[(1'h1):(1'h1)] : (wire1226 <= reg1193[(2'h2):(2'h2)])),
              reg1175,
              reg1326[(4'he):(3'h7)]}))
        begin
          for (forvar1343 = (1'h0); (forvar1343 < (3'h6)); forvar1343 = (forvar1343 + (1'h1)))
            begin
              reg1344 <= wire1007[(2'h2):(1'h1)];
              reg1345 = ($unsigned(reg1033[(4'hd):(1'h0)]) ?
                  reg1076[(2'h2):(1'h1)] : $signed($unsigned($signed((reg1056 ?
                      reg1197 : reg1092)))));
              reg1346 = (-$signed(($unsigned(((8'hb5) < reg1122)) ?
                  reg1102 : ((reg1012 || (8'ha6)) ?
                      (reg1241 ? reg1308 : (8'hbd)) : (reg1344 <<< (7'h54))))));
              reg1347 = (reg1189[(1'h0):(1'h0)] ?
                  $signed((reg1151 ?
                      {$unsigned(reg1146)} : (&(8'ha6)))) : $signed(reg1338[(4'h9):(3'h4)]));
              reg1348 = (reg1117[(3'h6):(1'h0)] ?
                  (!reg1027[(1'h1):(1'h0)]) : reg1144[(2'h2):(2'h2)]);
              reg1349 = $unsigned(reg1034);
            end
          reg1350 = (({reg1102} ?
                  ($signed((reg1071 ? reg1329 : (8'hbc))) ?
                      (~|(reg1179 ^ (7'h48))) : $signed($unsigned(reg1088))) : reg1193) ?
              (reg1041[(3'h6):(2'h3)] << $signed(((+reg1319) >>> $unsigned(reg1246)))) : (!$unsigned($unsigned(reg1340[(3'h5):(1'h0)]))));
          reg1351 = ((&reg1048) ?
              ((($signed((8'hba)) ? (+(8'hb7)) : (7'h45)) == $signed({reg1158,
                  (8'haa),
                  reg1112})) <<< (((reg1332 && reg1172) & reg1142[(1'h0):(1'h0)]) ?
                  reg1152 : (~|$signed(reg1222)))) : (~&(~&$signed(reg1013[(2'h2):(1'h1)]))));
          for (forvar1352 = (1'h0); (forvar1352 < (2'h3)); forvar1352 = (forvar1352 + (1'h1)))
            begin
              reg1353 = (^($unsigned(reg1238[(3'h6):(2'h2)]) ?
                  $unsigned($unsigned((^~reg1331))) : reg1237));
            end
          for (forvar1354 = (1'h0); (forvar1354 < (1'h0)); forvar1354 = (forvar1354 + (1'h1)))
            begin
              reg1355 <= (~|(reg1263 ?
                  (8'hb9) : $unsigned({reg1235[(5'h13):(5'h13)],
                      $signed(reg1112),
                      $signed(reg1219)})));
              reg1356 = ((reg1326 ?
                  (~&((reg1218 ? reg1155 : reg1145) ?
                      $signed((8'hb8)) : reg1301)) : reg1183[(4'h9):(3'h7)]) > $signed(((^$signed(reg1179)) ?
                  ((reg1316 ? (8'hbf) : reg1077) ?
                      reg1351 : (|reg1086)) : (wire1231 > reg1337[(3'h6):(3'h6)]))));
              reg1357 <= (reg1175[(3'h5):(3'h5)] < $unsigned({{reg1034[(3'h4):(2'h2)],
                      reg1086}}));
              reg1358 <= $unsigned((((forvar1352[(4'hd):(4'ha)] != reg1293) >> ({reg1353,
                  reg1238,
                  reg1156} >= (~^reg1333))) && $signed($signed((reg1323 ?
                  reg1189 : (7'h53))))));
              reg1359 <= (~|((~^$signed((~reg1015))) >> (+($signed(reg1222) ?
                  reg1013 : $unsigned(reg1012)))));
            end
          reg1360 <= reg1094[(2'h2):(2'h2)];
          reg1361 <= (^~$signed(reg1329[(5'h16):(5'h12)]));
        end
      else
        begin
          reg1343 = (~&(7'h48));
          reg1345 = $signed(((reg1149 | (reg1013[(5'h10):(4'hf)] ^ reg1326[(4'he):(4'hd)])) != {reg1112[(2'h3):(2'h3)]}));
          reg1346 = $unsigned(reg1198[(4'hb):(3'h6)]);
          if ((8'hb4))
            begin
              reg1352 <= ((~&reg1356) ?
                  ((reg1049[(2'h2):(2'h2)] ?
                      {(reg1035 * reg1251)} : $signed((reg1055 ?
                          reg1089 : (7'h50)))) ~^ (reg1344[(5'h16):(4'hf)] ?
                      {{reg1187, reg1198}} : (~|(reg1093 ?
                          (8'h9f) : reg1349)))) : reg1032);
              reg1353 = reg1307;
              reg1354 = reg1094[(4'h9):(4'h9)];
            end
          else
            begin
              reg1347 = (reg1350 < $signed($unsigned(reg1167)));
              reg1348 = ($unsigned((reg1193 ~^ reg1321[(1'h0):(1'h0)])) > reg1070[(3'h4):(2'h3)]);
              reg1352 <= reg1034;
              reg1355 <= ((wire1007 <<< ((~^(reg1092 ?
                  reg1055 : wire1228)) * wire1231[(2'h2):(1'h0)])) > (-($signed(reg1218) ?
                  $unsigned($signed((7'h4a))) : reg1272)));
              reg1357 <= ($signed((reg1100 ?
                  ({reg1360,
                      reg1359,
                      reg1245} >> (8'hae)) : (+$unsigned(reg1038)))) * (&reg1319[(3'h6):(3'h6)]));
              reg1358 <= reg1035[(4'hd):(2'h2)];
            end
        end
      reg1362 = $signed((~(|$unsigned($unsigned(reg1361)))));
      reg1363 <= (&($unsigned(((reg1236 ? (8'hae) : reg1238) ?
              $signed((7'h57)) : $unsigned(reg1191))) ?
          reg1227 : (reg1193[(1'h1):(1'h0)] ?
              reg1041 : ($signed(reg1334) | (&wire1229)))));
    end
  assign wire1364 = {(($signed($unsigned(reg1099)) ?
                            $unsigned(reg1025[(3'h4):(2'h3)]) : (((7'h41) ?
                                    reg1336 : reg1192) ?
                                $signed(reg1165) : (~(7'h4f)))) && (reg1269[(5'h18):(4'ha)] ^~ $unsigned((^wire1228)))),
                        (~|reg1269[(4'he):(1'h1)]),
                        (~^reg1145)};
  always
    @(posedge clk) begin
      if ((~&reg1122))
        begin
          for (forvar1365 = (1'h0); (forvar1365 < (1'h1)); forvar1365 = (forvar1365 + (1'h1)))
            begin
              reg1366 <= ((reg1298 & (8'h9c)) && (!{($unsigned(reg1070) < (reg1245 ?
                      reg1124 : reg1293)),
                  reg1156[(2'h3):(2'h2)],
                  reg1301[(3'h5):(3'h4)]}));
              reg1367 <= (reg1117 & reg1344);
              reg1368 <= (^~$unsigned(reg1269));
              reg1369 = reg1301[(3'h4):(2'h2)];
              reg1370 <= ((~^$signed($signed((^wire1006)))) >> (!((^~$signed(reg1194)) << reg1155[(2'h3):(2'h2)])));
            end
          reg1371 = (((((~|reg1279) << reg1313[(1'h0):(1'h0)]) ?
                  reg1161[(4'h8):(1'h1)] : $unsigned((reg1335 ?
                      (8'hb6) : reg1015))) ?
              reg1049 : reg1352) < (($signed((reg1191 ?
              reg1077 : reg1189)) << reg1052) | wire1082));
          if ({$unsigned(reg1122)})
            begin
              reg1372 <= $unsigned((reg1188[(1'h1):(1'h0)] <<< (reg1191 ?
                  reg1118 : $signed({reg1358, reg1206}))));
              reg1373 <= (~^$unsigned($signed((8'hac))));
              reg1374 = $signed((~|$signed({$signed(wire1228)})));
              reg1375 <= (reg1259 ?
                  {(~|$unsigned($unsigned(reg1096))),
                      reg1289[(1'h1):(1'h0)]} : (~$unsigned(reg1043[(3'h7):(2'h3)])));
            end
          else
            begin
              reg1374 = ({((~(^reg1324)) ?
                      $unsigned(((7'h54) ?
                          reg1066 : (8'ha7))) : reg1203[(1'h1):(1'h0)])} * (((reg1361 ?
                  reg1191 : $unsigned(reg1144)) | (~|$unsigned(reg1139))) * reg1197));
              reg1376 = reg1204;
              reg1377 = (~|{(~$signed($unsigned(reg1094))),
                  reg1148,
                  {{$unsigned(reg1136)},
                      {reg1259, (reg1369 >> (7'h42)), $unsigned(reg1124)},
                      reg1055}});
              reg1378 = $signed($signed((+$unsigned((reg1074 ?
                  reg1361 : reg1334)))));
              reg1379 = (-reg1377);
              reg1380 <= $unsigned(reg1086[(2'h2):(1'h1)]);
              reg1381 <= ({(((reg1159 | reg1102) ?
                              (8'hb6) : (reg1298 ? reg1268 : (8'h9f))) ?
                          ((|reg1086) ?
                              reg1204 : (reg1219 == (8'haf))) : ((forvar1365 ?
                              reg1043 : reg1259) >= (reg1133 * reg1100))),
                      reg1188[(1'h1):(1'h0)]} ?
                  reg1196 : reg1218);
            end
          reg1382 <= reg1339[(3'h5):(3'h5)];
          reg1383 = {(|{((reg1237 <<< reg1101) ?
                      ((7'h56) >>> reg1136) : (+reg1204))}),
              ({((reg1266 - reg1042) & reg1118[(5'h1c):(5'h16)])} ?
                  (((reg1301 ? reg1368 : reg1357) ?
                          (reg1093 <= reg1106) : (reg1245 <= reg1172)) ?
                      ((|reg1074) - (reg1142 ?
                          reg1359 : reg1197)) : ((^~reg1161) ?
                          (reg1216 > (8'ha7)) : reg1193[(3'h7):(3'h7)])) : reg1381)};
          for (forvar1384 = (1'h0); (forvar1384 < (3'h4)); forvar1384 = (forvar1384 + (1'h1)))
            begin
              reg1385 = (+$unsigned($signed(reg1379)));
              reg1386 <= reg1237[(2'h3):(2'h2)];
              reg1387 = $signed((reg1246[(3'h7):(1'h1)] ?
                  wire1230[(3'h4):(1'h1)] : ($signed((~^reg1378)) ?
                      reg1149[(5'h13):(3'h4)] : ($signed((8'hbe)) >> (reg1286 ?
                          reg1218 : (7'h4d))))));
              reg1388 <= (((~&(~|$unsigned(reg1197))) == reg1334[(2'h2):(1'h0)]) ?
                  reg1363[(4'ha):(1'h1)] : $signed(($unsigned((^~wire1226)) << (reg1279[(1'h1):(1'h0)] + reg1142[(2'h2):(2'h2)]))));
              reg1389 = ((($signed((reg1106 ? reg1266 : reg1158)) != ((reg1267 ?
                          reg1314 : (8'h9c)) ?
                      reg1197 : $unsigned(reg1048))) && $signed(reg1358)) ?
                  reg1156 : reg1286[(4'hb):(4'hb)]);
              reg1390 <= (reg1089[(5'h10):(3'h5)] ?
                  reg1241 : reg1361[(1'h1):(1'h0)]);
              reg1391 = (~reg1289[(1'h1):(1'h1)]);
            end
          reg1392 = $unsigned(wire1230[(5'h11):(5'h11)]);
        end
      else
        begin
          reg1365 <= reg1380;
          for (forvar1366 = (1'h0); (forvar1366 < (1'h1)); forvar1366 = (forvar1366 + (1'h1)))
            begin
              reg1369 = reg1251[(2'h3):(1'h0)];
              reg1371 = $signed((&reg1049));
              reg1372 <= (!$unsigned(reg1314));
              reg1374 = reg1315[(3'h5):(1'h0)];
            end
          reg1375 <= (($signed(((&forvar1365) ? $signed(reg1100) : {reg1159})) ?
              {reg1126[(3'h4):(2'h3)],
                  (7'h4c)} : reg1386[(4'h8):(1'h0)]) & wire1226[(5'h12):(4'he)]);
        end
      for (forvar1393 = (1'h0); (forvar1393 < (3'h4)); forvar1393 = (forvar1393 + (1'h1)))
        begin
          for (forvar1394 = (1'h0); (forvar1394 < (2'h2)); forvar1394 = (forvar1394 + (1'h1)))
            begin
              reg1395 <= $unsigned($unsigned(reg1177));
            end
          reg1396 = $unsigned((^$unsigned(reg1070[(4'hf):(4'ha)])));
          for (forvar1397 = (1'h0); (forvar1397 < (1'h1)); forvar1397 = (forvar1397 + (1'h1)))
            begin
              reg1398 = (({(reg1263[(5'h14):(4'hf)] ?
                              (~&reg1258) : (wire1007 ? wire1230 : (8'hb6)))} ?
                      $unsigned(((reg1142 || wire1228) ?
                          $signed(reg1204) : $signed(reg1070))) : $signed((reg1339[(2'h3):(2'h2)] ?
                          (~|reg1374) : (~reg1184)))) ?
                  (((reg1155 > (reg1179 <<< (8'hb6))) <<< reg1389) ?
                      {$signed((reg1259 ^~ (7'h54))),
                          (!{reg1086, reg1307}),
                          reg1292} : ((-reg1193) ?
                          (^~((7'h4a) ?
                              wire1006 : reg1050)) : reg1298[(3'h5):(2'h2)])) : ({{reg1194,
                          $unsigned(reg1396)}} ^ reg1267[(4'ha):(2'h2)]));
              reg1399 = reg1388[(4'ha):(1'h1)];
              reg1400 <= $unsigned((reg1382 ?
                  $unsigned($signed($signed(reg1352))) : wire1231));
              reg1401 <= $signed(reg1122[(4'h9):(2'h3)]);
              reg1402 <= $signed($signed(wire1230[(4'h9):(2'h2)]));
            end
        end
    end
endmodule