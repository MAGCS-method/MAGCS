(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param1025 = {(8'hb2), ((({(8'hb8), (8'hb7)} < (~(7'h41))) ? {((7'h40) ? (8'h9c) : (8'haf))} : {((7'h4a) ? (8'hb7) : (8'hb2))}) ? ({((8'h9f) ? (8'ha5) : (8'hae))} || (~(&(8'ha2)))) : ((8'hb0) & (((8'hb2) - (7'h40)) ? (|(7'h44)) : ((8'h9d) ^~ (8'ha9)))))}, 
parameter param1026 = (param1025 ? (7'h44) : (|{(-(param1025 <= param1025))})))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h137):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire0;
  input wire [(5'h18):(1'h0)] wire1;
  input wire signed [(5'h10):(1'h0)] wire2;
  input wire signed [(3'h7):(1'h0)] wire3;
  wire signed [(2'h2):(1'h0)] wire1024;
  wire [(5'h17):(1'h0)] wire1023;
  wire [(5'h14):(1'h0)] wire22;
  wire [(5'h14):(1'h0)] wire1021;
  reg signed [(2'h3):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg18 = (1'h0);
  reg [(5'h17):(1'h0)] reg13 = (1'h0);
  reg [(4'hb):(1'h0)] reg11 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg21 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar16 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar14 = (1'h0);
  reg [(5'h14):(1'h0)] reg12 = (1'h0);
  reg [(5'h10):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar9 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg7 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4 = (1'h0);
  assign y = {wire1024,
                 wire1023,
                 wire22,
                 wire1021,
                 reg19,
                 reg18,
                 reg13,
                 reg11,
                 reg6,
                 reg21,
                 reg20,
                 reg17,
                 forvar16,
                 reg15,
                 forvar14,
                 reg12,
                 reg10,
                 forvar9,
                 reg8,
                 reg7,
                 reg5,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (3'h4)); forvar4 = (forvar4 + (1'h1)))
        begin
          if ((wire2[(4'hd):(3'h5)] != ((~^{wire1,
              (wire3 == wire1)}) & (({wire1} + ((8'hb8) ? (8'hb5) : wire3)) ?
              (&$signed(forvar4)) : wire3))))
            begin
              reg5 = $signed($unsigned({(((7'h40) ? wire3 : wire2) ?
                      {forvar4, forvar4} : (wire2 ? wire1 : wire0)),
                  ((wire2 ? wire0 : wire1) > (wire2 ? (8'hb0) : forvar4))}));
              reg6 <= $unsigned((^forvar4[(1'h1):(1'h0)]));
              reg7 = $signed($signed({(|(!forvar4)),
                  {forvar4, (wire0 ? forvar4 : reg6)}}));
              reg8 = (^(forvar4 ?
                  wire2 : ($unsigned((reg7 > forvar4)) || $signed((wire0 < wire1)))));
            end
          else
            begin
              reg5 = (~&($signed((((8'hb8) ? reg6 : (7'h42)) == {(8'h9d),
                      reg6})) ?
                  (~|reg6) : $signed(wire2)));
              reg6 <= (~|$signed(wire1[(4'he):(4'h8)]));
            end
          for (forvar9 = (1'h0); (forvar9 < (1'h0)); forvar9 = (forvar9 + (1'h1)))
            begin
              reg10 = wire2;
              reg11 <= $unsigned(wire3);
            end
          reg12 = wire0[(3'h4):(3'h4)];
          reg13 <= reg12;
          for (forvar14 = (1'h0); (forvar14 < (3'h4)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 = ($unsigned(wire1) + $signed(($signed($unsigned(reg11)) ?
                  forvar4 : ($unsigned(wire0) ?
                      $signed(forvar4) : (reg5 >>> wire3)))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar16 = (1'h0); (forvar16 < (2'h3)); forvar16 = (forvar16 + (1'h1)))
        begin
          reg17 = $signed((~&$unsigned(wire1[(4'hd):(4'hb)])));
          reg18 <= $signed($signed((forvar16 - $unsigned($signed(forvar16)))));
        end
      reg19 <= ($signed($signed(wire2[(4'ha):(3'h4)])) ?
          reg17 : (wire2 ?
              (($signed(wire1) > {wire2}) ^~ (-forvar16[(4'h8):(3'h4)])) : (~$unsigned((8'h9d)))));
    end
  always
    @(posedge clk) begin
      reg20 = {((8'h9d) ?
              wire1[(5'h11):(5'h11)] : ((reg13 ?
                  reg19[(1'h1):(1'h0)] : (8'ha4)) << {(reg19 >= reg6),
                  {reg6}}))};
      reg21 = reg13[(3'h4):(2'h3)];
    end
  assign wire22 = (($unsigned({(~&wire0)}) >> reg18[(3'h7):(3'h7)]) | (8'hb2));
  module23 #() modinst1022 (wire1021, clk, wire22, wire2, reg13, wire0, reg11);
  assign wire1023 = $unsigned(((8'had) == {(((8'hba) ?
                            wire1021 : wire3) ^~ wire2[(2'h3):(1'h1)])}));
  assign wire1024 = ((reg6 ~^ (~^(^{reg11,
                        (8'ha0)}))) || (wire0[(4'hb):(2'h2)] ?
                        ($signed((wire22 ? wire2 : wire1023)) ?
                            (reg19 ?
                                (wire22 ?
                                    wire1023 : (8'ha3)) : wire3) : (8'hb2)) : {$signed((reg19 ?
                                (8'ha8) : wire22)),
                            wire1021[(4'hf):(1'h1)]}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module23  (y, clk, wire28, wire27, wire26, wire25, wire24);
  output wire [(32'h6b0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire28;
  input wire [(4'hf):(1'h0)] wire27;
  input wire signed [(5'h11):(1'h0)] wire26;
  input wire [(5'h15):(1'h0)] wire25;
  input wire [(4'hb):(1'h0)] wire24;
  wire [(5'h11):(1'h0)] wire956;
  wire signed [(5'h15):(1'h0)] wire955;
  wire signed [(4'he):(1'h0)] wire922;
  wire signed [(5'h13):(1'h0)] wire921;
  wire [(4'hc):(1'h0)] wire919;
  wire signed [(5'h15):(1'h0)] wire243;
  wire [(3'h6):(1'h0)] wire241;
  reg [(4'hb):(1'h0)] reg1015 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1014 = (1'h0);
  reg [(4'he):(1'h0)] reg1013 = (1'h0);
  reg [(5'h14):(1'h0)] reg1008 = (1'h0);
  reg [(5'h18):(1'h0)] reg1006 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1004 = (1'h0);
  reg [(4'hb):(1'h0)] reg1001 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1000 = (1'h0);
  reg [(3'h7):(1'h0)] reg999 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg996 = (1'h0);
  reg [(5'h16):(1'h0)] reg995 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg993 = (1'h0);
  reg [(5'h11):(1'h0)] reg992 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg990 = (1'h0);
  reg [(2'h3):(1'h0)] reg986 = (1'h0);
  reg [(4'hb):(1'h0)] reg976 = (1'h0);
  reg [(5'h16):(1'h0)] reg974 = (1'h0);
  reg [(4'he):(1'h0)] reg971 = (1'h0);
  reg [(5'h15):(1'h0)] reg969 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg968 = (1'h0);
  reg [(2'h3):(1'h0)] reg961 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg958 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg954 = (1'h0);
  reg [(5'h11):(1'h0)] reg953 = (1'h0);
  reg [(3'h5):(1'h0)] reg949 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg948 = (1'h0);
  reg [(4'he):(1'h0)] reg943 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg938 = (1'h0);
  reg [(4'h9):(1'h0)] reg934 = (1'h0);
  reg [(3'h7):(1'h0)] reg933 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg931 = (1'h0);
  reg [(4'hb):(1'h0)] reg930 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg929 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg928 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg924 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg54 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg53 = (1'h0);
  reg [(3'h7):(1'h0)] reg51 = (1'h0);
  reg [(4'h8):(1'h0)] reg48 = (1'h0);
  reg [(3'h7):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg46 = (1'h0);
  reg [(4'hd):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg39 = (1'h0);
  reg [(5'h12):(1'h0)] reg38 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg37 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg33 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg31 = (1'h0);
  reg [(5'h11):(1'h0)] reg30 = (1'h0);
  reg [(4'ha):(1'h0)] reg29 = (1'h0);
  reg [(4'hd):(1'h0)] reg1020 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1019 = (1'h0);
  reg [(4'hf):(1'h0)] reg1018 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1015 = (1'h0);
  reg [(4'he):(1'h0)] reg1017 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1016 = (1'h0);
  reg [(2'h3):(1'h0)] reg1012 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1011 = (1'h0);
  reg [(5'h13):(1'h0)] reg1010 = (1'h0);
  reg [(3'h5):(1'h0)] reg1009 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1007 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1005 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1003 = (1'h0);
  reg [(4'h8):(1'h0)] reg1002 = (1'h0);
  reg [(4'ha):(1'h0)] forvar995 = (1'h0);
  reg [(5'h13):(1'h0)] reg998 = (1'h0);
  reg [(2'h2):(1'h0)] reg997 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg994 = (1'h0);
  reg [(3'h5):(1'h0)] reg991 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg989 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg988 = (1'h0);
  reg [(5'h11):(1'h0)] forvar987 = (1'h0);
  reg [(4'he):(1'h0)] reg985 = (1'h0);
  reg signed [(4'he):(1'h0)] reg984 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg983 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar982 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg981 = (1'h0);
  reg [(4'h9):(1'h0)] reg980 = (1'h0);
  reg [(3'h4):(1'h0)] reg979 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg978 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg977 = (1'h0);
  reg [(5'h14):(1'h0)] forvar975 = (1'h0);
  reg [(5'h14):(1'h0)] reg973 = (1'h0);
  reg [(3'h4):(1'h0)] reg972 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar970 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar967 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar966 = (1'h0);
  reg [(4'he):(1'h0)] reg965 = (1'h0);
  reg [(3'h4):(1'h0)] reg964 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg963 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg962 = (1'h0);
  reg [(5'h12):(1'h0)] reg959 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar958 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg960 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar959 = (1'h0);
  reg [(5'h17):(1'h0)] reg957 = (1'h0);
  reg [(4'h9):(1'h0)] reg952 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg951 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg950 = (1'h0);
  reg [(4'ha):(1'h0)] reg947 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg946 = (1'h0);
  reg [(4'hf):(1'h0)] forvar945 = (1'h0);
  reg [(5'h15):(1'h0)] forvar944 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg942 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg941 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg940 = (1'h0);
  reg [(5'h15):(1'h0)] reg939 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg937 = (1'h0);
  reg [(5'h18):(1'h0)] reg936 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg935 = (1'h0);
  reg [(4'he):(1'h0)] reg932 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg927 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg926 = (1'h0);
  reg [(5'h11):(1'h0)] reg925 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar924 = (1'h0);
  reg [(3'h4):(1'h0)] reg52 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg50 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg49 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg45 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg36 = (1'h0);
  reg [(4'he):(1'h0)] reg35 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg34 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar32 = (1'h0);
  assign y = {wire956,
                 wire955,
                 wire922,
                 wire921,
                 wire919,
                 wire243,
                 wire241,
                 reg1015,
                 reg1014,
                 reg1013,
                 reg1008,
                 reg1006,
                 reg1004,
                 reg1001,
                 reg1000,
                 reg999,
                 reg996,
                 reg995,
                 reg993,
                 reg992,
                 reg990,
                 reg986,
                 reg976,
                 reg974,
                 reg971,
                 reg969,
                 reg968,
                 reg961,
                 reg958,
                 reg954,
                 reg953,
                 reg949,
                 reg948,
                 reg943,
                 reg938,
                 reg934,
                 reg933,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 reg924,
                 reg54,
                 reg53,
                 reg51,
                 reg48,
                 reg47,
                 reg46,
                 reg44,
                 reg42,
                 reg41,
                 reg39,
                 reg38,
                 reg37,
                 reg33,
                 reg31,
                 reg30,
                 reg29,
                 reg1020,
                 reg1019,
                 reg1018,
                 forvar1015,
                 reg1017,
                 reg1016,
                 reg1012,
                 reg1011,
                 reg1010,
                 reg1009,
                 reg1007,
                 reg1005,
                 reg1003,
                 reg1002,
                 forvar995,
                 reg998,
                 reg997,
                 reg994,
                 reg991,
                 reg989,
                 reg988,
                 forvar987,
                 reg985,
                 reg984,
                 reg983,
                 forvar982,
                 reg981,
                 reg980,
                 reg979,
                 reg978,
                 reg977,
                 forvar975,
                 reg973,
                 reg972,
                 forvar970,
                 forvar967,
                 forvar966,
                 reg965,
                 reg964,
                 reg963,
                 reg962,
                 reg959,
                 forvar958,
                 reg960,
                 forvar959,
                 reg957,
                 reg952,
                 reg951,
                 reg950,
                 reg947,
                 reg946,
                 forvar945,
                 forvar944,
                 reg942,
                 reg941,
                 reg940,
                 reg939,
                 reg937,
                 reg936,
                 reg935,
                 reg932,
                 reg927,
                 reg926,
                 reg925,
                 forvar924,
                 reg52,
                 reg50,
                 reg49,
                 reg45,
                 reg43,
                 reg40,
                 reg36,
                 reg35,
                 reg32,
                 reg34,
                 forvar32,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ({($signed($unsigned(wire24)) ?
              wire27[(4'h9):(1'h1)] : $unsigned(((+(8'h9f)) ?
                  $unsigned(wire28) : ((8'hb5) - wire27))))})
        begin
          reg29 <= (&{$signed(wire27)});
          reg30 <= $unsigned(($signed((|wire27[(3'h5):(3'h5)])) ?
              (((!wire25) ?
                  (wire28 == wire28) : {wire26}) > wire28[(1'h0):(1'h0)]) : reg29));
          reg31 <= ($signed((reg30 ?
                  {$signed(reg29),
                      (wire27 ?
                          (8'hbf) : wire28)} : $unsigned($signed(wire24)))) ?
              (reg29 ^~ (&wire24[(1'h1):(1'h1)])) : wire28[(5'h13):(4'hf)]);
          for (forvar32 = (1'h0); (forvar32 < (1'h0)); forvar32 = (forvar32 + (1'h1)))
            begin
              reg33 <= wire26[(4'ha):(3'h4)];
            end
          reg34 = (forvar32[(4'hf):(4'hc)] ?
              (~&wire25[(2'h3):(2'h3)]) : ($signed(wire28) ?
                  wire28 : ((forvar32[(5'h17):(3'h5)] ?
                          ((8'ha4) & (8'hbd)) : (reg29 ? forvar32 : wire27)) ?
                      wire27[(4'h8):(2'h3)] : $signed((+wire28)))));
        end
      else
        begin
          if ({(^~$signed(wire24))})
            begin
              reg32 = (wire27[(4'ha):(4'h9)] ^ $unsigned($unsigned($signed({reg29}))));
              reg33 <= $signed(reg29[(1'h1):(1'h0)]);
              reg34 = (~^((reg30[(2'h3):(2'h2)] & $signed((^wire25))) << (!$signed($signed(reg29)))));
            end
          else
            begin
              reg32 = (reg34 ?
                  reg29[(4'h9):(3'h6)] : ((&reg30) ?
                      $signed(forvar32[(2'h2):(2'h2)]) : (^~$unsigned($unsigned(wire26)))));
              reg34 = (reg29 ~^ reg34);
              reg35 = ((reg34[(5'h10):(1'h0)] && wire27[(4'h9):(1'h1)]) ?
                  (wire28[(1'h0):(1'h0)] ?
                      wire24[(2'h3):(2'h2)] : ({reg32[(1'h0):(1'h0)],
                              {wire24, wire27}} ?
                          forvar32 : $signed((8'hb5)))) : reg29);
              reg36 = $signed(((-reg29) ~^ $unsigned($unsigned(((7'h4a) ?
                  wire26 : reg35)))));
              reg37 <= (8'ha9);
            end
          if ((~^$unsigned(reg37[(1'h1):(1'h1)])))
            begin
              reg38 <= {reg33};
              reg39 <= reg30[(1'h1):(1'h0)];
            end
          else
            begin
              reg38 <= $unsigned(((((~&(8'ha8)) ?
                  wire26 : ((8'h9d) ? reg29 : reg33)) + reg31) ^ (~(8'h9d))));
              reg39 <= ($signed($signed($unsigned((~&reg38)))) ?
                  (~(8'ha9)) : $signed($signed((+(reg38 != reg30)))));
              reg40 = $unsigned($unsigned(reg30[(2'h2):(1'h1)]));
              reg41 <= {(reg37[(1'h1):(1'h1)] ^~ {((reg36 ? reg34 : reg34) ?
                          (reg40 ? reg33 : reg32) : {(8'ha1)}),
                      $signed(reg38)})};
              reg42 <= (^~(-reg37));
            end
          if (((((&reg29) != {$signed(reg35), (reg42 ? reg42 : wire26)}) ?
                  $signed(reg40) : (reg33 ?
                      $signed((~|(8'hba))) : $unsigned(reg37))) ?
              ($unsigned({{reg36, reg42}, $signed(reg39)}) ?
                  {$unsigned((&wire24)),
                      reg29} : $signed($signed($unsigned(reg36)))) : $unsigned($signed(forvar32))))
            begin
              reg43 = (^$signed((^~(reg42[(2'h3):(2'h3)] ?
                  ((8'ha8) <<< reg34) : $unsigned(reg38)))));
              reg44 <= $unsigned((7'h40));
              reg45 = ((((~(reg44 ? (8'ha3) : reg39)) ?
                      ((reg30 ? (8'ha2) : reg31) < $signed(reg41)) : reg29) ?
                  reg33 : reg33[(3'h6):(1'h0)]) - ({$unsigned($unsigned(reg40))} ?
                  wire28[(1'h0):(1'h0)] : ({(reg40 ? (8'hb8) : (8'haa)),
                          reg34} ?
                      ((reg37 < reg40) == wire26[(4'hd):(3'h7)]) : reg43)));
              reg46 <= ($signed((&(!reg34[(5'h10):(5'h10)]))) > reg40);
              reg47 <= (&(8'haf));
            end
          else
            begin
              reg44 <= (({((forvar32 ? reg30 : reg39) ~^ reg44)} ?
                      $unsigned(($signed(wire24) ?
                          wire28 : (^~reg33))) : reg39[(1'h0):(1'h0)]) ?
                  $unsigned(((~&$signed(wire24)) ?
                      $signed(((7'h45) && reg42)) : {(reg36 ? (8'had) : reg34),
                          (wire28 ?
                              wire26 : forvar32)})) : wire26[(4'hd):(3'h4)]);
              reg45 = $signed(($unsigned($signed($unsigned(wire25))) ?
                  $signed((~^reg34[(4'hd):(4'h8)])) : reg46));
            end
          if ((($signed($signed((wire28 <<< reg41))) * $signed($signed(wire27[(3'h4):(2'h3)]))) ?
              reg43 : {(^({(8'h9d), reg40} ~^ reg41)), reg38}))
            begin
              reg48 <= ($signed($unsigned(((reg47 ^ reg36) ?
                  (|(8'haa)) : reg47))) <= (|$unsigned(reg34)));
              reg49 = reg32[(1'h1):(1'h1)];
              reg50 = reg32[(1'h0):(1'h0)];
              reg51 <= (^reg36[(5'h12):(4'hb)]);
              reg52 = ((!$signed((wire24 ?
                      {reg48, (7'h44)} : reg41[(5'h15):(5'h15)]))) ?
                  (+(|(&(8'ha4)))) : (~^(reg36[(3'h4):(2'h2)] ?
                      (reg47[(2'h3):(2'h2)] ? reg35 : reg43) : reg36)));
            end
          else
            begin
              reg49 = forvar32;
              reg51 <= $unsigned($unsigned($signed(reg31)));
            end
        end
      reg53 <= {reg51[(3'h7):(1'h0)]};
      reg54 <= reg43;
    end
  module55 #() modinst242 (.wire57(reg30), .wire59(reg29), .y(wire241), .wire60(reg41), .wire58(reg48), .clk(clk), .wire56(reg46));
  assign wire243 = $signed(($signed(((+reg54) && (8'haf))) ?
                       (reg29 && reg48) : wire26[(1'h0):(1'h0)]));
  module244 #() modinst920 (.wire245(reg47), .wire246(wire27), .wire249(wire26), .clk(clk), .wire248(reg53), .wire247(reg46), .y(wire919));
  assign wire921 = $unsigned(($signed(reg37[(2'h3):(2'h3)]) & wire27));
  module385 #() modinst923 (.wire387(reg38), .wire388(wire243), .wire389(wire25), .y(wire922), .clk(clk), .wire386(reg48));
  always
    @(posedge clk) begin
      if ((8'hb8))
        begin
          reg924 <= ((reg44 ^ ($unsigned(reg46) >= (~|(wire921 == wire922)))) ^~ $unsigned(reg31));
        end
      else
        begin
          for (forvar924 = (1'h0); (forvar924 < (2'h2)); forvar924 = (forvar924 + (1'h1)))
            begin
              reg925 = ($unsigned($signed(reg42)) ?
                  {(8'ha6)} : (^$unsigned(($signed(reg53) ^ $signed(reg44)))));
              reg926 = (~^$signed(reg44));
              reg927 = $signed((reg42 <= (!(+reg30))));
              reg928 <= {(~|reg33[(4'h8):(3'h7)])};
              reg929 <= reg39[(3'h4):(3'h4)];
            end
        end
      reg930 <= (~reg33);
    end
  always
    @(posedge clk) begin
      reg931 <= (8'ha4);
    end
  always
    @(posedge clk) begin
      reg932 = (!($signed(reg51[(3'h4):(1'h1)]) <= reg931));
      if ((~^{$signed($unsigned((&reg53))),
          ($signed($signed(wire921)) == reg54[(4'h9):(3'h5)])}))
        begin
          if (wire24[(4'ha):(3'h4)])
            begin
              reg933 <= $unsigned($unsigned((~^$signed((reg39 < reg931)))));
              reg934 <= reg51[(2'h2):(1'h1)];
              reg935 = wire922;
              reg936 = (!(~^(~|$unsigned(reg39[(1'h1):(1'h0)]))));
            end
          else
            begin
              reg933 <= reg38[(1'h1):(1'h0)];
              reg935 = $signed((~|{wire28, {$signed(reg51), (-reg931)}}));
              reg936 = reg29;
              reg937 = wire921[(4'h8):(3'h4)];
            end
          if (((reg42 ?
                  $signed(reg929) : ((^reg933[(3'h5):(3'h4)]) ?
                      $unsigned(reg936[(4'ha):(4'h8)]) : ($signed((8'ha5)) | $unsigned(reg47)))) ?
              (reg935 ?
                  wire243[(4'hc):(3'h4)] : {(wire24 ?
                          {reg932} : reg935[(3'h5):(1'h1)])}) : (((((8'hba) ?
                              reg928 : (7'h46)) ?
                          (reg935 ? wire241 : reg934) : reg930[(3'h4):(1'h0)]) ?
                      ((8'hbc) + $signed(wire25)) : ((+(8'ha6)) & (reg54 ?
                          wire243 : reg41))) ?
                  ($signed($unsigned(reg933)) != wire243) : reg30)))
            begin
              reg938 <= {$signed(reg44),
                  $signed($unsigned($signed($signed(reg30))))};
              reg939 = $signed(($unsigned(({reg33, reg31} ?
                      (reg44 != wire25) : (^~reg53))) ?
                  (reg46[(5'h12):(5'h11)] ?
                      (7'h42) : wire28[(3'h4):(1'h0)]) : (&reg937[(4'ha):(4'h8)])));
            end
          else
            begin
              reg939 = $unsigned(reg935[(4'hb):(3'h6)]);
              reg940 = (8'h9d);
              reg941 = (8'ha5);
            end
          reg942 = reg934[(2'h3):(1'h0)];
          reg943 <= $signed((reg941 ^ $signed((~&wire26[(4'ha):(1'h1)]))));
        end
      else
        begin
          reg933 <= (reg47 ~^ (reg30 ?
              wire25[(4'ha):(3'h6)] : ($unsigned($unsigned(reg37)) | reg941)));
        end
    end
  always
    @(posedge clk) begin
      for (forvar944 = (1'h0); (forvar944 < (1'h0)); forvar944 = (forvar944 + (1'h1)))
        begin
          for (forvar945 = (1'h0); (forvar945 < (1'h0)); forvar945 = (forvar945 + (1'h1)))
            begin
              reg946 = ((8'hb8) ? $signed(reg37) : $unsigned(wire26));
              reg947 = {($unsigned(reg33) <= ({reg47, reg47} ?
                      (&reg37[(1'h1):(1'h0)]) : wire25))};
              reg948 <= reg933;
            end
          reg949 <= reg39[(2'h3):(2'h2)];
          reg950 = $signed(reg46[(3'h7):(3'h6)]);
          reg951 = (8'h9c);
          reg952 = {wire922[(2'h3):(2'h2)],
              {((+(reg48 && (8'hab))) - ((&reg48) | $unsigned(reg928))),
                  (|reg928[(3'h5):(2'h2)])}};
        end
      reg953 <= $signed(reg946);
      reg954 <= $unsigned({{reg42, reg949}});
    end
  assign wire955 = $signed($signed({(wire243 ?
                           $unsigned(reg37) : reg934[(3'h6):(3'h6)]),
                       (7'h4a)}));
  assign wire956 = {(8'hab),
                       (!({{(8'h9e), reg954}} << (wire922[(1'h1):(1'h1)] ?
                           (~reg30) : reg948[(4'h8):(1'h0)])))};
  always
    @(posedge clk) begin
      if ({wire921[(5'h12):(1'h1)]})
        begin
          reg957 = reg44[(2'h2):(1'h0)];
          reg958 <= ((reg934 ?
              wire241 : {(((7'h4a) <<< (7'h45)) ?
                      reg46[(4'he):(3'h6)] : (reg39 ?
                          reg933 : (8'hb3)))}) + $unsigned(reg931[(5'h17):(4'hc)]));
          for (forvar959 = (1'h0); (forvar959 < (1'h0)); forvar959 = (forvar959 + (1'h1)))
            begin
              reg960 = $signed($signed(reg29));
              reg961 <= (^$signed(reg46));
            end
        end
      else
        begin
          reg957 = $unsigned(reg933);
          for (forvar958 = (1'h0); (forvar958 < (3'h4)); forvar958 = (forvar958 + (1'h1)))
            begin
              reg959 = $signed((({$signed(reg958)} ?
                      (reg46 ^~ (reg954 ? reg51 : reg938)) : ((~^reg47) ?
                          (reg928 ? reg960 : (8'hb9)) : (~|reg51))) ?
                  (wire955 ^ wire28[(5'h10):(3'h7)]) : $unsigned((~|(-reg924)))));
              reg960 = ((~&($signed({(8'hb0), reg53}) ?
                      (reg37[(1'h1):(1'h1)] ?
                          (reg48 ~^ reg938) : (+reg42)) : (~&{(7'h44)}))) ?
                  reg948[(4'hb):(3'h7)] : ((($unsigned((8'haf)) <<< (~wire25)) ?
                      $signed((reg931 ?
                          (8'ha5) : wire28)) : (8'hb7)) <= reg29));
              reg962 = (({reg54[(1'h1):(1'h1)],
                      reg47} >= reg928[(4'hd):(4'hc)]) ?
                  (^(7'h47)) : $signed($signed($signed((reg948 ?
                      reg958 : reg948)))));
            end
          reg963 = (($signed(reg933[(3'h4):(2'h3)]) != $unsigned($signed((reg51 ?
              reg53 : wire922)))) ^~ (((reg948[(4'ha):(3'h4)] & $signed(reg42)) >>> wire24[(1'h0):(1'h0)]) ?
              (((reg929 ^~ (8'haf)) ? $signed(wire919) : (~&wire28)) ?
                  $unsigned($signed(reg33)) : $unsigned($signed(forvar959))) : reg961));
        end
    end
  always
    @(posedge clk) begin
      reg964 = $signed((({$unsigned(wire24)} ~^ {wire956[(3'h4):(2'h2)]}) ?
          reg44[(4'h8):(3'h6)] : (reg928 >> ($unsigned(wire919) * (wire241 & reg51)))));
      reg965 = {wire25,
          $signed(($unsigned((8'hbb)) ?
              reg961[(2'h3):(2'h3)] : $signed({reg943, reg933})))};
      for (forvar966 = (1'h0); (forvar966 < (1'h0)); forvar966 = (forvar966 + (1'h1)))
        begin
          for (forvar967 = (1'h0); (forvar967 < (1'h1)); forvar967 = (forvar967 + (1'h1)))
            begin
              reg968 <= ($signed(reg44[(2'h3):(1'h0)]) ?
                  reg47 : $unsigned(((reg933 ?
                      {reg46,
                          forvar967} : (^~reg931)) <<< reg924[(2'h3):(2'h2)])));
              reg969 <= $unsigned(((reg53[(4'ha):(3'h4)] | $signed((~&reg47))) ?
                  ($signed({wire956}) ?
                      ($unsigned(reg42) ?
                          (~&reg934) : (reg53 ? wire26 : wire922)) : (!(wire24 ?
                          (8'h9f) : wire956))) : $unsigned($unsigned(reg53[(4'hb):(4'h9)]))));
            end
          for (forvar970 = (1'h0); (forvar970 < (2'h2)); forvar970 = (forvar970 + (1'h1)))
            begin
              reg971 <= ((~$signed(reg51[(3'h7):(2'h2)])) ?
                  (((~(~^reg924)) ~^ $signed(reg51[(3'h4):(3'h4)])) >> $signed((~|$signed(reg928)))) : reg948);
              reg972 = reg928;
              reg973 = (((+($unsigned(reg971) + (reg51 ^~ reg934))) * reg38) << reg30[(4'he):(2'h3)]);
              reg974 <= ($signed($unsigned(({reg39} > $unsigned(reg972)))) ~^ ($unsigned((~^forvar966)) ?
                  reg44[(4'hd):(3'h7)] : ($unsigned(forvar967[(1'h1):(1'h0)]) ?
                      (^wire26[(2'h3):(1'h0)]) : $unsigned({forvar966,
                          reg51}))));
            end
          for (forvar975 = (1'h0); (forvar975 < (1'h1)); forvar975 = (forvar975 + (1'h1)))
            begin
              reg976 <= forvar966[(5'h11):(4'hc)];
              reg977 = reg931[(4'hd):(4'h8)];
            end
          reg978 = {$signed(reg48)};
        end
    end
  always
    @(posedge clk) begin
      if (reg971[(3'h5):(1'h0)])
        begin
          reg979 = reg933;
        end
      else
        begin
          reg979 = reg969[(4'hc):(2'h3)];
          if (reg47)
            begin
              reg980 = (^(($unsigned(reg31[(3'h5):(2'h2)]) ?
                      ($unsigned(reg42) < reg949[(2'h2):(2'h2)]) : $unsigned((reg33 ?
                          reg938 : reg974))) ?
                  $unsigned(($unsigned(reg33) + reg30)) : reg948));
              reg981 = {$unsigned((reg933[(1'h1):(1'h0)] >> reg47[(2'h3):(1'h1)]))};
            end
          else
            begin
              reg980 = (-$signed($unsigned(wire26)));
            end
          for (forvar982 = (1'h0); (forvar982 < (1'h0)); forvar982 = (forvar982 + (1'h1)))
            begin
              reg983 = reg981;
              reg984 = reg38;
              reg985 = (^~(~&wire26));
              reg986 <= reg31;
            end
        end
      if (($unsigned((($signed(reg47) ?
                  (reg953 | reg974) : $unsigned(wire955)) ?
              (wire25[(3'h4):(2'h2)] ?
                  $unsigned(wire919) : (reg930 <<< (8'hb0))) : $unsigned(wire25[(5'h10):(4'hc)]))) ?
          reg37 : reg931))
        begin
          for (forvar987 = (1'h0); (forvar987 < (2'h3)); forvar987 = (forvar987 + (1'h1)))
            begin
              reg988 = ((wire955 ?
                      (($signed(reg938) ?
                              wire956[(1'h0):(1'h0)] : (reg33 - reg961)) ?
                          reg53 : (wire921 ?
                              reg938[(1'h1):(1'h0)] : (reg943 ^ reg29))) : wire28) ?
                  ($signed(reg47[(3'h4):(1'h1)]) ?
                      (^$unsigned(reg46[(3'h6):(1'h0)])) : (8'hb0)) : $unsigned({(((8'ha6) ?
                              reg41 : reg984) ?
                          (&reg980) : wire26),
                      reg961[(2'h2):(1'h0)]}));
              reg989 = reg953[(4'h9):(4'h8)];
            end
          if (reg38)
            begin
              reg990 <= ($unsigned(((+reg929[(3'h6):(3'h4)]) | reg44[(2'h2):(2'h2)])) ^ $unsigned($signed($signed((reg44 >>> wire26)))));
              reg991 = reg47;
              reg992 <= $signed(($unsigned(reg991[(1'h1):(1'h0)]) ?
                  $signed($unsigned($signed(forvar987))) : $signed(wire28[(3'h4):(2'h3)])));
              reg993 <= wire243[(4'hd):(2'h3)];
              reg994 = $signed($signed(reg53[(4'h8):(2'h2)]));
            end
          else
            begin
              reg991 = ($unsigned({({reg984, wire26} ^~ (~&reg979))}) ?
                  wire241[(2'h3):(1'h0)] : (reg994[(2'h2):(1'h1)] ?
                      {reg54[(3'h6):(1'h0)]} : {(8'hab),
                          reg929[(3'h7):(3'h6)]}));
              reg994 = ($unsigned(wire243[(5'h12):(4'he)]) >= reg991[(2'h3):(1'h0)]);
              reg995 <= (~^(7'h47));
            end
          if ($unsigned((reg930[(4'hb):(3'h4)] || (8'ha7))))
            begin
              reg996 <= ((8'hb9) < $signed((|($unsigned(reg29) ?
                  $signed(wire27) : (reg953 ? reg928 : reg33)))));
              reg997 = (~^$unsigned({(8'hbb)}));
              reg998 = wire24[(3'h4):(1'h0)];
              reg999 <= {{reg53[(3'h5):(3'h5)], wire25}};
            end
          else
            begin
              reg996 <= ((reg48 ?
                      $unsigned({(-forvar987),
                          (reg54 ? forvar982 : wire919)}) : $unsigned(reg53)) ?
                  ($signed(reg948) ?
                      (($unsigned(reg979) ^ (reg31 ^ (8'hb3))) ?
                          reg999 : $signed(forvar982)) : ($unsigned(((8'haa) - (8'ha0))) ?
                          ($signed(reg943) ?
                              reg930 : (reg994 ?
                                  wire955 : wire24)) : $signed(reg41))) : $signed(wire955));
              reg999 <= reg928;
              reg1000 <= $unsigned(($signed((^~reg985)) ^ wire27[(3'h5):(3'h5)]));
              reg1001 <= reg38[(3'h7):(1'h1)];
            end
        end
      else
        begin
          for (forvar987 = (1'h0); (forvar987 < (1'h1)); forvar987 = (forvar987 + (1'h1)))
            begin
              reg990 <= $signed((((reg31[(2'h3):(1'h1)] << $unsigned(reg981)) != $signed(reg46)) ?
                  (($unsigned(wire922) ?
                      reg990 : $unsigned((7'h45))) <<< ((reg961 | reg38) ?
                      reg992 : (-reg931))) : (^((8'h9c) ?
                      $signed(reg1000) : $signed(reg929)))));
              reg992 <= wire956[(4'hc):(2'h2)];
              reg993 <= ($unsigned($unsigned($unsigned($unsigned((8'ha4))))) << (($unsigned((!(8'ha7))) ?
                      ($unsigned(forvar982) ~^ $signed(reg954)) : reg31[(1'h1):(1'h1)]) ?
                  $unsigned((7'h4a)) : $signed(reg988)));
              reg994 = $unsigned($unsigned(($signed($signed(reg961)) ?
                  reg995 : reg54)));
            end
          for (forvar995 = (1'h0); (forvar995 < (1'h0)); forvar995 = (forvar995 + (1'h1)))
            begin
              reg996 <= ((~|(^((8'hb2) >>> $signed(wire243)))) * ($unsigned((~|wire27[(3'h6):(2'h3)])) << reg997[(1'h0):(1'h0)]));
              reg999 <= $signed(reg39[(2'h3):(2'h3)]);
            end
          reg1002 = wire24;
          reg1003 = ((!(((~&reg1001) && reg989) ?
                  {$signed(reg39), ((8'hb1) ? reg992 : wire241)} : reg53)) ?
              (((7'h45) ? reg990 : forvar982) ?
                  (~&{(~|reg988),
                      (reg54 & wire955)}) : (+reg969[(5'h14):(3'h6)])) : (^$unsigned(($unsigned(forvar995) ?
                  wire956 : $signed(reg958)))));
          if ($signed((reg928 ?
              reg997[(1'h0):(1'h0)] : {$signed((reg933 ? reg42 : (8'ha0)))})))
            begin
              reg1004 <= $unsigned(($signed((reg995 ?
                      (reg985 && forvar982) : reg981)) ?
                  ($signed($unsigned(reg54)) >= $unsigned(reg1003)) : $signed($unsigned((&reg943)))));
              reg1005 = $signed($unsigned($signed($signed((wire922 ~^ reg933)))));
              reg1006 <= $unsigned(reg992);
              reg1007 = $signed($signed({$unsigned((reg924 ?
                      reg995 : reg934))}));
            end
          else
            begin
              reg1005 = wire956[(4'h9):(3'h7)];
              reg1006 <= $signed($unsigned({$signed((reg1006 & reg39)),
                  ($unsigned(reg979) + reg983[(3'h4):(3'h4)])}));
              reg1008 <= (|wire956[(4'hd):(3'h4)]);
            end
        end
      reg1009 = $unsigned($signed((!(~|(reg54 <<< (8'hac))))));
      if ((~|$signed(reg996[(3'h5):(1'h1)])))
        begin
          reg1010 = $unsigned($signed(((!(reg995 ^ wire922)) > ((forvar987 >= reg971) || (reg948 ?
              reg1003 : reg949)))));
          if ((&reg1001[(4'ha):(3'h4)]))
            begin
              reg1011 = (-({(forvar982 ?
                      (reg42 ? reg997 : reg984) : (&(8'ha9))),
                  (8'ha7)} ^~ (+reg995[(5'h15):(1'h0)])));
              reg1012 = reg988[(2'h2):(2'h2)];
            end
          else
            begin
              reg1011 = (8'ha3);
              reg1013 <= (^~wire28[(5'h12):(4'hf)]);
              reg1014 <= reg989[(3'h4):(2'h3)];
              reg1015 <= (reg47[(1'h1):(1'h1)] == ((reg997[(1'h1):(1'h0)] * reg928) || $unsigned($signed(reg47))));
              reg1016 = $signed($signed(reg980[(1'h0):(1'h0)]));
            end
          reg1017 = $unsigned({((8'hbc) ? (~|wire27) : (~(|forvar982)))});
        end
      else
        begin
          reg1013 <= reg989;
          reg1014 <= ($unsigned(reg938[(1'h0):(1'h0)]) ^ (~&reg1005));
          for (forvar1015 = (1'h0); (forvar1015 < (1'h0)); forvar1015 = (forvar1015 + (1'h1)))
            begin
              reg1016 = $signed(reg1015);
              reg1017 = $unsigned($unsigned($unsigned({reg51[(3'h6):(3'h4)]})));
              reg1018 = (((^$signed((reg1012 ? reg928 : reg928))) ?
                  {(reg992[(3'h4):(1'h0)] ? ((7'h47) >= reg949) : (~|reg998)),
                      reg38[(3'h7):(3'h4)]} : (reg1015 ?
                      reg971 : $signed((reg949 ?
                          forvar987 : wire919)))) ^~ reg994);
              reg1019 = (&(~&((wire922 ?
                      $unsigned(reg1011) : $unsigned(reg949)) ?
                  wire919 : $unsigned($signed(reg953)))));
            end
          reg1020 = (~($signed((+((8'h9d) ^~ (8'hab)))) | $signed($unsigned($signed(reg961)))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module244
#(parameter param917 = (!(~^{(((7'h42) ? (8'ha2) : (8'hb2)) ? {(8'h9f), (8'hbc)} : ((8'hbb) ? (8'hab) : (7'h46)))})), 
parameter param918 = param917)
(y, clk, wire245, wire246, wire247, wire248, wire249);
  output wire [(32'h89e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire245;
  input wire [(4'hf):(1'h0)] wire246;
  input wire signed [(5'h12):(1'h0)] wire247;
  input wire signed [(4'hb):(1'h0)] wire248;
  input wire signed [(4'hc):(1'h0)] wire249;
  wire signed [(3'h4):(1'h0)] wire915;
  wire [(5'h10):(1'h0)] wire676;
  wire signed [(5'h13):(1'h0)] wire675;
  wire [(4'he):(1'h0)] wire674;
  wire [(5'h14):(1'h0)] wire671;
  wire [(4'hb):(1'h0)] wire250;
  wire [(4'hd):(1'h0)] wire322;
  wire signed [(3'h6):(1'h0)] wire323;
  wire [(5'h17):(1'h0)] wire324;
  wire signed [(4'hb):(1'h0)] wire325;
  wire signed [(2'h2):(1'h0)] wire326;
  wire [(5'h12):(1'h0)] wire357;
  wire signed [(5'h15):(1'h0)] wire358;
  wire [(5'h15):(1'h0)] wire359;
  wire signed [(5'h15):(1'h0)] wire361;
  wire signed [(3'h4):(1'h0)] wire362;
  wire [(3'h5):(1'h0)] wire656;
  reg [(2'h2):(1'h0)] reg384 = (1'h0);
  reg [(4'hf):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg382 = (1'h0);
  reg [(4'he):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg377 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg374 = (1'h0);
  reg [(5'h10):(1'h0)] reg373 = (1'h0);
  reg [(5'h12):(1'h0)] reg372 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg368 = (1'h0);
  reg [(4'he):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg364 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg356 = (1'h0);
  reg [(4'h9):(1'h0)] reg355 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg352 = (1'h0);
  reg [(4'h8):(1'h0)] reg350 = (1'h0);
  reg [(5'h14):(1'h0)] reg349 = (1'h0);
  reg [(5'h18):(1'h0)] reg348 = (1'h0);
  reg [(4'h9):(1'h0)] reg344 = (1'h0);
  reg [(5'h18):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg335 = (1'h0);
  reg [(3'h4):(1'h0)] reg332 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg330 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg320 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg314 = (1'h0);
  reg [(4'hd):(1'h0)] reg311 = (1'h0);
  reg [(5'h14):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg299 = (1'h0);
  reg [(5'h15):(1'h0)] reg298 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg296 = (1'h0);
  reg [(5'h10):(1'h0)] reg295 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg286 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg285 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg283 = (1'h0);
  reg [(3'h5):(1'h0)] reg280 = (1'h0);
  reg [(2'h2):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg274 = (1'h0);
  reg [(5'h12):(1'h0)] reg273 = (1'h0);
  reg [(3'h5):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg269 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg263 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg260 = (1'h0);
  reg [(5'h10):(1'h0)] reg259 = (1'h0);
  reg [(5'h16):(1'h0)] reg258 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg257 = (1'h0);
  reg [(3'h7):(1'h0)] reg255 = (1'h0);
  reg [(3'h7):(1'h0)] reg254 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg251 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg659 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg663 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg665 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg668 = (1'h0);
  reg [(5'h10):(1'h0)] reg669 = (1'h0);
  reg [(5'h11):(1'h0)] reg673 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg672 = (1'h0);
  reg signed [(4'he):(1'h0)] reg670 = (1'h0);
  reg [(4'hf):(1'h0)] reg667 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg666 = (1'h0);
  reg [(4'hf):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg662 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg661 = (1'h0);
  reg [(4'ha):(1'h0)] reg660 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar658 = (1'h0);
  reg [(5'h12):(1'h0)] reg380 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg379 = (1'h0);
  reg [(4'he):(1'h0)] forvar378 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg376 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg375 = (1'h0);
  reg [(4'he):(1'h0)] reg370 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg371 = (1'h0);
  reg [(4'hf):(1'h0)] forvar370 = (1'h0);
  reg [(5'h10):(1'h0)] reg369 = (1'h0);
  reg [(4'h9):(1'h0)] reg366 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar365 = (1'h0);
  reg [(5'h18):(1'h0)] forvar363 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg360 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg354 = (1'h0);
  reg [(5'h18):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar351 = (1'h0);
  reg [(4'he):(1'h0)] forvar347 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar346 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg340 = (1'h0);
  reg [(5'h15):(1'h0)] reg339 = (1'h0);
  reg [(5'h12):(1'h0)] reg338 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg337 = (1'h0);
  reg [(5'h12):(1'h0)] reg336 = (1'h0);
  reg [(2'h2):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg333 = (1'h0);
  reg [(4'h8):(1'h0)] reg331 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg329 = (1'h0);
  reg [(4'h9):(1'h0)] reg328 = (1'h0);
  reg [(4'hf):(1'h0)] forvar327 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg321 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar318 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg317 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg316 = (1'h0);
  reg [(2'h2):(1'h0)] forvar315 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg313 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg309 = (1'h0);
  reg [(4'h8):(1'h0)] reg308 = (1'h0);
  reg [(5'h18):(1'h0)] forvar306 = (1'h0);
  reg [(4'hf):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg302 = (1'h0);
  reg [(5'h15):(1'h0)] reg301 = (1'h0);
  reg [(5'h12):(1'h0)] reg297 = (1'h0);
  reg [(4'ha):(1'h0)] reg294 = (1'h0);
  reg [(5'h12):(1'h0)] reg293 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg292 = (1'h0);
  reg signed [(4'he):(1'h0)] reg291 = (1'h0);
  reg [(5'h14):(1'h0)] reg290 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar289 = (1'h0);
  reg [(3'h7):(1'h0)] reg288 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg287 = (1'h0);
  reg [(4'hc):(1'h0)] forvar285 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg284 = (1'h0);
  reg [(4'hf):(1'h0)] forvar284 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg282 = (1'h0);
  reg [(4'hb):(1'h0)] reg281 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg277 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar266 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg265 = (1'h0);
  reg [(2'h3):(1'h0)] reg272 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg270 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg268 = (1'h0);
  reg [(4'hb):(1'h0)] reg267 = (1'h0);
  reg [(3'h5):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar265 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg261 = (1'h0);
  reg [(3'h5):(1'h0)] reg256 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar253 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar252 = (1'h0);
  assign y = {wire915,
                 wire676,
                 wire675,
                 wire674,
                 wire671,
                 wire250,
                 wire322,
                 wire323,
                 wire324,
                 wire325,
                 wire326,
                 wire357,
                 wire358,
                 wire359,
                 wire361,
                 wire362,
                 wire656,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg377,
                 reg374,
                 reg373,
                 reg372,
                 reg368,
                 reg367,
                 reg364,
                 reg356,
                 reg355,
                 reg352,
                 reg350,
                 reg349,
                 reg348,
                 reg344,
                 reg341,
                 reg335,
                 reg332,
                 reg330,
                 reg320,
                 reg319,
                 reg314,
                 reg311,
                 reg307,
                 reg305,
                 reg303,
                 reg300,
                 reg299,
                 reg298,
                 reg296,
                 reg295,
                 reg286,
                 reg285,
                 reg283,
                 reg280,
                 reg278,
                 reg275,
                 reg274,
                 reg273,
                 reg271,
                 reg269,
                 reg263,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg255,
                 reg254,
                 reg251,
                 reg659,
                 reg663,
                 reg665,
                 reg668,
                 reg669,
                 reg673,
                 reg672,
                 reg670,
                 reg667,
                 reg666,
                 reg664,
                 reg662,
                 reg661,
                 reg660,
                 forvar658,
                 reg380,
                 reg379,
                 forvar378,
                 reg376,
                 reg375,
                 reg370,
                 reg371,
                 forvar370,
                 reg369,
                 reg366,
                 forvar365,
                 forvar363,
                 reg360,
                 reg354,
                 reg353,
                 forvar351,
                 forvar347,
                 forvar346,
                 reg345,
                 reg343,
                 reg342,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg334,
                 reg333,
                 reg331,
                 reg329,
                 reg328,
                 forvar327,
                 reg321,
                 forvar318,
                 reg317,
                 reg316,
                 forvar315,
                 reg313,
                 reg312,
                 reg310,
                 reg309,
                 reg308,
                 forvar306,
                 reg304,
                 reg302,
                 reg301,
                 reg297,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 forvar289,
                 reg288,
                 reg287,
                 forvar285,
                 reg284,
                 forvar284,
                 reg282,
                 reg281,
                 reg279,
                 reg277,
                 reg276,
                 forvar266,
                 reg265,
                 reg272,
                 reg270,
                 reg268,
                 reg267,
                 reg266,
                 forvar265,
                 reg264,
                 reg262,
                 reg261,
                 reg256,
                 forvar253,
                 forvar252,
                 (1'h0)};
  assign wire250 = ((wire247[(4'h8):(1'h1)] && {($signed((8'ha3)) <= (~^wire249))}) + (wire245 ?
                       (wire248[(1'h1):(1'h0)] ?
                           ({(8'ha0), wire248} ?
                               $unsigned(wire249) : (wire247 ?
                                   wire246 : (8'hb7))) : (~wire249)) : wire249));
  always
    @(posedge clk) begin
      reg251 <= wire248;
      for (forvar252 = (1'h0); (forvar252 < (1'h0)); forvar252 = (forvar252 + (1'h1)))
        begin
          for (forvar253 = (1'h0); (forvar253 < (3'h4)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 <= forvar252;
              reg255 <= forvar253;
              reg256 = forvar252[(1'h1):(1'h0)];
              reg257 <= (~(+$signed((~|(wire248 + reg255)))));
              reg258 <= $unsigned($unsigned(reg254[(1'h1):(1'h1)]));
            end
          if ($unsigned((+$signed(($signed(reg251) * forvar252)))))
            begin
              reg259 <= ($signed($signed(forvar253)) ?
                  reg258 : wire250[(4'ha):(1'h1)]);
              reg260 <= reg251[(1'h0):(1'h0)];
              reg261 = $signed(wire250);
              reg262 = $unsigned($unsigned(((^~$signed(reg257)) <= $signed((^~wire245)))));
            end
          else
            begin
              reg259 <= reg260;
              reg260 <= ((wire249 ?
                  reg259[(4'h8):(3'h6)] : ($signed($signed(forvar253)) ?
                      (8'hbc) : $signed(wire246[(1'h1):(1'h1)]))) | wire250[(2'h3):(2'h3)]);
              reg263 <= $unsigned($signed(reg262));
            end
        end
      reg264 = $signed({(+($signed(wire249) ?
              $unsigned((7'h4a)) : $unsigned(reg257)))});
      if ($signed($signed((((-wire246) != (wire246 && reg254)) ?
          $unsigned((~|reg263)) : $signed(reg261[(4'hf):(1'h1)])))))
        begin
          for (forvar265 = (1'h0); (forvar265 < (2'h2)); forvar265 = (forvar265 + (1'h1)))
            begin
              reg266 = reg259;
              reg267 = reg255;
              reg268 = forvar252;
            end
          if ($signed(((reg257 ^~ $signed((reg263 ? reg257 : reg254))) ?
              {$signed(reg257),
                  (~&$unsigned(wire245))} : ($signed(wire246[(3'h7):(3'h6)]) ^~ {reg266[(2'h3):(2'h2)],
                  $unsigned(reg254)}))))
            begin
              reg269 <= $signed({$unsigned((forvar252 ? {reg258} : {reg257})),
                  (((^~wire247) <= ((8'ha3) ? reg260 : forvar252)) ?
                      (~|$unsigned(forvar265)) : reg266[(1'h1):(1'h1)])});
              reg270 = $unsigned((reg263[(4'hb):(4'h9)] | $signed(reg258[(4'hb):(3'h7)])));
              reg271 <= reg254;
              reg272 = (~|(8'ha6));
            end
          else
            begin
              reg269 <= (&{(^reg259)});
            end
        end
      else
        begin
          reg265 = ((+($unsigned($signed(reg268)) ?
              ($unsigned(reg257) ?
                  (reg271 * reg257) : (reg271 ?
                      forvar265 : (8'hbc))) : reg268[(4'ha):(1'h0)])) >>> $unsigned((($signed(wire248) ?
              reg272 : {wire246}) >= $unsigned(forvar253[(2'h2):(2'h2)]))));
          for (forvar266 = (1'h0); (forvar266 < (1'h1)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg269 <= (-forvar253);
              reg270 = ({(~|(+(~&reg263))),
                      (reg263[(4'hf):(4'hb)] != $signed({wire245, reg263}))} ?
                  reg257 : ((7'h45) ?
                      $unsigned(reg256) : $signed({$unsigned(wire245)})));
              reg271 <= (reg268 ?
                  (~|$signed(((forvar266 < reg266) == reg257))) : {reg264,
                      forvar252[(1'h0):(1'h0)]});
              reg272 = {{wire247, reg270}};
            end
          if (($signed((reg256[(2'h2):(1'h0)] ?
                  reg269[(3'h7):(3'h7)] : $signed($unsigned((7'h41))))) ?
              ((reg251[(1'h0):(1'h0)] ?
                  (forvar252 ?
                      (reg251 <<< reg266) : (~wire245)) : (~|$signed(reg260))) && $signed((forvar253 < reg265[(4'hd):(1'h1)]))) : (($signed((wire250 ^~ reg251)) ?
                      reg272[(2'h3):(1'h1)] : $signed((forvar266 < reg256))) ?
                  wire246 : $signed((+(wire247 >= (7'h4a)))))))
            begin
              reg273 <= $signed(reg256[(3'h4):(2'h3)]);
              reg274 <= (($unsigned(($signed(reg256) ?
                      $unsigned(reg262) : (reg273 ? reg263 : (8'hb6)))) ?
                  (($unsigned(reg267) >>> reg269[(4'hc):(3'h5)]) ?
                      ({reg268,
                          reg272} < $unsigned(reg255)) : reg258[(4'hb):(3'h4)]) : reg264[(4'hc):(3'h4)]) != $unsigned($unsigned($unsigned(wire249))));
              reg275 <= reg270[(1'h1):(1'h0)];
              reg276 = ($signed($signed(reg258)) >= (+$unsigned(reg261[(5'h14):(2'h2)])));
            end
          else
            begin
              reg276 = $unsigned((reg268[(4'ha):(4'h8)] ?
                  $unsigned(reg264[(2'h2):(2'h2)]) : (reg266[(1'h1):(1'h0)] != (!(reg264 ?
                      reg254 : (7'h40))))));
              reg277 = $unsigned(reg274);
              reg278 <= (reg273[(4'hd):(4'hd)] ?
                  wire249[(3'h4):(2'h3)] : ($unsigned($unsigned(((8'ha6) & (7'h43)))) ?
                      reg267 : reg273[(3'h7):(1'h0)]));
              reg279 = $signed(reg260);
              reg280 <= $unsigned(($unsigned({((8'hbe) ?
                      reg273 : wire246)}) * reg271[(2'h2):(1'h0)]));
            end
          reg281 = wire250[(1'h1):(1'h0)];
        end
      reg282 = ($unsigned((^reg269)) < reg254);
    end
  always
    @(posedge clk) begin
      if ((reg259[(5'h10):(3'h7)] * ($signed((~^wire246)) ?
          (~&(~$unsigned(wire246))) : $unsigned($signed((reg271 != reg259))))))
        begin
          reg283 <= (~reg257[(3'h7):(1'h0)]);
          for (forvar284 = (1'h0); (forvar284 < (1'h1)); forvar284 = (forvar284 + (1'h1)))
            begin
              reg285 <= (wire250 ?
                  ((reg251[(1'h1):(1'h1)] >> reg280) && ((^~wire249) ?
                      $unsigned($signed(reg259)) : ((reg254 ? reg260 : reg259) ?
                          $signed(reg271) : (8'ha0)))) : (8'hab));
              reg286 <= reg285;
            end
        end
      else
        begin
          reg284 = reg285;
          for (forvar285 = (1'h0); (forvar285 < (2'h2)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg287 = {(+(reg286 ?
                      $signed({reg271,
                          wire249}) : $signed($unsigned(forvar284))))};
              reg288 = ((!(({reg280} ? reg255 : {(7'h40)}) ?
                      (^~$unsigned(reg286)) : (wire250[(4'h9):(3'h6)] < (8'hb2)))) ?
                  (({reg286[(4'hb):(3'h4)], wire246} ?
                      (|reg273[(4'hc):(4'hc)]) : (~&wire249)) | $unsigned({$unsigned(reg275)})) : $unsigned($signed(forvar284[(1'h1):(1'h1)])));
            end
          for (forvar289 = (1'h0); (forvar289 < (2'h3)); forvar289 = (forvar289 + (1'h1)))
            begin
              reg290 = ((($signed(reg284) == $unsigned(wire250[(4'h9):(2'h3)])) ?
                  (^reg255) : forvar284[(3'h6):(2'h3)]) <= $unsigned((($signed((7'h40)) ?
                  $unsigned(reg263) : reg251) ^~ reg274[(4'h9):(3'h7)])));
              reg291 = (~&$unsigned((+(^wire246))));
              reg292 = reg274[(1'h0):(1'h0)];
              reg293 = reg269;
            end
          reg294 = ($unsigned(wire245[(2'h2):(2'h2)]) >= forvar284);
        end
    end
  always
    @(posedge clk) begin
      if (($unsigned({$unsigned(reg263)}) < reg269[(5'h13):(3'h7)]))
        begin
          reg295 <= $signed((~&{$signed($signed((8'hb8))),
              ((reg271 | wire247) ? (-reg275) : reg273)}));
          reg296 <= $unsigned(wire250[(3'h6):(2'h2)]);
          if ((reg286[(4'h8):(1'h0)] ?
              (8'hb7) : (reg296[(4'hb):(3'h7)] ^~ reg259[(1'h1):(1'h0)])))
            begin
              reg297 = reg275;
            end
          else
            begin
              reg298 <= $unsigned(reg269[(5'h13):(2'h2)]);
              reg299 <= {((reg298[(4'hc):(1'h1)] ?
                          reg280 : ($unsigned(wire246) - (reg274 << reg258))) ?
                      reg258 : (wire248 << ($signed(reg283) || (^reg296)))),
                  $unsigned({($unsigned(wire245) ?
                          $signed(reg273) : reg254[(2'h3):(1'h1)]),
                      reg280})};
              reg300 <= $unsigned(reg280);
              reg301 = reg280;
              reg302 = (((|((wire247 ^ wire246) ?
                  (reg255 - (7'h46)) : reg273)) >= $signed($signed(reg257))) - $unsigned((|{(8'had)})));
            end
          reg303 <= (!$signed(reg297[(3'h7):(3'h4)]));
          reg304 = reg258[(4'hf):(3'h4)];
        end
      else
        begin
          reg297 = $unsigned($signed((((~^(7'h4a)) ?
              $unsigned(wire249) : $signed(wire245)) - ({reg297, reg295} ?
              (wire246 ^~ reg301) : (^reg296)))));
          reg301 = (~|$unsigned((~{$signed(wire246)})));
          reg303 <= reg297[(4'hf):(2'h2)];
          reg305 <= (reg259[(4'ha):(3'h6)] ?
              $signed(reg271[(3'h4):(3'h4)]) : $unsigned({reg296,
                  reg259[(1'h1):(1'h0)]}));
        end
      for (forvar306 = (1'h0); (forvar306 < (1'h1)); forvar306 = (forvar306 + (1'h1)))
        begin
          if (reg257[(1'h1):(1'h1)])
            begin
              reg307 <= (!((reg274 && $signed($unsigned(reg305))) ?
                  ((&reg296) & wire249[(4'hb):(3'h5)]) : $signed(wire249)));
              reg308 = reg295[(2'h2):(1'h0)];
              reg309 = forvar306[(5'h12):(3'h5)];
              reg310 = $unsigned($signed(((&((8'hac) << (8'hab))) ?
                  (~^reg303[(3'h6):(3'h4)]) : (&{(7'h41), reg302}))));
            end
          else
            begin
              reg307 <= $signed((reg254 ?
                  {$signed((|reg254)),
                      reg260[(2'h3):(2'h2)]} : $signed(($signed(reg275) ?
                      reg263 : reg278[(2'h2):(1'h1)]))));
              reg311 <= reg297[(4'hf):(3'h4)];
              reg312 = (wire250[(4'h9):(3'h7)] ? {reg260} : reg263);
              reg313 = reg310[(1'h0):(1'h0)];
              reg314 <= ((8'ha0) <= $signed((reg280 >= (~|$signed(reg309)))));
            end
          for (forvar315 = (1'h0); (forvar315 < (1'h1)); forvar315 = (forvar315 + (1'h1)))
            begin
              reg316 = (($unsigned(((~^reg310) ?
                  (|reg301) : (~&reg283))) ^~ $unsigned($unsigned((reg308 + reg297)))) <<< (reg308[(3'h4):(1'h0)] ?
                  reg283[(4'h9):(1'h0)] : ((!(^~(8'haf))) ?
                      ($signed(wire246) ?
                          $unsigned((8'hbc)) : (reg278 ?
                              reg296 : reg269)) : $signed((wire246 << reg298)))));
            end
          reg317 = wire246[(3'h6):(3'h4)];
          for (forvar318 = (1'h0); (forvar318 < (1'h0)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg319 <= reg305;
            end
          reg320 <= (-reg310);
        end
      reg321 = reg319;
    end
  assign wire322 = reg257[(4'h9):(1'h0)];
  assign wire323 = (^~(+(!{$signed((7'h42)), (wire247 < reg298)})));
  assign wire324 = $unsigned($unsigned((-$unsigned($signed((8'hbd))))));
  assign wire325 = reg295[(4'hb):(2'h3)];
  assign wire326 = (~&(reg303 ^ $signed($signed(wire325))));
  always
    @(posedge clk) begin
      for (forvar327 = (1'h0); (forvar327 < (1'h0)); forvar327 = (forvar327 + (1'h1)))
        begin
          reg328 = (reg251[(3'h6):(2'h2)] ?
              $signed((wire324 - $signed(reg314[(1'h1):(1'h0)]))) : ((wire249 ?
                  $signed((reg285 ?
                      reg299 : reg314)) : (~|reg295)) - ($signed($signed(wire245)) + forvar327[(3'h6):(3'h5)])));
        end
      reg329 = reg328;
      if ({((($unsigned(wire246) << {reg285,
              reg298}) ^~ $unsigned({reg259})) < ((~(8'hb2)) > $unsigned((reg260 || reg295)))),
          {reg274}})
        begin
          reg330 <= reg311;
          if ($unsigned(($unsigned((reg298 - $unsigned((8'haa)))) ?
              wire324[(3'h4):(2'h2)] : {reg271})))
            begin
              reg331 = reg254[(3'h5):(3'h5)];
              reg332 <= reg303[(1'h0):(1'h0)];
              reg333 = reg332;
              reg334 = reg330[(3'h4):(2'h2)];
            end
          else
            begin
              reg332 <= ((|$unsigned($signed(reg295))) ?
                  reg271 : (wire323[(3'h5):(1'h1)] ? wire326 : wire250));
              reg335 <= (^~$unsigned((^(wire249[(4'hb):(1'h1)] ?
                  (^wire325) : reg330))));
            end
          reg336 = {((wire323 << reg263) <= $signed((~|(reg298 < reg263))))};
          if (($signed($unsigned($signed(reg283))) ?
              (($signed((reg257 ?
                  reg332 : reg280)) < ($unsigned((8'hb2)) ^~ reg295)) ^~ (($unsigned(reg258) != reg300[(4'hf):(4'hc)]) ?
                  ($signed(wire245) ^~ (reg296 ?
                      (8'ha4) : wire246)) : wire326[(2'h2):(1'h0)])) : ($signed($unsigned($unsigned(reg285))) + wire326)))
            begin
              reg337 = $unsigned((reg307 ?
                  {reg320} : {$signed($signed(reg300)), (~(~wire324))}));
              reg338 = (7'h43);
              reg339 = ({reg257, (&reg332)} ?
                  $unsigned(($signed((reg280 || reg337)) ?
                      ((8'hac) ?
                          (~|reg299) : $signed(reg320)) : reg275[(4'he):(4'h8)])) : {(reg298 == (8'h9d))});
              reg340 = $unsigned((reg251 ?
                  ((((8'ha3) ? reg278 : reg269) ?
                      {wire249} : {reg254}) == wire324[(5'h14):(1'h1)]) : ({reg273[(4'he):(3'h6)],
                          $signed(wire249)} ?
                      (~^$unsigned(wire247)) : (7'h46))));
            end
          else
            begin
              reg341 <= (&reg271[(2'h2):(1'h1)]);
            end
          reg342 = (({reg335} <= (reg269[(5'h13):(4'hf)] + $unsigned(reg330[(2'h3):(1'h0)]))) - (8'h9c));
        end
      else
        begin
          if (reg331[(3'h5):(3'h4)])
            begin
              reg330 <= $unsigned({(~^$signed($signed(reg255))),
                  (((reg286 ? wire250 : wire324) ?
                      (8'haa) : ((8'haa) | reg296)) ^ reg269)});
            end
          else
            begin
              reg331 = ((|((^~(reg263 ? reg295 : reg298)) ?
                  $signed((reg259 ?
                      reg299 : reg269)) : {(~^reg341)})) & {reg275,
                  $unsigned(reg340[(2'h2):(2'h2)])});
              reg332 <= reg295;
              reg333 = (^(^~reg274[(4'hf):(2'h2)]));
              reg335 <= ($unsigned((8'ha2)) ?
                  (((((8'hb1) << reg255) - (^reg319)) ?
                          reg258[(5'h13):(5'h12)] : $signed($unsigned(reg319))) ?
                      (reg260[(3'h4):(1'h1)] > (!reg271)) : {($signed(wire245) < reg259[(4'ha):(4'h8)])}) : reg263[(4'he):(4'hd)]);
              reg336 = $signed(reg337);
            end
          reg337 = (^~$unsigned($unsigned($signed((reg260 ~^ wire248)))));
          reg341 <= ($unsigned(($unsigned((wire248 ?
                  reg286 : reg285)) >> {$signed(forvar327), reg341})) ?
              $unsigned($signed($signed(reg328))) : (^{($signed(reg286) ?
                      (reg283 ? reg269 : (8'hbe)) : (reg298 ? reg296 : reg263)),
                  (|reg280)}));
          if ($unsigned((7'h46)))
            begin
              reg342 = $unsigned((($unsigned(reg331[(3'h5):(2'h3)]) <<< (!(|reg299))) ?
                  (~&(-(~&wire250))) : $unsigned($signed(wire247))));
              reg343 = (wire246[(4'hb):(2'h3)] ?
                  ($signed(($signed(reg260) ~^ (reg330 | reg258))) ?
                      {(reg338 ?
                              $signed(reg337) : ((8'ha5) > reg271))} : $signed(($unsigned(reg332) ?
                          ((7'h46) >= reg319) : $signed(reg339)))) : reg280);
              reg344 <= $signed($signed((reg255[(2'h2):(1'h0)] & ((reg255 ~^ wire326) ?
                  (7'h45) : reg331[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg344 <= ($unsigned((((reg342 & (8'hbf)) ?
                      reg311[(2'h3):(2'h3)] : (reg255 | reg273)) ?
                  (~^(&wire247)) : ($unsigned(reg298) <= wire326))) >>> (((reg341 * (|reg271)) > (wire247 * {reg259})) <= ($signed(reg340[(4'h8):(4'h8)]) == (reg255[(3'h4):(2'h2)] ~^ $unsigned(forvar327)))));
              reg345 = $signed((~&(~^$unsigned($signed(wire247)))));
            end
        end
      for (forvar346 = (1'h0); (forvar346 < (1'h0)); forvar346 = (forvar346 + (1'h1)))
        begin
          for (forvar347 = (1'h0); (forvar347 < (3'h4)); forvar347 = (forvar347 + (1'h1)))
            begin
              reg348 <= (reg275[(3'h5):(3'h5)] != reg336);
              reg349 <= (!$signed((($signed(reg255) - (wire325 || reg348)) >= $unsigned((~reg285)))));
              reg350 <= $unsigned(({reg335} | reg338));
            end
          for (forvar351 = (1'h0); (forvar351 < (2'h2)); forvar351 = (forvar351 + (1'h1)))
            begin
              reg352 <= $signed((+$signed((+$unsigned(reg254)))));
              reg353 = reg339[(5'h12):(2'h3)];
              reg354 = $unsigned($unsigned(reg319[(1'h0):(1'h0)]));
            end
          reg355 <= reg260[(1'h0):(1'h0)];
        end
      reg356 <= reg329;
    end
  assign wire357 = (8'ha5);
  assign wire358 = $signed(wire246[(4'h9):(2'h2)]);
  assign wire359 = reg335;
  always
    @(posedge clk) begin
      reg360 = reg251[(1'h1):(1'h0)];
    end
  assign wire361 = {$unsigned({($unsigned(reg269) ^ (wire325 ?
                               reg251 : reg283)),
                           ((|reg299) || $unsigned(wire324))})};
  assign wire362 = $unsigned(reg311);
  always
    @(posedge clk) begin
      for (forvar363 = (1'h0); (forvar363 < (3'h4)); forvar363 = (forvar363 + (1'h1)))
        begin
          reg364 <= (&reg285[(1'h0):(1'h0)]);
          for (forvar365 = (1'h0); (forvar365 < (3'h4)); forvar365 = (forvar365 + (1'h1)))
            begin
              reg366 = (-reg311[(1'h1):(1'h1)]);
              reg367 <= wire322;
              reg368 <= wire248;
            end
        end
      reg369 = (({reg254[(3'h4):(1'h0)]} < reg255) << ($signed(($unsigned(reg269) <= $signed(reg269))) <= {$signed(wire357)}));
      if ((&$signed(wire249[(4'h8):(4'h8)])))
        begin
          for (forvar370 = (1'h0); (forvar370 < (2'h2)); forvar370 = (forvar370 + (1'h1)))
            begin
              reg371 = reg364;
              reg372 <= (~reg366);
            end
          reg373 <= {reg274,
              ((reg307 ? reg320 : $unsigned($unsigned(reg286))) ?
                  reg305[(4'ha):(1'h1)] : $signed($signed((reg314 ?
                      (7'h41) : reg280))))};
        end
      else
        begin
          if ((+((~{reg303}) ?
              $signed((+$signed(reg371))) : wire361[(5'h13):(4'hf)])))
            begin
              reg370 = (~({(reg348[(3'h7):(2'h2)] != (wire245 ?
                      (7'h48) : wire245))} >= reg278[(2'h2):(2'h2)]));
              reg371 = ($signed(wire359) || reg274[(4'h8):(2'h2)]);
              reg372 <= {((8'hba) == forvar363[(5'h15):(1'h1)]),
                  (|((~|$signed(reg364)) && $unsigned((wire362 ?
                      reg332 : reg373))))};
              reg373 <= ((~&(((reg314 ? reg271 : reg305) >= {reg341,
                      wire247}) | $signed((reg271 ? reg348 : reg355)))) ?
                  ((8'hbd) ?
                      (+($unsigned(reg271) * $signed(reg271))) : ({reg259} >> (((7'h47) != reg286) ?
                          $unsigned((8'hb9)) : $unsigned(reg275)))) : $signed(wire323[(3'h5):(1'h1)]));
              reg374 <= reg283[(2'h2):(1'h0)];
            end
          else
            begin
              reg370 = (8'ha8);
              reg371 = (reg369 <= $unsigned(reg319));
              reg375 = (^~{$unsigned(reg370[(4'hd):(3'h5)]),
                  ($unsigned($signed(reg320)) - {(7'h46), reg271})});
              reg376 = {$signed({(wire248[(1'h0):(1'h0)] ?
                          ((8'ha6) >> reg370) : (reg259 ? reg368 : reg341))}),
                  {{$unsigned((8'hbd))}}};
            end
          reg377 <= (reg350 >= ($unsigned($signed($unsigned(reg286))) ?
              {((~wire250) ? $signed(reg254) : (+(8'hb3)))} : $signed(reg258)));
          for (forvar378 = (1'h0); (forvar378 < (1'h1)); forvar378 = (forvar378 + (1'h1)))
            begin
              reg379 = reg296[(4'he):(4'hd)];
              reg380 = reg352;
              reg381 <= reg254;
              reg382 <= (reg274[(5'h13):(2'h3)] >> reg352[(3'h7):(3'h4)]);
              reg383 <= $signed({reg285,
                  (forvar363 ? $unsigned(reg283) : reg283)});
            end
        end
      reg384 <= (reg352 ?
          reg299 : (~&($unsigned(reg295) ?
              ($unsigned(reg332) ~^ (reg300 >>> reg364)) : (reg355 ?
                  $unsigned(reg372) : $unsigned(reg257)))));
    end
  module385 #() modinst657 (.wire387(reg372), .wire389(wire359), .y(wire656), .clk(clk), .wire386(reg314), .wire388(reg298));
  always
    @(posedge clk) begin
      for (forvar658 = (1'h0); (forvar658 < (1'h1)); forvar658 = (forvar658 + (1'h1)))
        begin
          reg659 <= reg382;
          reg660 = (8'had);
          if ((((reg271[(1'h1):(1'h0)] ? reg341 : ((!reg273) << reg271)) ?
              (^~{(!(8'haa))}) : $signed(((reg280 ?
                  reg341 : reg275) <= $unsigned(reg382)))) <<< $unsigned((((wire322 ?
              (7'h41) : reg341) + (reg377 ? (8'ha9) : reg273)) != reg356))))
            begin
              reg661 = reg355[(2'h2):(1'h1)];
              reg662 = (+((((reg274 ? reg295 : reg348) ?
                          {reg278} : $unsigned((8'hb0))) ?
                      (~^(reg381 >= reg335)) : $unsigned((wire359 ?
                          reg344 : reg255))) ?
                  ((~|reg259) ?
                      (reg305[(4'hf):(4'h9)] <<< (^reg260)) : reg320[(4'hd):(3'h5)]) : {$signed((wire323 ?
                          reg271 : wire357)),
                      (reg364 ?
                          $signed(reg298) : (wire246 ? reg273 : wire248))}));
              reg663 <= $signed($signed($unsigned(reg298[(3'h5):(2'h2)])));
              reg664 = (~|(&(+($signed((8'ha4)) ?
                  (reg273 ? reg659 : reg350) : wire324))));
            end
          else
            begin
              reg661 = $signed({reg383[(3'h6):(1'h0)],
                  (~&((&reg368) - $unsigned(reg335)))});
              reg663 <= (~|$unsigned(((wire248 ? wire656 : reg286) ?
                  $signed($signed((8'h9d))) : reg299[(5'h17):(1'h0)])));
              reg665 <= ($signed(($signed((reg381 ? reg285 : reg286)) ?
                  $signed($unsigned(reg377)) : {reg377})) ^~ (($unsigned(reg295[(4'hd):(4'ha)]) <= $signed((wire247 ?
                  (8'hb6) : (8'hb7)))) >>> (~reg300[(3'h6):(2'h3)])));
              reg666 = reg257;
            end
          reg667 = $signed(reg269);
          if (reg330)
            begin
              reg668 <= ((!$signed($unsigned($unsigned(reg384)))) > $signed(wire247[(4'h8):(3'h4)]));
              reg669 <= $unsigned($signed(({((8'hb3) > wire325),
                      $signed(reg283)} ?
                  $unsigned($signed(reg352)) : (!$signed((8'ha3))))));
              reg670 = (reg667 >= (8'h9c));
            end
          else
            begin
              reg670 = (reg296 ?
                  (!(($signed(reg367) ? (&reg285) : (&(8'h9e))) ?
                      ($signed(reg263) ?
                          reg251 : $unsigned(wire656)) : wire656)) : ($signed(($unsigned(reg372) ?
                      (reg251 ? reg298 : reg344) : (^~reg278))) - (&(8'hb7))));
            end
        end
    end
  assign wire671 = ((^reg273) < {((~|((7'h48) && reg349)) ?
                           (~^{reg263, (8'hba)}) : reg280[(2'h3):(2'h3)]),
                       reg356[(1'h1):(1'h1)]});
  always
    @(posedge clk) begin
      reg672 = $unsigned($unsigned(({reg273} ?
          wire357[(3'h5):(2'h2)] : reg280[(2'h2):(1'h1)])));
      reg673 = {wire361,
          ({{reg274, $unsigned(wire248)}} ?
              (($signed(reg300) >>> (reg364 ? (8'haa) : (7'h40))) ?
                  reg305[(2'h3):(2'h2)] : wire361) : $signed(reg344))};
    end
  assign wire674 = $signed((-((-$unsigned(reg356)) ?
                       (!$unsigned(reg383)) : reg303)));
  assign wire675 = (~(~^((reg381[(4'hb):(1'h0)] || (~|reg663)) ?
                       (^~(reg659 ? (8'h9c) : reg335)) : (-{reg341}))));
  assign wire676 = $unsigned(reg381[(1'h1):(1'h1)]);
  module677 #() modinst916 (wire915, clk, reg372, reg348, reg320, reg341, reg286);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module55
#(parameter param239 = (~&(((((8'haf) >= (8'h9e)) ^ (~&(8'haf))) ? (7'h48) : (8'had)) ? ({((8'hae) ? (8'hab) : (7'h42))} && (((7'h49) ? (7'h43) : (8'hbb)) ? (8'hb4) : ((8'h9f) ? (8'h9f) : (7'h41)))) : {((8'hbb) + (^~(8'ha5))), (((8'h9e) ? (8'hae) : (7'h45)) ? {(8'ha7), (8'ha6)} : ((7'h41) <<< (8'hb7)))})), 
parameter param240 = param239)
(y, clk, wire60, wire59, wire58, wire57, wire56);
  output wire [(32'h31c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire60;
  input wire signed [(3'h5):(1'h0)] wire59;
  input wire [(2'h3):(1'h0)] wire58;
  input wire signed [(5'h11):(1'h0)] wire57;
  input wire signed [(4'hc):(1'h0)] wire56;
  wire [(4'hb):(1'h0)] wire216;
  wire signed [(5'h13):(1'h0)] wire215;
  wire signed [(5'h14):(1'h0)] wire213;
  wire [(5'h11):(1'h0)] wire72;
  reg signed [(4'h8):(1'h0)] reg237 = (1'h0);
  reg [(5'h14):(1'h0)] reg234 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg233 = (1'h0);
  reg [(5'h15):(1'h0)] reg231 = (1'h0);
  reg [(3'h7):(1'h0)] reg230 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg229 = (1'h0);
  reg [(5'h16):(1'h0)] reg227 = (1'h0);
  reg [(3'h5):(1'h0)] reg226 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg224 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg219 = (1'h0);
  reg [(2'h2):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg88 = (1'h0);
  reg [(4'h8):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg81 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg80 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg68 = (1'h0);
  reg [(3'h4):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg62 = (1'h0);
  reg [(3'h4):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg238 = (1'h0);
  reg [(5'h14):(1'h0)] reg236 = (1'h0);
  reg signed [(4'he):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg232 = (1'h0);
  reg [(5'h10):(1'h0)] reg228 = (1'h0);
  reg [(5'h12):(1'h0)] forvar222 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg220 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg218 = (1'h0);
  reg [(3'h7):(1'h0)] forvar217 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg92 = (1'h0);
  reg [(2'h3):(1'h0)] reg91 = (1'h0);
  reg [(5'h18):(1'h0)] forvar90 = (1'h0);
  reg [(2'h3):(1'h0)] reg89 = (1'h0);
  reg [(5'h14):(1'h0)] reg87 = (1'h0);
  reg [(5'h10):(1'h0)] forvar85 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg84 = (1'h0);
  reg signed [(4'he):(1'h0)] reg83 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg82 = (1'h0);
  reg [(5'h15):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg77 = (1'h0);
  reg [(4'h9):(1'h0)] forvar75 = (1'h0);
  reg [(3'h5):(1'h0)] reg74 = (1'h0);
  reg [(4'h8):(1'h0)] reg73 = (1'h0);
  reg [(5'h18):(1'h0)] reg71 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg70 = (1'h0);
  reg [(4'he):(1'h0)] reg69 = (1'h0);
  reg [(4'ha):(1'h0)] forvar64 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg65 = (1'h0);
  reg [(5'h15):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg63 = (1'h0);
  assign y = {wire216,
                 wire215,
                 wire213,
                 wire72,
                 reg237,
                 reg234,
                 reg233,
                 reg231,
                 reg230,
                 reg229,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg221,
                 reg219,
                 reg85,
                 reg88,
                 reg86,
                 reg81,
                 reg80,
                 reg76,
                 reg68,
                 reg67,
                 reg66,
                 reg62,
                 reg61,
                 reg238,
                 reg236,
                 reg235,
                 reg232,
                 reg228,
                 forvar222,
                 reg220,
                 reg218,
                 forvar217,
                 reg92,
                 reg91,
                 forvar90,
                 reg89,
                 reg87,
                 forvar85,
                 reg84,
                 reg83,
                 reg82,
                 reg79,
                 reg78,
                 reg77,
                 forvar75,
                 reg74,
                 reg73,
                 reg71,
                 reg70,
                 reg69,
                 forvar64,
                 reg65,
                 reg64,
                 reg63,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg61 <= {$unsigned($unsigned($signed($signed(wire59)))),
          (-$unsigned((&$signed(wire57))))};
      if ((~&wire58[(2'h2):(1'h0)]))
        begin
          if (wire60[(2'h3):(1'h0)])
            begin
              reg62 <= (~^(wire57[(4'hc):(1'h0)] ?
                  $signed(($signed(wire56) ?
                      reg61 : (^~reg61))) : wire60[(3'h5):(3'h5)]));
              reg63 = {wire57,
                  ($signed((~^{wire58, wire60})) ?
                      ({$signed(wire57), wire56} ?
                          wire57 : $unsigned(wire58)) : $signed(wire57[(4'hb):(2'h2)]))};
              reg64 = $unsigned($unsigned($unsigned((^{reg62, (8'had)}))));
              reg65 = $unsigned((~^(8'hb4)));
              reg66 <= reg63[(3'h5):(2'h3)];
            end
          else
            begin
              reg63 = $unsigned($signed(((~(8'hb4)) ?
                  reg63[(3'h6):(1'h1)] : reg61)));
              reg66 <= wire60;
            end
        end
      else
        begin
          reg63 = $unsigned($unsigned((((~wire59) ?
              wire58 : (wire58 ?
                  wire60 : reg63)) << ($signed(wire59) < (reg63 << wire59)))));
          for (forvar64 = (1'h0); (forvar64 < (2'h3)); forvar64 = (forvar64 + (1'h1)))
            begin
              reg66 <= wire56[(4'hb):(4'hb)];
              reg67 <= $unsigned(reg64[(4'hb):(2'h3)]);
              reg68 <= $signed($signed($unsigned($signed($unsigned(reg62)))));
              reg69 = ((wire57[(2'h2):(2'h2)] ?
                  (~&$signed($unsigned(reg67))) : {({wire56, reg64} ?
                          wire57 : (~^reg64))}) & (!((reg64 && (-(8'haa))) ^ (-reg63[(4'hc):(4'h9)]))));
              reg70 = {reg61, $unsigned(wire57[(3'h7):(2'h3)])};
            end
        end
      reg71 = (reg62[(5'h10):(3'h4)] ?
          reg63 : $unsigned($signed((~&$unsigned(wire60)))));
    end
  assign wire72 = (~&reg68);
  always
    @(posedge clk) begin
      reg73 = $signed(wire60[(3'h6):(3'h6)]);
      reg74 = wire56;
      for (forvar75 = (1'h0); (forvar75 < (3'h4)); forvar75 = (forvar75 + (1'h1)))
        begin
          reg76 <= $signed(wire72);
          if ((((+reg66) <= ($unsigned((reg62 >= reg66)) + $signed((+wire59)))) ?
              wire57[(4'hf):(4'he)] : $signed(reg67[(1'h0):(1'h0)])))
            begin
              reg77 = ($unsigned((8'ha2)) ?
                  wire57[(5'h10):(4'h9)] : ((reg66 ?
                      $signed(((8'h9e) ?
                          (8'hb0) : wire59)) : ($unsigned(wire56) ?
                          (wire72 == reg76) : (~^wire58))) ~^ $unsigned($unsigned((~^reg74)))));
              reg78 = reg77[(5'h17):(4'hf)];
              reg79 = (($unsigned(((wire59 ? (8'ha2) : reg77) || reg67)) ?
                      $signed((~reg76[(1'h1):(1'h0)])) : $signed(wire57[(3'h4):(2'h2)])) ?
                  reg77 : (+(reg61[(1'h1):(1'h0)] * ($unsigned(reg78) == (reg62 ?
                      reg73 : reg67)))));
              reg80 <= ($unsigned({forvar75[(4'h8):(3'h4)]}) ?
                  {$signed((!(reg74 >= forvar75))),
                      ($signed(reg77[(5'h15):(3'h4)]) < ((~|(7'h49)) >= (reg67 ?
                          (8'hb1) : wire60)))} : reg74[(1'h1):(1'h0)]);
              reg81 <= (+{reg80, $signed(reg76[(1'h1):(1'h1)])});
            end
          else
            begin
              reg80 <= reg62;
            end
          reg82 = (!(|wire58[(2'h3):(2'h2)]));
          reg83 = (~$unsigned(wire56[(2'h2):(1'h0)]));
        end
    end
  always
    @(posedge clk) begin
      reg84 = $signed((reg80 <<< ((wire60 <<< (wire60 << wire57)) ?
          reg81[(3'h7):(3'h6)] : ($signed(wire57) & $signed(reg81)))));
      if ($signed($signed(((reg62 << (wire56 > wire72)) ?
          wire56[(4'h8):(1'h1)] : wire57))))
        begin
          for (forvar85 = (1'h0); (forvar85 < (1'h0)); forvar85 = (forvar85 + (1'h1)))
            begin
              reg86 <= (8'hb7);
              reg87 = {(8'hb1)};
              reg88 <= wire58;
              reg89 = $unsigned({(^reg68[(4'h9):(2'h2)]), (reg66 == reg76)});
            end
        end
      else
        begin
          reg85 <= $signed((reg76 ?
              $unsigned(wire58) : $signed($signed((|(8'ha0))))));
          reg87 = reg80[(1'h0):(1'h0)];
        end
      for (forvar90 = (1'h0); (forvar90 < (3'h4)); forvar90 = (forvar90 + (1'h1)))
        begin
          if ((&(&wire72)))
            begin
              reg91 = (8'h9e);
            end
          else
            begin
              reg91 = $signed(($signed(((~^reg67) + ((7'h40) != reg89))) >>> ((&reg91) ?
                  reg66 : ($signed(reg84) ~^ reg80))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg92 = wire57;
    end
  module93 #() modinst214 (.wire94(reg88), .wire97(wire57), .clk(clk), .wire95(wire56), .y(wire213), .wire96(reg68));
  assign wire215 = wire213;
  assign wire216 = wire56;
  always
    @(posedge clk) begin
      for (forvar217 = (1'h0); (forvar217 < (1'h1)); forvar217 = (forvar217 + (1'h1)))
        begin
          if ((|((&(7'h46)) ?
              reg76 : (~&($signed(wire59) | reg66[(4'h8):(3'h6)])))))
            begin
              reg218 = (-wire215[(2'h2):(1'h1)]);
              reg219 <= (reg218 ? (7'h4a) : reg86[(3'h5):(1'h0)]);
              reg220 = ((((7'h48) ~^ $signed((wire57 ? wire58 : (7'h45)))) ?
                  wire215[(4'hd):(2'h2)] : (({wire216} ?
                      wire59 : (7'h46)) | ((reg218 <<< reg81) ^ (wire59 == reg62)))) ^~ reg219[(1'h0):(1'h0)]);
            end
          else
            begin
              reg219 <= $signed({reg76, reg81[(4'h8):(3'h5)]});
            end
          reg221 <= reg86[(1'h0):(1'h0)];
          for (forvar222 = (1'h0); (forvar222 < (2'h3)); forvar222 = (forvar222 + (1'h1)))
            begin
              reg223 <= reg67[(2'h3):(2'h2)];
              reg224 <= {{$unsigned($unsigned((forvar217 ? (8'hb6) : wire57))),
                      (($unsigned((8'hb1)) <<< reg86) ?
                          reg88 : (&(reg221 <= (8'hb8))))}};
              reg225 <= forvar217;
              reg226 <= (wire58 == {$signed(reg225)});
              reg227 <= $signed($signed((~^((~reg76) == (|reg68)))));
            end
        end
      reg228 = {(+({(reg85 ? (8'hb2) : reg225), reg223} ?
              reg220[(1'h1):(1'h0)] : {(wire213 ~^ reg76),
                  ((8'hb9) ? wire213 : reg226)}))};
      reg229 <= reg88[(5'h13):(3'h5)];
      if (reg220[(3'h5):(2'h3)])
        begin
          reg230 <= reg226;
          if ((+reg76))
            begin
              reg231 <= (~&$unsigned(wire60[(2'h2):(1'h1)]));
              reg232 = ((^{$signed((reg223 ?
                      reg220 : (8'ha8)))}) <= $unsigned($unsigned($signed((reg68 ^ wire60)))));
              reg233 <= ($signed($unsigned((!$signed(reg227)))) >>> reg223);
              reg234 <= (reg220 ? reg219[(4'hd):(4'ha)] : ((8'ha7) + reg86));
              reg235 = $unsigned({reg220,
                  (((reg67 ? forvar217 : wire58) ~^ reg68[(3'h7):(3'h6)]) ?
                      $signed({forvar222, reg233}) : reg218)});
            end
          else
            begin
              reg231 <= reg220;
              reg233 <= ({$signed($unsigned(reg226[(1'h1):(1'h0)]))} != (7'h47));
              reg234 <= wire57;
              reg235 = ((reg66 >= ((!reg232) >= (8'ha7))) ?
                  (8'ha3) : {$signed(reg228[(3'h4):(3'h4)])});
            end
          reg236 = $signed($signed($signed((~|forvar222[(4'h8):(3'h5)]))));
          reg237 <= (-$signed((~^(((8'ha2) ? reg220 : reg233) ?
              $signed((8'ha8)) : ((8'ha9) ? (8'hb4) : wire57)))));
          if (reg67[(2'h3):(1'h0)])
            begin
              reg238 = (~&reg237);
            end
          else
            begin
              reg238 = $unsigned({((reg223 ? {(8'ha1)} : ((8'hbb) | reg223)) ?
                      (^$unsigned(reg223)) : reg68),
                  ($signed((wire56 ? reg234 : forvar222)) ?
                      forvar222[(2'h3):(1'h0)] : ((!(8'ha1)) ?
                          (wire72 ^~ reg218) : $signed(reg226)))});
            end
        end
      else
        begin
          reg230 <= $signed($signed($unsigned($signed($unsigned(reg66)))));
          if (forvar217[(2'h2):(1'h0)])
            begin
              reg232 = (wire58 ?
                  (reg225 + {(((8'hbe) ? reg221 : (7'h47)) << (wire215 ?
                          (8'ha9) : reg228)),
                      reg218[(5'h12):(3'h5)]}) : (reg229[(1'h1):(1'h0)] >= reg66));
              reg235 = wire215[(5'h12):(3'h5)];
            end
          else
            begin
              reg231 <= ($signed((($unsigned(reg219) || (wire213 || (8'ha5))) ?
                      (^wire56[(4'hb):(4'h8)]) : (-{reg233, wire216}))) ?
                  ((~^$signed($unsigned(reg68))) == reg220) : $unsigned($unsigned(reg66[(4'hd):(1'h1)])));
              reg232 = (~^$unsigned($signed(reg232[(3'h7):(2'h2)])));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module93  (y, clk, wire97, wire96, wire95, wire94);
  output wire [(32'h5b8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire97;
  input wire signed [(5'h18):(1'h0)] wire96;
  input wire [(3'h5):(1'h0)] wire95;
  input wire signed [(4'h9):(1'h0)] wire94;
  wire signed [(4'hc):(1'h0)] wire178;
  wire signed [(4'hf):(1'h0)] wire177;
  wire [(4'ha):(1'h0)] wire176;
  reg signed [(3'h5):(1'h0)] reg199 = (1'h0);
  reg [(4'hb):(1'h0)] reg209 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg208 = (1'h0);
  reg [(2'h3):(1'h0)] reg207 = (1'h0);
  reg signed [(4'he):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg202 = (1'h0);
  reg [(4'hb):(1'h0)] reg200 = (1'h0);
  reg [(5'h11):(1'h0)] reg196 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg194 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg191 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg189 = (1'h0);
  reg [(4'hd):(1'h0)] reg188 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg185 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg182 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg179 = (1'h0);
  reg [(4'hd):(1'h0)] reg171 = (1'h0);
  reg [(5'h18):(1'h0)] reg167 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg161 = (1'h0);
  reg [(4'hc):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg159 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg156 = (1'h0);
  reg [(5'h18):(1'h0)] reg154 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg151 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg150 = (1'h0);
  reg [(4'hb):(1'h0)] reg149 = (1'h0);
  reg [(4'hd):(1'h0)] reg147 = (1'h0);
  reg [(2'h2):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg143 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg142 = (1'h0);
  reg [(3'h4):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg135 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg134 = (1'h0);
  reg [(5'h14):(1'h0)] reg126 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg123 = (1'h0);
  reg [(5'h18):(1'h0)] reg122 = (1'h0);
  reg [(3'h7):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg114 = (1'h0);
  reg [(5'h13):(1'h0)] reg113 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg112 = (1'h0);
  reg [(5'h14):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg109 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg108 = (1'h0);
  reg [(4'h9):(1'h0)] reg107 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg100 = (1'h0);
  reg [(5'h11):(1'h0)] reg212 = (1'h0);
  reg [(2'h2):(1'h0)] reg211 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg206 = (1'h0);
  reg [(3'h5):(1'h0)] reg205 = (1'h0);
  reg [(4'hb):(1'h0)] reg204 = (1'h0);
  reg [(4'hd):(1'h0)] reg201 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar199 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg198 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg197 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg195 = (1'h0);
  reg [(3'h7):(1'h0)] forvar194 = (1'h0);
  reg [(5'h15):(1'h0)] reg193 = (1'h0);
  reg [(4'ha):(1'h0)] reg192 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar187 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg186 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg184 = (1'h0);
  reg signed [(4'he):(1'h0)] reg183 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg181 = (1'h0);
  reg [(3'h7):(1'h0)] reg180 = (1'h0);
  reg [(5'h17):(1'h0)] forvar179 = (1'h0);
  reg [(5'h14):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar174 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg173 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar170 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg169 = (1'h0);
  reg [(5'h13):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg164 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg163 = (1'h0);
  reg [(3'h6):(1'h0)] forvar162 = (1'h0);
  reg [(4'hd):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg157 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg155 = (1'h0);
  reg [(2'h3):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg152 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg146 = (1'h0);
  reg [(5'h15):(1'h0)] forvar144 = (1'h0);
  reg [(4'h8):(1'h0)] reg140 = (1'h0);
  reg [(3'h7):(1'h0)] forvar139 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg137 = (1'h0);
  reg [(5'h15):(1'h0)] reg136 = (1'h0);
  reg [(5'h16):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg132 = (1'h0);
  reg [(3'h5):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg129 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg128 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg124 = (1'h0);
  reg [(5'h16):(1'h0)] reg121 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg120 = (1'h0);
  reg [(3'h6):(1'h0)] forvar117 = (1'h0);
  reg [(3'h4):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar115 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg111 = (1'h0);
  reg [(5'h12):(1'h0)] forvar106 = (1'h0);
  reg [(5'h14):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar99 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar98 = (1'h0);
  assign y = {wire178,
                 wire177,
                 wire176,
                 reg199,
                 reg209,
                 reg208,
                 reg207,
                 reg203,
                 reg202,
                 reg200,
                 reg196,
                 reg194,
                 reg191,
                 reg189,
                 reg188,
                 reg185,
                 reg182,
                 reg179,
                 reg171,
                 reg167,
                 reg166,
                 reg161,
                 reg160,
                 reg159,
                 reg156,
                 reg154,
                 reg151,
                 reg150,
                 reg149,
                 reg147,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg135,
                 reg134,
                 reg126,
                 reg125,
                 reg123,
                 reg122,
                 reg119,
                 reg118,
                 reg114,
                 reg113,
                 reg112,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg105,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg212,
                 reg211,
                 reg210,
                 reg206,
                 reg205,
                 reg204,
                 reg201,
                 forvar199,
                 reg198,
                 reg197,
                 reg195,
                 forvar194,
                 reg193,
                 reg192,
                 reg190,
                 forvar187,
                 reg186,
                 reg184,
                 reg183,
                 reg181,
                 reg180,
                 forvar179,
                 reg175,
                 forvar174,
                 reg173,
                 reg172,
                 forvar170,
                 reg169,
                 reg168,
                 reg165,
                 reg164,
                 reg163,
                 forvar162,
                 reg158,
                 reg157,
                 reg155,
                 reg153,
                 reg152,
                 reg148,
                 reg146,
                 forvar144,
                 reg140,
                 forvar139,
                 reg138,
                 reg137,
                 reg136,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg124,
                 reg121,
                 reg120,
                 forvar117,
                 reg116,
                 forvar115,
                 reg111,
                 forvar106,
                 reg104,
                 forvar99,
                 forvar98,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar98 = (1'h0); (forvar98 < (2'h3)); forvar98 = (forvar98 + (1'h1)))
        begin
          for (forvar99 = (1'h0); (forvar99 < (1'h1)); forvar99 = (forvar99 + (1'h1)))
            begin
              reg100 <= ({(wire95 ?
                          wire97[(4'hb):(2'h3)] : ({wire94,
                              wire95} <<< wire95[(3'h4):(2'h2)]))} ?
                  $signed((~(&$signed(forvar98)))) : wire94);
              reg101 <= $unsigned($signed((+(forvar99 ^~ $signed(wire97)))));
              reg102 <= forvar99;
              reg103 <= (wire96 ?
                  reg101[(1'h1):(1'h1)] : (wire96 ?
                      ($unsigned(forvar98[(3'h6):(1'h0)]) ^ $signed($signed(wire94))) : (((^(8'ha7)) || (~^wire96)) >> wire97)));
            end
          reg104 = (-wire95);
          reg105 <= (~(!$unsigned((forvar98 - (&forvar99)))));
        end
      for (forvar106 = (1'h0); (forvar106 < (2'h2)); forvar106 = (forvar106 + (1'h1)))
        begin
          if (wire97)
            begin
              reg107 <= (wire95[(3'h5):(3'h5)] ?
                  ($signed(reg105) ?
                      (forvar99 ?
                          $signed({(8'ha7),
                              wire95}) : $signed(wire97[(4'hc):(3'h7)])) : (~&{$signed(reg103),
                          (~reg105)})) : $unsigned({$signed({wire95}),
                      forvar106}));
              reg108 <= $signed((({(~|reg101),
                      $signed(reg105)} >> ($signed(forvar106) ?
                      reg101[(1'h1):(1'h0)] : (reg104 > (8'hb9)))) ?
                  (((forvar106 >> reg104) ?
                      $signed(wire96) : $signed(forvar98)) > {wire97,
                      $signed(reg100)}) : $signed(reg100)));
              reg109 <= $signed(((reg101[(3'h5):(1'h0)] >> {reg104[(3'h7):(2'h2)],
                      reg100}) ?
                  forvar106[(4'h9):(3'h6)] : $unsigned(({reg103} ?
                      forvar99 : {(7'h40), wire97}))));
              reg110 <= $signed(reg103[(1'h1):(1'h1)]);
              reg111 = (wire96 + (~|$signed($unsigned((-reg102)))));
            end
          else
            begin
              reg107 <= ($signed(({$unsigned(wire94)} >>> ($unsigned(forvar106) == forvar98))) - $unsigned((^((~&reg108) ?
                  $signed(forvar99) : $signed(reg108)))));
              reg108 <= wire96[(4'hd):(3'h7)];
            end
          reg112 <= (~((|(reg104 ?
              reg109 : reg110[(5'h10):(4'hd)])) >> (^{(8'hb0)})));
          reg113 <= reg104;
          reg114 <= $unsigned($unsigned((reg100[(3'h6):(1'h0)] ?
              $unsigned($signed(wire95)) : forvar98[(1'h1):(1'h1)])));
          for (forvar115 = (1'h0); (forvar115 < (1'h1)); forvar115 = (forvar115 + (1'h1)))
            begin
              reg116 = (reg114 ?
                  $unsigned((~(~$signed(reg100)))) : ({(((8'hab) ?
                                  (8'ha0) : reg100) ?
                              (7'h4a) : $signed((8'ha2))),
                          ({reg104, forvar99} ?
                              (forvar98 ?
                                  reg111 : reg104) : $unsigned(forvar98))} ?
                      reg103[(2'h3):(1'h0)] : reg104[(5'h11):(2'h2)]));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar117 = (1'h0); (forvar117 < (1'h1)); forvar117 = (forvar117 + (1'h1)))
        begin
          if ($unsigned((^~wire94)))
            begin
              reg118 <= ({$signed((~|$unsigned((8'ha4))))} <<< $signed($signed($signed($signed((8'h9e))))));
              reg119 <= ((^(forvar117[(2'h3):(1'h1)] << {$signed(reg110)})) >= reg109);
              reg120 = (!$unsigned(($unsigned({reg102}) > $signed(reg101[(4'hd):(4'hd)]))));
              reg121 = (~^$signed(wire95));
            end
          else
            begin
              reg120 = reg101[(5'h16):(4'ha)];
              reg121 = reg109;
              reg122 <= reg120;
              reg123 <= reg113[(3'h7):(3'h4)];
            end
          reg124 = reg107[(1'h1):(1'h0)];
        end
      if (($unsigned(reg102[(1'h1):(1'h0)]) ?
          $unsigned($unsigned({wire96[(5'h18):(5'h14)]})) : {{($signed(wire94) ?
                      (wire96 - reg110) : $unsigned(wire97))},
              $signed((reg101 ? $signed(reg112) : $unsigned(reg124)))}))
        begin
          if (reg113[(2'h3):(2'h2)])
            begin
              reg125 <= ($signed($unsigned((reg120[(2'h2):(1'h0)] || (forvar117 ~^ reg110)))) ?
                  (!$unsigned($unsigned(reg102))) : ((7'h45) ?
                      $unsigned((~&$signed(reg119))) : (8'hab)));
              reg126 <= wire95[(2'h2):(2'h2)];
              reg127 = {reg103};
            end
          else
            begin
              reg127 = reg102[(3'h5):(1'h1)];
              reg128 = $unsigned(reg127[(2'h2):(1'h0)]);
              reg129 = (8'hb6);
            end
          if (reg100[(3'h5):(1'h0)])
            begin
              reg130 = (^reg105[(1'h1):(1'h0)]);
              reg131 = (~|reg127[(2'h3):(1'h0)]);
              reg132 = $unsigned($signed($signed((~(wire94 + wire94)))));
              reg133 = (!reg131);
            end
          else
            begin
              reg130 = reg131;
              reg131 = reg128;
            end
        end
      else
        begin
          reg125 <= {(!(~&$signed(reg128)))};
          reg126 <= (($signed($unsigned(reg132)) ?
                  reg103 : (((reg127 ? reg122 : reg112) ?
                          {reg131, forvar117} : (reg121 ? reg131 : reg132)) ?
                      reg120 : (reg131 ?
                          reg113[(3'h6):(3'h5)] : $signed(reg129)))) ?
              $signed((reg121 < (((7'h49) ? reg119 : reg100) << {(8'hb2),
                  reg124}))) : $signed((($unsigned((8'h9f)) ?
                  reg123 : $unsigned(reg105)) + $signed((reg122 ?
                  reg103 : wire95)))));
          if ($unsigned($unsigned((reg129[(2'h3):(2'h3)] ?
              $signed($signed((8'hba))) : $unsigned((|reg130))))))
            begin
              reg127 = (($signed((+reg133[(4'h8):(2'h3)])) ?
                      (($unsigned(reg122) <<< $unsigned((7'h41))) >>> (^~$unsigned(reg129))) : {{(!wire97)},
                          (reg102[(3'h5):(2'h3)] <<< (reg122 ?
                              forvar117 : (8'hba)))}) ?
                  {($unsigned({reg132}) ?
                          $unsigned({(7'h46), reg110}) : (((8'ha3) ?
                                  (7'h4a) : reg107) ?
                              wire96[(4'hb):(1'h1)] : (reg118 ?
                                  wire94 : reg108))),
                      (+((~^reg125) ?
                          reg127 : $unsigned(reg105)))} : $signed((reg108[(1'h0):(1'h0)] ?
                      reg120 : ({reg120} - (|(8'ha1))))));
              reg128 = (+wire94[(3'h6):(3'h4)]);
              reg134 <= (~reg120[(3'h5):(1'h1)]);
              reg135 <= reg130[(4'he):(4'ha)];
            end
          else
            begin
              reg127 = reg119;
              reg134 <= $signed({($unsigned(reg113[(4'hc):(4'h9)]) ?
                      reg121 : $unsigned((reg121 ? reg102 : forvar117)))});
              reg135 <= ($signed({($unsigned((8'hba)) - $unsigned(reg103))}) ?
                  ((reg102 ? reg100[(1'h0):(1'h0)] : (&wire96)) ?
                      $unsigned($unsigned((reg123 ?
                          forvar117 : reg122))) : $unsigned(reg119[(2'h2):(1'h0)])) : $unsigned((reg108[(3'h4):(2'h2)] - $signed({reg130}))));
              reg136 = {($signed($unsigned($signed(reg129))) ?
                      (+$unsigned($unsigned(reg126))) : $signed(reg125)),
                  reg131};
              reg137 = ($unsigned(($unsigned($signed(wire96)) ?
                  reg110 : $unsigned((reg102 ?
                      reg128 : reg114)))) << (({$unsigned(reg135)} ?
                      reg136 : $unsigned((~|reg101))) ?
                  reg128 : {reg102, {$signed(reg124), reg102}}));
            end
          reg138 = ((~|((8'hbe) ?
              (reg103 ?
                  $unsigned(reg103) : (reg131 ?
                      wire95 : reg129)) : $signed((reg131 ?
                  wire96 : reg113)))) | $unsigned(reg131));
          for (forvar139 = (1'h0); (forvar139 < (1'h0)); forvar139 = (forvar139 + (1'h1)))
            begin
              reg140 = $signed(reg120[(4'h8):(1'h0)]);
              reg141 <= (+($signed((~^reg109)) ^~ reg100));
              reg142 <= {(^$unsigned((7'h48))), reg137};
              reg143 <= ({$unsigned(wire95[(1'h1):(1'h0)]), reg113} ?
                  (+{(|(reg124 ? reg136 : reg127)),
                      {$signed(reg122)}}) : {reg100[(2'h2):(1'h0)]});
            end
        end
      if (wire95[(2'h2):(1'h0)])
        begin
          reg144 <= (reg105 ?
              $unsigned((($signed(forvar139) > reg107) || reg107)) : reg135);
        end
      else
        begin
          for (forvar144 = (1'h0); (forvar144 < (3'h4)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 <= $signed(reg109[(5'h12):(4'ha)]);
            end
          if ($signed($unsigned((^~reg130[(4'hf):(4'hf)]))))
            begin
              reg146 = reg101;
            end
          else
            begin
              reg147 <= ($signed((+reg146)) ?
                  (($signed($signed(reg110)) ?
                          $unsigned(((8'hac) ^~ reg130)) : $unsigned($unsigned(reg123))) ?
                      {((wire94 ? reg107 : reg146) ?
                              $unsigned((8'h9e)) : (reg114 ? reg138 : reg127)),
                          $unsigned((reg100 ?
                              reg114 : reg146))} : (!reg113)) : $unsigned($unsigned($signed((8'hb3)))));
              reg148 = $signed($unsigned(({(forvar139 >> reg112)} || $unsigned($signed(reg127)))));
              reg149 <= ({($signed(reg128[(1'h1):(1'h1)]) ?
                          reg108[(2'h2):(1'h1)] : ($unsigned(reg134) | (reg105 != wire95)))} ?
                  reg120[(3'h5):(3'h5)] : $unsigned($signed((8'hb5))));
              reg150 <= (^~$unsigned(($unsigned(reg147[(1'h0):(1'h0)]) ?
                  ((8'hb6) < $signed(reg142)) : wire94[(4'h9):(3'h5)])));
              reg151 <= (^~$unsigned(reg119[(3'h4):(2'h3)]));
            end
          reg152 = (({{$unsigned((8'h9f))}, $unsigned($signed(reg121))} ?
                  $unsigned($unsigned((reg109 * reg113))) : $signed({(reg132 != reg118)})) ?
              reg135[(2'h3):(2'h2)] : ($signed(reg126) ?
                  {forvar144} : reg127[(2'h3):(1'h1)]));
          reg153 = $signed($unsigned($signed($signed($unsigned(reg112)))));
          if (reg122)
            begin
              reg154 <= (~|reg148);
              reg155 = ($signed($unsigned((reg141[(2'h3):(2'h2)] ?
                      $unsigned(reg124) : (reg143 ? reg108 : reg145)))) ?
                  reg103[(4'hb):(3'h4)] : (reg143 ?
                      ((reg135 != reg102[(3'h4):(1'h0)]) <= ((forvar117 <<< forvar117) ?
                          (reg125 <<< reg152) : ((8'hb5) ?
                              reg108 : (7'h40)))) : (!(forvar144[(5'h15):(4'he)] ?
                          (!reg144) : (forvar139 + reg107)))));
              reg156 <= $signed({{reg136, $signed({reg142})}});
              reg157 = forvar139[(3'h7):(3'h7)];
              reg158 = (~&{$signed(reg142[(1'h1):(1'h1)]),
                  (+((~|reg142) * (reg141 ? reg105 : reg141)))});
            end
          else
            begin
              reg154 <= ($signed(reg102) & (~^(~reg101)));
              reg156 <= (reg129[(3'h6):(3'h5)] ^ (~(forvar117 ?
                  $unsigned($signed((8'hae))) : (^~(+reg113)))));
              reg159 <= $unsigned((^~wire94[(1'h0):(1'h0)]));
              reg160 <= (!$signed((reg112[(1'h0):(1'h0)] <= (reg124[(5'h11):(4'hc)] ?
                  (~reg149) : reg121))));
              reg161 <= ($signed(forvar144) - ((reg107[(2'h3):(2'h2)] | ((&reg138) ?
                  reg142[(1'h1):(1'h1)] : $unsigned(wire95))) * (($signed(reg159) ~^ reg114) ?
                  reg137 : $signed((+reg140)))));
            end
        end
      if (reg107[(3'h4):(1'h0)])
        begin
          for (forvar162 = (1'h0); (forvar162 < (2'h2)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg163 = reg121;
              reg164 = reg131[(2'h2):(1'h0)];
              reg165 = $signed((reg125[(2'h2):(2'h2)] ^~ {(8'ha0)}));
            end
          reg166 <= (reg142[(2'h3):(2'h2)] > reg105);
          reg167 <= reg148[(3'h4):(1'h0)];
        end
      else
        begin
          for (forvar162 = (1'h0); (forvar162 < (3'h4)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg166 <= (-reg103);
              reg168 = ($signed($unsigned($signed(reg150))) ?
                  (~wire95[(2'h2):(2'h2)]) : reg141);
              reg169 = ((reg112 ?
                      $signed((-{reg149,
                          reg119})) : (+$unsigned($unsigned(reg128)))) ?
                  (~^reg143[(3'h5):(1'h1)]) : reg152);
            end
          for (forvar170 = (1'h0); (forvar170 < (2'h3)); forvar170 = (forvar170 + (1'h1)))
            begin
              reg171 <= reg143;
              reg172 = reg160;
              reg173 = $signed($unsigned(reg152));
            end
          for (forvar174 = (1'h0); (forvar174 < (3'h4)); forvar174 = (forvar174 + (1'h1)))
            begin
              reg175 = $unsigned(reg141[(2'h3):(1'h0)]);
            end
        end
    end
  assign wire176 = ($unsigned($unsigned({$signed(reg145)})) - (reg109[(5'h12):(4'hc)] ^~ (&reg150)));
  assign wire177 = reg156[(4'he):(4'h8)];
  assign wire178 = $unsigned($signed(reg113[(4'he):(4'h9)]));
  always
    @(posedge clk) begin
      if (wire95[(1'h1):(1'h0)])
        begin
          for (forvar179 = (1'h0); (forvar179 < (1'h0)); forvar179 = (forvar179 + (1'h1)))
            begin
              reg180 = $unsigned((($unsigned({reg103}) != (8'ha6)) ?
                  reg118 : $signed(((&reg159) || (~reg171)))));
              reg181 = $signed({{$unsigned($unsigned(reg118)),
                      {$unsigned(reg107)}},
                  ($signed((reg159 ?
                      wire94 : reg105)) - $unsigned($signed((8'ha6))))});
            end
        end
      else
        begin
          if ((~^reg156[(4'hd):(3'h7)]))
            begin
              reg179 <= ((($unsigned({reg150, wire94}) ?
                          ($signed(reg135) ?
                              (reg103 + (8'h9d)) : ((8'ha8) >> reg151)) : (|(~^reg150))) ?
                      reg156 : (reg171[(3'h5):(2'h2)] ? (7'h46) : wire95)) ?
                  $signed({(reg150[(4'h9):(4'h9)] || reg112[(2'h3):(1'h1)])}) : (wire176 >> ((8'haf) ?
                      (&reg154[(4'ha):(1'h0)]) : ((~&wire176) >= reg122))));
              reg182 <= $unsigned((+reg122));
              reg183 = (((&{$unsigned(reg142),
                  ((7'h49) >> reg182)}) ~^ (((~^reg181) ~^ $signed(reg154)) + ({reg166,
                  wire177} != (wire177 + reg141)))) ^ (8'h9c));
              reg184 = forvar179[(5'h13):(4'h8)];
            end
          else
            begin
              reg180 = reg114[(4'hc):(4'hb)];
              reg182 <= $signed(reg181);
              reg183 = $signed(reg151);
              reg184 = ((($signed(((8'ha5) ?
                      wire178 : reg167)) >>> $unsigned(reg154[(3'h6):(1'h1)])) && wire176) ?
                  $signed((8'ha9)) : $unsigned(((8'hb8) ?
                      $signed((reg182 & reg145)) : {reg145[(1'h0):(1'h0)],
                          $unsigned(reg107)})));
              reg185 <= {$signed(reg110),
                  ((($unsigned(reg183) ?
                      $unsigned(wire97) : ((8'h9c) ?
                          forvar179 : reg113)) <<< reg167) ^ ($unsigned((reg145 ?
                          reg171 : (7'h49))) ?
                      ({reg167, reg108} ?
                          (~^reg113) : {(8'hb2),
                              reg108}) : $signed(reg112[(2'h3):(1'h0)])))};
            end
          reg186 = reg185[(1'h0):(1'h0)];
          for (forvar187 = (1'h0); (forvar187 < (2'h3)); forvar187 = (forvar187 + (1'h1)))
            begin
              reg188 <= (+reg144[(5'h13):(3'h6)]);
              reg189 <= $unsigned((-$unsigned((&reg166))));
              reg190 = $unsigned(reg114[(4'hf):(3'h7)]);
              reg191 <= $unsigned((wire178[(4'hb):(3'h6)] ?
                  reg119[(1'h0):(1'h0)] : $signed($unsigned((+reg189)))));
              reg192 = ((((~|(reg189 + reg144)) ?
                          ($signed((8'hab)) ?
                              reg191 : (reg126 <= reg113)) : $unsigned(reg110)) ?
                      (8'hbd) : $unsigned((reg144[(4'hb):(1'h0)] ?
                          (reg105 ? forvar179 : wire96) : {reg181,
                              forvar179}))) ?
                  (7'h42) : reg191);
            end
          reg193 = $unsigned(reg147);
        end
      if (($signed($unsigned((8'had))) >>> reg156))
        begin
          for (forvar194 = (1'h0); (forvar194 < (2'h2)); forvar194 = (forvar194 + (1'h1)))
            begin
              reg195 = reg160[(3'h7):(3'h5)];
            end
        end
      else
        begin
          if ($signed((wire97[(3'h4):(2'h2)] ?
              (($signed(reg145) ? wire97 : (reg142 ? reg192 : reg112)) ?
                  ((^~reg123) ? reg123 : (reg114 >> reg161)) : ({forvar194} ?
                      reg142 : (~|reg195))) : reg190)))
            begin
              reg194 <= {(+reg122[(5'h11):(2'h2)])};
              reg195 = $unsigned(((($signed(reg149) ?
                      $signed(reg143) : (7'h45)) << {wire177, (8'haf)}) ?
                  reg159 : ($unsigned($unsigned(reg135)) >>> {reg105,
                      $unsigned(reg103)})));
              reg196 <= (~|(!forvar194[(3'h6):(1'h1)]));
              reg197 = reg186[(5'h10):(3'h4)];
            end
          else
            begin
              reg195 = $unsigned(reg161[(3'h6):(2'h3)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg198 = $signed(reg141);
      if ((~&$signed((((reg110 ?
          reg102 : (7'h44)) > $signed(reg182)) <<< {wire178[(4'hb):(3'h7)]}))))
        begin
          for (forvar199 = (1'h0); (forvar199 < (1'h0)); forvar199 = (forvar199 + (1'h1)))
            begin
              reg200 <= $unsigned(reg143);
              reg201 = reg167[(4'he):(4'h9)];
              reg202 <= (~|wire96);
            end
          if (reg100[(4'hc):(4'hc)])
            begin
              reg203 <= ($unsigned((($signed(reg191) ^~ forvar199) || $unsigned($unsigned(wire97)))) - (reg150[(4'hc):(4'ha)] * ($unsigned(reg196[(4'h8):(3'h4)]) ?
                  reg202[(2'h2):(1'h0)] : {$signed(reg149)})));
              reg204 = (8'hbb);
            end
          else
            begin
              reg203 <= $signed((reg160 && $unsigned((-reg142[(1'h0):(1'h0)]))));
            end
          if (($signed($signed($signed($signed((7'h44))))) ?
              (^~$signed(({reg159} ?
                  $signed(wire96) : (reg182 && reg147)))) : reg196))
            begin
              reg205 = reg134;
              reg206 = (($unsigned(($signed(wire97) ?
                  (&reg145) : reg122[(4'hf):(3'h7)])) + (reg150 >= $unsigned(reg143[(1'h0):(1'h0)]))) != $signed(reg171[(4'hb):(3'h6)]));
              reg207 <= (~^$unsigned(reg189));
              reg208 <= $signed({$signed(reg194)});
              reg209 <= (8'hac);
            end
          else
            begin
              reg207 <= (8'haa);
            end
        end
      else
        begin
          reg199 <= wire94;
        end
      reg210 = reg126;
      reg211 = (($unsigned((&$unsigned(reg147))) ?
          wire96 : $unsigned(($unsigned(reg147) ?
              reg105 : $unsigned((8'ha0))))) ^~ {(~^$signed((-(8'hac))))});
      reg212 = reg134;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module677  (y, clk, wire682, wire681, wire680, wire679, wire678);
  output wire [(32'hb90):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire682;
  input wire signed [(5'h18):(1'h0)] wire681;
  input wire signed [(4'ha):(1'h0)] wire680;
  input wire signed [(5'h18):(1'h0)] wire679;
  input wire [(5'h11):(1'h0)] wire678;
  wire [(4'h9):(1'h0)] wire799;
  wire [(3'h5):(1'h0)] wire776;
  wire [(4'h8):(1'h0)] wire736;
  wire signed [(3'h5):(1'h0)] wire719;
  reg signed [(3'h6):(1'h0)] reg913 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg912 = (1'h0);
  reg [(5'h17):(1'h0)] reg910 = (1'h0);
  reg [(3'h7):(1'h0)] reg909 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg907 = (1'h0);
  reg [(5'h18):(1'h0)] reg905 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg902 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg901 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg898 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg894 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg891 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg890 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg887 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg884 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg883 = (1'h0);
  reg [(5'h15):(1'h0)] reg882 = (1'h0);
  reg [(3'h6):(1'h0)] reg876 = (1'h0);
  reg [(4'hd):(1'h0)] reg869 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg867 = (1'h0);
  reg [(5'h14):(1'h0)] reg866 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg864 = (1'h0);
  reg [(5'h11):(1'h0)] reg860 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg859 = (1'h0);
  reg [(5'h12):(1'h0)] reg851 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg849 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg848 = (1'h0);
  reg [(3'h6):(1'h0)] reg846 = (1'h0);
  reg [(3'h6):(1'h0)] reg840 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg838 = (1'h0);
  reg [(5'h10):(1'h0)] reg836 = (1'h0);
  reg [(4'hf):(1'h0)] reg835 = (1'h0);
  reg [(4'hd):(1'h0)] reg833 = (1'h0);
  reg [(3'h6):(1'h0)] reg831 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg828 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg826 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg825 = (1'h0);
  reg [(5'h10):(1'h0)] reg821 = (1'h0);
  reg [(5'h12):(1'h0)] reg820 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg813 = (1'h0);
  reg [(2'h3):(1'h0)] reg812 = (1'h0);
  reg [(5'h17):(1'h0)] reg810 = (1'h0);
  reg [(4'hc):(1'h0)] reg808 = (1'h0);
  reg [(5'h16):(1'h0)] reg807 = (1'h0);
  reg [(2'h3):(1'h0)] reg806 = (1'h0);
  reg [(4'ha):(1'h0)] reg800 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg794 = (1'h0);
  reg [(2'h3):(1'h0)] reg792 = (1'h0);
  reg [(5'h14):(1'h0)] reg791 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg790 = (1'h0);
  reg [(3'h4):(1'h0)] reg786 = (1'h0);
  reg signed [(4'he):(1'h0)] reg785 = (1'h0);
  reg [(5'h10):(1'h0)] reg781 = (1'h0);
  reg [(4'hf):(1'h0)] reg773 = (1'h0);
  reg [(4'h9):(1'h0)] reg772 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg768 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg764 = (1'h0);
  reg [(3'h6):(1'h0)] reg763 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg762 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg761 = (1'h0);
  reg [(4'h8):(1'h0)] reg757 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg755 = (1'h0);
  reg [(5'h10):(1'h0)] reg753 = (1'h0);
  reg [(2'h2):(1'h0)] reg752 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg750 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg747 = (1'h0);
  reg [(5'h18):(1'h0)] reg746 = (1'h0);
  reg [(2'h2):(1'h0)] reg743 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg742 = (1'h0);
  reg [(4'hc):(1'h0)] reg741 = (1'h0);
  reg [(4'ha):(1'h0)] reg740 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg735 = (1'h0);
  reg [(2'h2):(1'h0)] reg733 = (1'h0);
  reg [(3'h7):(1'h0)] reg731 = (1'h0);
  reg [(4'hf):(1'h0)] reg728 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg725 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg721 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg718 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg716 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg708 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg695 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg709 = (1'h0);
  reg [(4'he):(1'h0)] reg707 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg705 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg701 = (1'h0);
  reg [(3'h6):(1'h0)] reg699 = (1'h0);
  reg [(4'he):(1'h0)] reg698 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg697 = (1'h0);
  reg [(4'he):(1'h0)] reg694 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg692 = (1'h0);
  reg [(4'he):(1'h0)] reg690 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg687 = (1'h0);
  reg [(3'h6):(1'h0)] reg686 = (1'h0);
  reg [(5'h15):(1'h0)] reg685 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg683 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg914 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg911 = (1'h0);
  reg [(4'h8):(1'h0)] reg908 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg906 = (1'h0);
  reg [(5'h12):(1'h0)] reg904 = (1'h0);
  reg [(4'hf):(1'h0)] forvar903 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg900 = (1'h0);
  reg [(5'h12):(1'h0)] forvar899 = (1'h0);
  reg [(5'h11):(1'h0)] forvar897 = (1'h0);
  reg [(2'h2):(1'h0)] reg895 = (1'h0);
  reg [(5'h10):(1'h0)] reg893 = (1'h0);
  reg [(4'h9):(1'h0)] reg892 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar889 = (1'h0);
  reg [(5'h17):(1'h0)] reg888 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar886 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg885 = (1'h0);
  reg [(5'h17):(1'h0)] reg881 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar880 = (1'h0);
  reg [(5'h13):(1'h0)] reg880 = (1'h0);
  reg [(5'h12):(1'h0)] reg879 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg878 = (1'h0);
  reg [(4'hf):(1'h0)] forvar877 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg875 = (1'h0);
  reg [(5'h13):(1'h0)] reg874 = (1'h0);
  reg [(2'h2):(1'h0)] reg873 = (1'h0);
  reg [(5'h17):(1'h0)] reg872 = (1'h0);
  reg [(3'h6):(1'h0)] reg871 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg870 = (1'h0);
  reg [(5'h12):(1'h0)] reg868 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg865 = (1'h0);
  reg [(5'h11):(1'h0)] forvar863 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg862 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar861 = (1'h0);
  reg [(2'h2):(1'h0)] reg858 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg857 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg856 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg855 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg854 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg853 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar852 = (1'h0);
  reg [(5'h16):(1'h0)] reg850 = (1'h0);
  reg [(5'h12):(1'h0)] forvar829 = (1'h0);
  reg [(4'hf):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg845 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg844 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg843 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar842 = (1'h0);
  reg [(5'h12):(1'h0)] reg841 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg839 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg837 = (1'h0);
  reg [(5'h10):(1'h0)] reg834 = (1'h0);
  reg [(3'h5):(1'h0)] reg832 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg830 = (1'h0);
  reg [(5'h17):(1'h0)] reg829 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg827 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg824 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg823 = (1'h0);
  reg [(2'h2):(1'h0)] reg822 = (1'h0);
  reg [(4'ha):(1'h0)] reg819 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg818 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg817 = (1'h0);
  reg [(4'h9):(1'h0)] reg816 = (1'h0);
  reg [(5'h17):(1'h0)] reg815 = (1'h0);
  reg [(4'hf):(1'h0)] forvar814 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar811 = (1'h0);
  reg signed [(4'he):(1'h0)] reg809 = (1'h0);
  reg [(3'h5):(1'h0)] forvar805 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg804 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg803 = (1'h0);
  reg [(4'he):(1'h0)] reg802 = (1'h0);
  reg [(4'hc):(1'h0)] forvar801 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg798 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg797 = (1'h0);
  reg [(4'hb):(1'h0)] reg796 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar795 = (1'h0);
  reg [(2'h2):(1'h0)] reg793 = (1'h0);
  reg [(3'h5):(1'h0)] reg789 = (1'h0);
  reg [(4'hf):(1'h0)] forvar788 = (1'h0);
  reg [(4'h9):(1'h0)] reg787 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg784 = (1'h0);
  reg [(5'h10):(1'h0)] reg783 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg782 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg780 = (1'h0);
  reg [(3'h7):(1'h0)] reg779 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg778 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg777 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg775 = (1'h0);
  reg [(5'h14):(1'h0)] reg774 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg771 = (1'h0);
  reg [(4'h8):(1'h0)] forvar770 = (1'h0);
  reg signed [(4'he):(1'h0)] reg769 = (1'h0);
  reg [(3'h5):(1'h0)] reg766 = (1'h0);
  reg [(5'h12):(1'h0)] reg765 = (1'h0);
  reg [(5'h16):(1'h0)] reg760 = (1'h0);
  reg [(4'he):(1'h0)] forvar759 = (1'h0);
  reg [(4'hf):(1'h0)] forvar758 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg756 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg754 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg751 = (1'h0);
  reg [(5'h17):(1'h0)] reg749 = (1'h0);
  reg [(5'h10):(1'h0)] forvar748 = (1'h0);
  reg [(3'h7):(1'h0)] reg745 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg744 = (1'h0);
  reg [(5'h16):(1'h0)] reg739 = (1'h0);
  reg [(5'h12):(1'h0)] forvar738 = (1'h0);
  reg [(3'h6):(1'h0)] forvar737 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg734 = (1'h0);
  reg [(3'h4):(1'h0)] reg732 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg730 = (1'h0);
  reg [(4'hf):(1'h0)] reg729 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg727 = (1'h0);
  reg [(4'h9):(1'h0)] forvar726 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg724 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg723 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg722 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg720 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg717 = (1'h0);
  reg [(4'hd):(1'h0)] reg715 = (1'h0);
  reg [(3'h6):(1'h0)] forvar714 = (1'h0);
  reg [(4'h9):(1'h0)] forvar713 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg712 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar694 = (1'h0);
  reg [(5'h15):(1'h0)] reg689 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg711 = (1'h0);
  reg [(3'h5):(1'h0)] reg710 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar708 = (1'h0);
  reg [(4'hd):(1'h0)] reg706 = (1'h0);
  reg [(5'h14):(1'h0)] reg704 = (1'h0);
  reg [(4'h9):(1'h0)] reg702 = (1'h0);
  reg signed [(4'he):(1'h0)] reg700 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg696 = (1'h0);
  reg [(5'h15):(1'h0)] forvar695 = (1'h0);
  reg [(4'h9):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg691 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar689 = (1'h0);
  reg [(4'ha):(1'h0)] reg688 = (1'h0);
  reg [(3'h7):(1'h0)] reg684 = (1'h0);
  assign y = {wire799,
                 wire776,
                 wire736,
                 wire719,
                 reg913,
                 reg912,
                 reg910,
                 reg909,
                 reg907,
                 reg905,
                 reg902,
                 reg901,
                 reg898,
                 reg896,
                 reg894,
                 reg891,
                 reg890,
                 reg887,
                 reg884,
                 reg883,
                 reg882,
                 reg876,
                 reg869,
                 reg867,
                 reg866,
                 reg864,
                 reg860,
                 reg859,
                 reg851,
                 reg849,
                 reg848,
                 reg846,
                 reg840,
                 reg838,
                 reg836,
                 reg835,
                 reg833,
                 reg831,
                 reg828,
                 reg826,
                 reg825,
                 reg821,
                 reg820,
                 reg813,
                 reg812,
                 reg810,
                 reg808,
                 reg807,
                 reg806,
                 reg800,
                 reg794,
                 reg792,
                 reg791,
                 reg790,
                 reg786,
                 reg785,
                 reg781,
                 reg773,
                 reg772,
                 reg768,
                 reg767,
                 reg764,
                 reg763,
                 reg762,
                 reg761,
                 reg757,
                 reg755,
                 reg753,
                 reg752,
                 reg750,
                 reg747,
                 reg746,
                 reg743,
                 reg742,
                 reg741,
                 reg740,
                 reg735,
                 reg733,
                 reg731,
                 reg728,
                 reg725,
                 reg721,
                 reg718,
                 reg716,
                 reg708,
                 reg695,
                 reg709,
                 reg707,
                 reg705,
                 reg703,
                 reg701,
                 reg699,
                 reg698,
                 reg697,
                 reg694,
                 reg692,
                 reg690,
                 reg687,
                 reg686,
                 reg685,
                 reg683,
                 reg914,
                 reg911,
                 reg908,
                 reg906,
                 reg904,
                 forvar903,
                 reg900,
                 forvar899,
                 forvar897,
                 reg895,
                 reg893,
                 reg892,
                 forvar889,
                 reg888,
                 forvar886,
                 reg885,
                 reg881,
                 forvar880,
                 reg880,
                 reg879,
                 reg878,
                 forvar877,
                 reg875,
                 reg874,
                 reg873,
                 reg872,
                 reg871,
                 reg870,
                 reg868,
                 reg865,
                 forvar863,
                 reg862,
                 forvar861,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 forvar852,
                 reg850,
                 forvar829,
                 reg847,
                 reg845,
                 reg844,
                 reg843,
                 forvar842,
                 reg841,
                 reg839,
                 reg837,
                 reg834,
                 reg832,
                 reg830,
                 reg829,
                 reg827,
                 reg824,
                 reg823,
                 reg822,
                 reg819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 forvar814,
                 forvar811,
                 reg809,
                 forvar805,
                 reg804,
                 reg803,
                 reg802,
                 forvar801,
                 reg798,
                 reg797,
                 reg796,
                 forvar795,
                 reg793,
                 reg789,
                 forvar788,
                 reg787,
                 reg784,
                 reg783,
                 reg782,
                 reg780,
                 reg779,
                 reg778,
                 reg777,
                 reg775,
                 reg774,
                 reg771,
                 forvar770,
                 reg769,
                 reg766,
                 reg765,
                 reg760,
                 forvar759,
                 forvar758,
                 reg756,
                 reg754,
                 reg751,
                 reg749,
                 forvar748,
                 reg745,
                 reg744,
                 reg739,
                 forvar738,
                 forvar737,
                 reg734,
                 reg732,
                 reg730,
                 reg729,
                 reg727,
                 forvar726,
                 reg724,
                 reg723,
                 reg722,
                 reg720,
                 reg717,
                 reg715,
                 forvar714,
                 forvar713,
                 reg712,
                 forvar694,
                 reg689,
                 reg711,
                 reg710,
                 forvar708,
                 reg706,
                 reg704,
                 reg702,
                 reg700,
                 reg696,
                 forvar695,
                 reg693,
                 reg691,
                 forvar689,
                 reg688,
                 reg684,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned(wire679[(3'h5):(2'h3)]))
        begin
          if (wire679[(4'h9):(1'h1)])
            begin
              reg683 <= ($signed((wire680 > wire678[(2'h3):(2'h3)])) == wire680[(1'h1):(1'h0)]);
            end
          else
            begin
              reg684 = $signed({$signed($unsigned((reg683 ^~ wire680)))});
              reg685 <= (wire678[(4'h9):(2'h2)] ?
                  (wire681 ?
                      (~(reg683[(1'h1):(1'h0)] + $signed(wire682))) : (+((reg684 ?
                              wire681 : wire681) ?
                          reg684[(2'h3):(2'h3)] : $unsigned(reg684)))) : $signed((wire681 ?
                      reg684[(3'h6):(3'h4)] : wire679)));
              reg686 <= ((reg685 ^~ (((wire678 >>> wire681) ?
                      wire678[(4'he):(4'ha)] : (~&reg684)) ?
                  {$unsigned(reg683)} : {$unsigned(wire680)})) + $unsigned((($unsigned(wire681) ?
                      wire678 : $unsigned(wire678)) ?
                  reg684 : ((-reg684) > reg685[(5'h11):(4'ha)]))));
              reg687 <= (^((~|(wire682[(4'hf):(3'h4)] ?
                  $unsigned(reg683) : wire678[(4'h9):(3'h6)])) >= wire681[(4'he):(4'hd)]));
              reg688 = $unsigned((wire680[(2'h2):(1'h1)] ?
                  (^~((+wire680) ?
                      {reg685} : $unsigned(wire679))) : $unsigned((-wire678[(1'h0):(1'h0)]))));
            end
        end
      else
        begin
          reg683 <= wire682[(4'hc):(4'h9)];
        end
      if ((^~(~&wire682[(3'h6):(1'h1)])))
        begin
          for (forvar689 = (1'h0); (forvar689 < (1'h0)); forvar689 = (forvar689 + (1'h1)))
            begin
              reg690 <= ($unsigned(wire680[(4'h9):(1'h1)]) ?
                  (~^$unsigned(reg684[(3'h7):(2'h2)])) : reg688);
              reg691 = (((^~reg686[(2'h2):(2'h2)]) ?
                  $unsigned(forvar689[(4'h8):(3'h7)]) : (&$unsigned((wire679 ^ wire682)))) && $unsigned($signed(reg685)));
              reg692 <= {(+wire679), $signed({(~^$signed(wire678))})};
              reg693 = $unsigned(wire682);
              reg694 <= (~|((((reg691 < wire682) <<< $unsigned(reg683)) ?
                      ((~&wire679) != ((8'ha1) ?
                          reg686 : reg690)) : $signed(reg691[(3'h5):(2'h2)])) ?
                  reg683[(2'h2):(1'h1)] : (($signed(reg688) << (8'hb2)) ?
                      (8'h9c) : (~&$unsigned(reg686)))));
            end
          for (forvar695 = (1'h0); (forvar695 < (1'h1)); forvar695 = (forvar695 + (1'h1)))
            begin
              reg696 = reg687;
              reg697 <= ((~((reg692[(1'h0):(1'h0)] & wire681) || $unsigned((wire678 >= forvar689)))) ?
                  ($unsigned((reg683[(3'h6):(3'h5)] < (+wire681))) ?
                      reg694 : (~^$unsigned($unsigned(reg687)))) : reg690);
              reg698 <= (~&(~(($unsigned(wire679) & $signed(forvar689)) < $signed((reg691 + reg688)))));
              reg699 <= reg690;
              reg700 = (~|wire679[(4'hc):(2'h3)]);
            end
          if (($signed($unsigned($signed(reg691))) != ($signed({((7'h4a) ?
                  wire678 : (8'h9d))}) ~^ forvar695[(4'h9):(4'h9)])))
            begin
              reg701 <= {$signed(reg687[(4'hc):(3'h5)]),
                  (^(&(wire678 ? reg684 : (reg692 || reg683))))};
              reg702 = wire680;
              reg703 <= $signed($unsigned((-((wire678 ?
                  wire682 : reg697) >> (wire679 * wire682)))));
              reg704 = (!$unsigned((8'hb3)));
            end
          else
            begin
              reg701 <= (+{(reg697 ?
                      reg687[(4'hf):(1'h1)] : ((reg690 ?
                          reg696 : reg696) < reg700))});
              reg702 = $unsigned(((~|reg692) * (($unsigned(reg687) ?
                  ((7'h49) && wire680) : $signed((7'h43))) <= (+(wire680 ?
                  wire679 : reg692)))));
              reg704 = ((8'h9c) + reg685);
              reg705 <= $signed($signed($unsigned((~|(&reg687)))));
            end
          if ($unsigned(reg698))
            begin
              reg706 = reg687;
              reg707 <= $signed((($unsigned($unsigned(reg691)) + reg700[(1'h1):(1'h1)]) * $signed((~^reg696[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg707 <= wire680[(1'h0):(1'h0)];
            end
          for (forvar708 = (1'h0); (forvar708 < (2'h2)); forvar708 = (forvar708 + (1'h1)))
            begin
              reg709 <= ((|(~|reg684)) ?
                  $unsigned((-$unsigned((reg705 ?
                      forvar708 : reg684)))) : (-wire682[(2'h2):(2'h2)]));
              reg710 = $signed($unsigned((+reg687[(3'h4):(1'h1)])));
              reg711 = {$signed(reg693)};
            end
        end
      else
        begin
          reg689 = reg711;
          if ((((|reg693) ?
                  reg691 : {(reg703[(4'hb):(2'h3)] ?
                          (!reg689) : (forvar708 != reg692)),
                      reg685[(2'h3):(1'h1)]}) ?
              (($signed((wire680 ?
                      forvar708 : (8'hae))) <<< ((|reg697) ^ (forvar689 >> reg707))) ?
                  $signed($signed(forvar695)) : reg693) : reg710))
            begin
              reg691 = ($unsigned(($signed({reg687, reg710}) <= $signed({reg703,
                      (7'h49)}))) ?
                  $signed(reg706[(2'h2):(1'h1)]) : $signed((^({wire680,
                      reg709} - (!reg696)))));
              reg693 = $unsigned($signed((^{(forvar695 > reg711),
                  (wire681 ? forvar708 : (8'ha2))})));
            end
          else
            begin
              reg691 = $unsigned($signed(({reg709,
                  reg700[(3'h4):(3'h4)]} || (!reg703))));
            end
          for (forvar694 = (1'h0); (forvar694 < (1'h1)); forvar694 = (forvar694 + (1'h1)))
            begin
              reg695 <= (^reg709[(2'h2):(1'h0)]);
              reg697 <= reg706;
              reg700 = $signed(reg698);
              reg702 = wire679;
              reg703 <= (~(forvar708 ?
                  {$signed((forvar708 ?
                          reg711 : (8'h9d)))} : reg683[(3'h4):(1'h0)]));
            end
          reg704 = {reg683};
          if (reg711[(1'h0):(1'h0)])
            begin
              reg705 <= (7'h47);
              reg707 <= {{reg710}};
              reg708 <= $unsigned(reg694[(3'h6):(2'h2)]);
            end
          else
            begin
              reg706 = ($unsigned((reg703[(3'h6):(1'h0)] ?
                      (~forvar689) : reg695)) ?
                  ($signed((8'hba)) < (^reg704[(4'h8):(4'h8)])) : reg691[(1'h0):(1'h0)]);
              reg707 <= ((($unsigned(reg693) ?
                  forvar689 : reg695[(1'h0):(1'h0)]) && ($unsigned($signed(reg684)) + $unsigned({reg692,
                  wire681}))) && (~^reg688));
              reg708 <= wire682;
              reg709 <= (~|$unsigned($unsigned($unsigned(reg704[(5'h12):(2'h3)]))));
            end
        end
      reg712 = (((($unsigned(wire682) + $signed((8'hbe))) ?
              (((8'hbe) == reg689) ?
                  (reg711 - reg702) : reg695) : (8'hb6)) + (-forvar695)) ?
          $signed(reg685[(4'hf):(3'h7)]) : (!reg707));
      for (forvar713 = (1'h0); (forvar713 < (2'h3)); forvar713 = (forvar713 + (1'h1)))
        begin
          for (forvar714 = (1'h0); (forvar714 < (1'h0)); forvar714 = (forvar714 + (1'h1)))
            begin
              reg715 = $unsigned((~forvar694[(5'h13):(5'h11)]));
            end
          reg716 <= ($signed(reg690) >>> ((^((+reg688) ?
              {reg688,
                  reg691} : (forvar713 && reg685))) == $unsigned(wire679)));
          reg717 = ((reg704[(3'h6):(3'h4)] ^ ({$unsigned(reg704),
              $unsigned(forvar714)} * (7'h44))) ^~ $signed((~|$signed((-forvar713)))));
          reg718 <= reg717;
        end
    end
  assign wire719 = (reg692[(3'h4):(2'h3)] - reg708);
  always
    @(posedge clk) begin
      reg720 = reg708;
      if ({(({$signed(wire679)} ?
              reg705[(1'h1):(1'h1)] : $signed(reg695[(3'h4):(1'h1)])) < wire719[(2'h3):(2'h2)])})
        begin
          reg721 <= reg709;
        end
      else
        begin
          if ($unsigned(reg686[(1'h0):(1'h0)]))
            begin
              reg722 = $signed(((+$signed($signed(reg708))) >= (+(^~(reg703 > reg709)))));
              reg723 = reg716[(3'h4):(2'h3)];
              reg724 = $signed((7'h40));
            end
          else
            begin
              reg722 = reg720[(1'h1):(1'h0)];
              reg725 <= (-$signed($unsigned(((reg718 < reg690) && (reg705 + wire679)))));
            end
          for (forvar726 = (1'h0); (forvar726 < (3'h4)); forvar726 = (forvar726 + (1'h1)))
            begin
              reg727 = reg698[(2'h2):(1'h1)];
              reg728 <= (((reg692[(1'h1):(1'h1)] < $signed((~&reg725))) << $signed(reg694)) ^ ((((reg725 ?
                      reg718 : (8'hac)) << {wire680,
                      reg720}) <= $signed(((8'haf) ? wire682 : reg699))) ?
                  $unsigned((wire679 <<< (reg707 >> wire680))) : (|$unsigned(((8'hb1) ?
                      reg686 : reg683)))));
            end
          reg729 = $unsigned($signed(((!reg716[(1'h1):(1'h1)]) ?
              reg685[(1'h0):(1'h0)] : {{reg724}, {reg694}})));
          if ($signed({wire682[(1'h1):(1'h1)], forvar726}))
            begin
              reg730 = $unsigned(wire678);
            end
          else
            begin
              reg730 = reg722;
              reg731 <= reg685[(5'h10):(2'h2)];
              reg732 = $signed($signed($unsigned((-(|wire681)))));
              reg733 <= ((~&(-(+$signed(reg685)))) ?
                  $signed(reg699[(1'h0):(1'h0)]) : reg725[(4'hc):(4'h8)]);
              reg734 = $unsigned((-(8'h9f)));
            end
          reg735 <= (reg690[(2'h3):(1'h0)] & forvar726[(1'h0):(1'h0)]);
        end
    end
  assign wire736 = {(8'h9f)};
  always
    @(posedge clk) begin
      for (forvar737 = (1'h0); (forvar737 < (2'h3)); forvar737 = (forvar737 + (1'h1)))
        begin
          for (forvar738 = (1'h0); (forvar738 < (3'h4)); forvar738 = (forvar738 + (1'h1)))
            begin
              reg739 = ((-$unsigned(wire681[(3'h6):(1'h1)])) ?
                  reg690[(1'h1):(1'h1)] : reg699);
              reg740 <= (~|$signed(reg739));
              reg741 <= ({reg709, reg699[(1'h0):(1'h0)]} >> (^~$signed((reg692 ?
                  ((8'hae) ? wire680 : reg731) : reg709))));
              reg742 <= ((reg697[(2'h2):(1'h0)] ?
                  (reg735 ~^ reg741) : ((!$unsigned((8'hb9))) << ((~&wire736) ^~ $unsigned(wire678)))) < (|(({reg739} ?
                  $unsigned(reg721) : reg687) >> (!reg705[(2'h3):(1'h1)]))));
            end
          if ($signed(($unsigned(wire680) ?
              (|($signed(reg728) ^ (reg733 ?
                  reg733 : reg709))) : $unsigned($signed({wire678, reg683})))))
            begin
              reg743 <= $unsigned($unsigned(((((8'hb5) >> reg705) + (reg721 ?
                      (8'hb9) : wire736)) ?
                  reg718 : ((forvar738 & wire736) ?
                      (-wire678) : (reg709 + wire719)))));
              reg744 = (((($unsigned(wire736) <= (^~reg725)) ?
                      reg685[(4'hd):(2'h2)] : reg695[(1'h1):(1'h0)]) ?
                  {reg716[(1'h1):(1'h1)]} : reg687) <= reg743[(2'h2):(2'h2)]);
              reg745 = reg744;
              reg746 <= wire679;
              reg747 <= (((~^({forvar738} ? (reg694 ^ reg685) : (~|(8'hb5)))) ?
                      ((^reg699[(2'h3):(1'h0)]) ?
                          (-(^~reg731)) : reg741[(4'h8):(2'h3)]) : {($unsigned((8'ha4)) != (wire679 < (8'ha6)))}) ?
                  (7'h43) : $signed((&reg741[(4'h8):(2'h3)])));
            end
          else
            begin
              reg744 = $signed(reg707[(4'h8):(3'h4)]);
            end
          for (forvar748 = (1'h0); (forvar748 < (3'h4)); forvar748 = (forvar748 + (1'h1)))
            begin
              reg749 = $unsigned((~$unsigned($signed({reg685}))));
              reg750 <= $signed(reg701);
              reg751 = (+reg716);
            end
          if ({reg733[(2'h2):(1'h0)], $signed(reg735)})
            begin
              reg752 <= reg695;
              reg753 <= (8'ha2);
            end
          else
            begin
              reg754 = (~reg690[(4'hd):(3'h7)]);
            end
          reg755 <= $unsigned($signed((&(!$unsigned(wire679)))));
        end
      reg756 = (reg716[(3'h4):(1'h1)] ?
          (reg745 & $unsigned(($signed(wire719) && (^forvar737)))) : $signed(forvar737[(1'h0):(1'h0)]));
      reg757 <= forvar737;
      for (forvar758 = (1'h0); (forvar758 < (1'h0)); forvar758 = (forvar758 + (1'h1)))
        begin
          for (forvar759 = (1'h0); (forvar759 < (3'h4)); forvar759 = (forvar759 + (1'h1)))
            begin
              reg760 = ({reg756[(1'h1):(1'h1)]} & $unsigned((8'haf)));
              reg761 <= $signed(reg690);
              reg762 <= {(^(+$unsigned(reg690[(4'hb):(3'h5)])))};
              reg763 <= reg718[(1'h1):(1'h0)];
            end
          if ($unsigned((($unsigned((&reg731)) + (((8'ha7) ? reg695 : reg754) ?
              {reg753} : ((8'ha8) ^~ reg687))) >= (~|reg761[(2'h2):(1'h0)]))))
            begin
              reg764 <= (|$signed($unsigned(({wire680} >> reg721))));
              reg765 = (~&$signed($signed(reg735)));
              reg766 = ((8'hb1) >> ((((~^reg733) ~^ (wire680 ?
                      reg698 : reg747)) <= $signed($unsigned(reg705))) ?
                  $unsigned((^$signed(reg742))) : (((reg718 ?
                          reg760 : reg701) * $unsigned((7'h46))) ?
                      forvar758[(1'h1):(1'h1)] : (8'ha3))));
              reg767 <= ($signed((reg747[(2'h3):(2'h2)] ?
                  ((wire678 ? reg701 : wire719) ?
                      reg756 : $signed(reg705)) : (^~reg749))) >= forvar758[(4'hd):(3'h6)]);
            end
          else
            begin
              reg765 = $unsigned(forvar737);
              reg767 <= $signed((((~&(reg685 ?
                  reg703 : (8'hb8))) + reg756[(4'h9):(3'h7)]) == $signed(reg718)));
              reg768 <= (($unsigned(reg709[(2'h2):(1'h0)]) ?
                  $signed((reg683[(4'hb):(3'h4)] ?
                      (~^reg721) : reg685[(2'h3):(2'h2)])) : $unsigned($unsigned(((8'hb5) - reg764)))) ^~ ((-reg747) & {((~^reg764) + ((8'hb2) - reg754)),
                  {(reg686 >>> reg685), (8'ha2)}}));
              reg769 = ($signed((((!reg743) ?
                          (wire719 ? reg739 : wire682) : (reg686 ?
                              reg750 : (8'ha0))) ?
                      ($unsigned(reg763) > (reg741 >>> reg761)) : ((wire679 < reg751) ?
                          (reg716 >>> forvar737) : reg747[(1'h0):(1'h0)]))) ?
                  $unsigned($signed(reg690)) : $unsigned((reg751[(3'h6):(1'h1)] ^~ $signed({reg683}))));
            end
          for (forvar770 = (1'h0); (forvar770 < (1'h1)); forvar770 = (forvar770 + (1'h1)))
            begin
              reg771 = reg761[(2'h2):(1'h0)];
              reg772 <= $unsigned(((reg725[(1'h1):(1'h1)] ? reg755 : reg753) ?
                  $signed($signed((reg735 * reg767))) : $unsigned((reg741 ?
                      (reg746 ? reg733 : reg747) : wire682[(5'h10):(1'h0)]))));
              reg773 <= reg692[(1'h0):(1'h0)];
              reg774 = reg728;
            end
        end
      reg775 = $unsigned(forvar759[(4'hc):(1'h0)]);
    end
  assign wire776 = reg764;
  always
    @(posedge clk) begin
      if ({(8'hb7)})
        begin
          reg777 = (8'hba);
          reg778 = reg716;
          if (reg735)
            begin
              reg779 = (({$signed((-reg755)),
                          $unsigned(wire682[(4'hb):(3'h5)])} ?
                      $signed(reg697[(2'h2):(1'h0)]) : reg747) ?
                  (~^$signed($signed(reg686[(1'h1):(1'h1)]))) : $unsigned((!$unsigned(reg773[(4'h8):(3'h5)]))));
              reg780 = (reg698 - (&$unsigned({reg731[(3'h5):(2'h2)]})));
            end
          else
            begin
              reg779 = reg698;
            end
          if (reg690)
            begin
              reg781 <= $signed(reg695[(1'h1):(1'h0)]);
            end
          else
            begin
              reg782 = $unsigned(($unsigned(reg708) ?
                  (($signed(reg752) >>> $signed(reg779)) ^ $unsigned({(8'hbc),
                      reg692})) : reg780));
              reg783 = (wire679[(4'he):(3'h5)] + reg683);
            end
          if ($signed(reg777[(1'h1):(1'h0)]))
            begin
              reg784 = $unsigned((^~$unsigned((~|(~|wire681)))));
              reg785 <= reg784;
            end
          else
            begin
              reg784 = (($signed((~|reg773[(4'hd):(4'h8)])) - $unsigned($signed(reg778[(1'h1):(1'h1)]))) || (reg705 ?
                  $unsigned(reg731) : {((!wire719) & (7'h40))}));
              reg785 <= reg683;
              reg786 <= ((~$signed(wire736[(3'h4):(2'h3)])) ?
                  $unsigned($signed($signed(reg683))) : wire736);
            end
        end
      else
        begin
          if ((8'hb4))
            begin
              reg781 <= reg764[(2'h3):(1'h1)];
              reg782 = (~^{(|wire678[(1'h1):(1'h0)])});
            end
          else
            begin
              reg777 = $signed(((&((|reg692) && reg697[(2'h2):(2'h2)])) ?
                  ($signed(wire719[(1'h0):(1'h0)]) + (7'h48)) : ($signed((wire736 ?
                      reg772 : wire776)) == reg772[(3'h4):(3'h4)])));
              reg781 <= $unsigned({(-(((8'haa) ? wire678 : reg705) > (8'hac))),
                  $signed($unsigned((reg698 ? reg716 : reg699)))});
              reg782 = (7'h40);
              reg783 = $signed($unsigned({reg685, $unsigned((8'hab))}));
              reg784 = (reg728 ?
                  $unsigned(((^~reg725[(2'h3):(2'h2)]) ?
                      reg687 : (reg718 + $unsigned(reg701)))) : (~|{(!(^wire681))}));
            end
          reg787 = (~&reg694[(2'h3):(1'h1)]);
          for (forvar788 = (1'h0); (forvar788 < (1'h1)); forvar788 = (forvar788 + (1'h1)))
            begin
              reg789 = ((reg701 ?
                      (~^((+reg773) + reg747)) : $signed(($unsigned(reg699) > $unsigned(forvar788)))) ?
                  $unsigned(($unsigned((!reg746)) ?
                      $signed((reg743 ?
                          reg733 : (7'h40))) : $unsigned((reg694 <<< reg753)))) : (&reg781[(3'h4):(2'h2)]));
              reg790 <= reg782;
              reg791 <= (8'h9d);
              reg792 <= (reg707 <= $unsigned(((~^wire736) - $signed($unsigned((8'haa))))));
            end
          reg793 = (reg780[(3'h7):(3'h4)] >>> (reg697[(2'h3):(2'h2)] >>> {{(reg755 ?
                      reg755 : reg694),
                  (+reg705)},
              ($signed(reg742) <= reg694)}));
          reg794 <= (~^$signed(forvar788));
        end
      for (forvar795 = (1'h0); (forvar795 < (1'h1)); forvar795 = (forvar795 + (1'h1)))
        begin
          reg796 = wire678[(3'h7):(1'h0)];
        end
      reg797 = reg753[(4'hb):(3'h7)];
      reg798 = reg708;
    end
  assign wire799 = ((reg716[(1'h0):(1'h0)] < reg792[(2'h3):(2'h2)]) <<< {(((reg683 == reg707) ?
                               reg781 : $unsigned(wire776)) ?
                           $unsigned(reg767) : $signed((&reg753))),
                       (^$unsigned((wire681 >= (8'hb5))))});
  always
    @(posedge clk) begin
      reg800 <= ($unsigned({{reg757, $signed(reg686)},
              wire776[(3'h5):(2'h2)]}) ?
          reg764[(3'h4):(1'h0)] : reg685);
      for (forvar801 = (1'h0); (forvar801 < (1'h0)); forvar801 = (forvar801 + (1'h1)))
        begin
          reg802 = $signed((($unsigned($unsigned(reg785)) != $unsigned(((8'hac) >= wire678))) ?
              (7'h45) : reg755));
          reg803 = reg772;
          reg804 = wire681[(3'h7):(3'h4)];
          for (forvar805 = (1'h0); (forvar805 < (2'h3)); forvar805 = (forvar805 + (1'h1)))
            begin
              reg806 <= reg716[(1'h1):(1'h1)];
            end
          if ((~(-($unsigned($unsigned(reg725)) || $signed({reg750})))))
            begin
              reg807 <= wire678[(3'h7):(2'h2)];
              reg808 <= {(8'hb0), (^~(reg728[(2'h3):(2'h3)] >= reg794))};
              reg809 = (8'hae);
            end
          else
            begin
              reg807 <= reg763;
            end
        end
      reg810 <= reg802[(4'ha):(1'h1)];
      for (forvar811 = (1'h0); (forvar811 < (3'h4)); forvar811 = (forvar811 + (1'h1)))
        begin
          reg812 <= wire736;
          reg813 <= ($unsigned($unsigned((~&{reg746}))) ?
              $signed($unsigned({(^~reg701), reg705})) : $signed((reg716 ?
                  (~&{reg690, (8'hb0)}) : reg728[(4'hb):(3'h5)])));
          for (forvar814 = (1'h0); (forvar814 < (2'h3)); forvar814 = (forvar814 + (1'h1)))
            begin
              reg815 = (($unsigned(($signed(reg728) ?
                      (+wire682) : $signed(reg683))) ?
                  reg698 : {(7'h46)}) != reg747);
              reg816 = ($unsigned({$unsigned($unsigned(reg792))}) == reg762);
              reg817 = (reg699 ?
                  (|(~^reg743)) : (reg752[(2'h2):(2'h2)] - $signed(((^reg815) + ((7'h41) ?
                      wire719 : reg747)))));
              reg818 = $signed(reg683);
            end
          if (reg750)
            begin
              reg819 = ($signed($signed((~|(reg728 ? reg817 : reg735)))) ?
                  reg804[(4'h8):(3'h7)] : (~|$unsigned((~(-reg755)))));
              reg820 <= $unsigned({$signed(((reg813 ?
                      reg703 : (8'h9c)) << (wire680 ~^ (8'h9d)))),
                  ($unsigned((reg686 ? wire682 : reg772)) ?
                      reg786 : $unsigned((|reg692)))});
              reg821 <= reg763;
            end
          else
            begin
              reg819 = $signed((reg740[(4'ha):(3'h5)] ?
                  {$unsigned(reg803),
                      ($signed(reg753) ? reg694 : (~forvar801))} : forvar805));
              reg822 = ($signed(reg820[(1'h0):(1'h0)]) || ((&reg755) ?
                  $unsigned(((wire776 ~^ (8'hb3)) ^~ reg816[(1'h0):(1'h0)])) : $unsigned(((reg731 == reg741) ?
                      reg721 : (&reg818)))));
              reg823 = reg822[(1'h1):(1'h0)];
              reg824 = $signed(reg815[(2'h3):(1'h0)]);
            end
          reg825 <= {reg694[(4'hd):(4'hb)],
              (~^(reg747 ?
                  ((reg752 || reg683) ?
                      (reg687 ?
                          reg716 : reg753) : (reg735 > reg708)) : $unsigned($unsigned(reg803))))};
        end
    end
  always
    @(posedge clk) begin
      if (((((+(-reg755)) ?
                  reg735 : (((8'ha3) ~^ reg768) ?
                      reg762[(1'h0):(1'h0)] : reg768[(2'h2):(2'h2)])) ?
              (~|(8'hb9)) : $unsigned(reg792[(2'h2):(1'h1)])) ?
          {$signed(reg701),
              (reg718[(1'h0):(1'h0)] ?
                  reg692 : (reg728[(2'h2):(2'h2)] ?
                      ((8'hbf) != reg753) : reg761[(1'h0):(1'h0)]))} : (-(+reg709[(2'h2):(2'h2)]))))
        begin
          reg826 <= ((8'haf) ?
              {{((reg705 ? reg683 : reg708) ? $unsigned(reg785) : wire799),
                      $unsigned((reg773 ?
                          wire679 : reg692))}} : $signed(reg742));
        end
      else
        begin
          reg827 = (8'h9f);
          reg828 <= wire682;
        end
      if (({($signed((wire736 ? reg683 : reg705)) ?
              reg694 : $unsigned((~|(8'haa)))),
          (($unsigned(reg810) ?
              (reg690 ~^ reg772) : (reg699 ?
                  reg742 : (8'hba))) | (~&(reg708 >>> reg791)))} == reg808))
        begin
          if (reg806)
            begin
              reg829 = (~|reg687[(4'he):(3'h5)]);
              reg830 = wire680[(2'h3):(2'h3)];
              reg831 <= (!$unsigned(reg830[(2'h2):(2'h2)]));
              reg832 = (($unsigned({((8'ha3) <<< reg800),
                          reg830[(3'h6):(3'h5)]}) ?
                      $signed($signed((reg701 == reg740))) : $signed((!wire776))) ?
                  {((((8'hbf) ? reg685 : reg763) >>> reg813) ?
                          $signed({reg762, reg785}) : (reg733 == {wire679,
                              reg740})),
                      reg830} : $unsigned($unsigned($unsigned($unsigned(reg785)))));
              reg833 <= ((reg683 & wire682) ?
                  (-(reg752[(2'h2):(1'h0)] ?
                      $unsigned(((8'hbd) <= reg820)) : ((^reg808) || ((8'hb9) ^~ reg757)))) : (~|((8'hbf) ?
                      {$unsigned(reg731)} : (8'hb3))));
            end
          else
            begin
              reg829 = $unsigned(reg716[(1'h0):(1'h0)]);
              reg830 = ($signed($unsigned(((wire680 ? (8'hb3) : reg731) ?
                      $unsigned(wire681) : (reg698 ? reg755 : reg781)))) ?
                  reg800[(4'h9):(3'h5)] : reg692[(1'h1):(1'h1)]);
              reg831 <= ($unsigned(($signed($unsigned(reg806)) - reg826)) ?
                  $signed($unsigned(reg755[(3'h4):(1'h0)])) : $unsigned($signed(((wire736 >= reg698) ^ (reg831 <<< reg761)))));
              reg833 <= ($signed((~|$unsigned((reg692 >>> reg742)))) + reg755);
            end
          if ({reg828[(4'h8):(4'h8)],
              $unsigned((((reg690 + (8'ha9)) ?
                  (reg755 ?
                      wire776 : reg828) : (^~reg716)) >> reg806[(1'h1):(1'h0)]))})
            begin
              reg834 = ((reg790[(4'h8):(2'h3)] ?
                      (^~$signed(reg768[(1'h0):(1'h0)])) : reg733[(1'h0):(1'h0)]) ?
                  reg820 : {(~&{$unsigned((8'hbd))}),
                      {{$signed(reg773), {(7'h43)}}}});
              reg835 <= reg829[(5'h15):(4'h8)];
              reg836 <= ($unsigned((reg698 || reg698[(1'h1):(1'h1)])) ?
                  reg703 : {reg692, reg810[(4'hb):(1'h0)]});
              reg837 = {$unsigned(reg705[(2'h3):(2'h3)])};
            end
          else
            begin
              reg834 = (|($signed(((reg791 * reg741) ?
                      $unsigned(reg808) : $unsigned(reg733))) ?
                  $unsigned($signed(reg763[(3'h6):(3'h5)])) : ({(reg728 ?
                          reg695 : reg705),
                      $signed(reg800)} ^~ reg740)));
              reg837 = ($signed($unsigned(((wire776 <<< reg753) >= $unsigned(reg728)))) ?
                  $unsigned($unsigned({(~^(7'h43))})) : (reg708[(3'h5):(1'h0)] << (($unsigned(reg695) || (reg703 || reg792)) ?
                      (reg707 - (8'haf)) : ((8'hae) ?
                          {(8'hb5), reg740} : (~reg836)))));
            end
          if ((~^(+(~|reg709))))
            begin
              reg838 <= (-(^~reg743));
            end
          else
            begin
              reg838 <= reg725;
              reg839 = ((^(!$unsigned((reg808 > reg791)))) ?
                  reg721[(2'h3):(1'h0)] : $unsigned(((~reg741[(3'h4):(1'h1)]) && $unsigned((+reg768)))));
              reg840 <= $unsigned(({{wire799,
                      (reg746 ? reg781 : (7'h41))}} && (&reg829)));
              reg841 = (reg832 ?
                  (reg709[(2'h2):(2'h2)] ?
                      (8'ha1) : $unsigned(reg692[(1'h1):(1'h0)])) : reg697[(3'h7):(3'h6)]);
            end
          for (forvar842 = (1'h0); (forvar842 < (2'h2)); forvar842 = (forvar842 + (1'h1)))
            begin
              reg843 = (((~|$unsigned(reg767)) ?
                  (!{$unsigned(reg750)}) : {((wire681 && reg721) || reg835[(4'h8):(1'h1)]),
                      $signed($unsigned(reg812))}) & wire799[(3'h6):(3'h4)]);
              reg844 = ($signed($signed(wire776)) ?
                  $unsigned(((~^{reg708}) ?
                      $unsigned((~reg746)) : {$unsigned(reg703)})) : reg835);
            end
          if (reg768[(1'h1):(1'h0)])
            begin
              reg845 = reg753;
            end
          else
            begin
              reg846 <= (((reg690[(3'h7):(3'h4)] ?
                  $signed((reg740 == reg833)) : (|(reg743 & reg820))) && {reg716[(1'h0):(1'h0)],
                  (reg733 ?
                      {reg735,
                          reg742} : reg750)}) && $unsigned($signed(({reg813} >> $signed(reg757)))));
              reg847 = $unsigned($signed(reg746));
            end
        end
      else
        begin
          for (forvar829 = (1'h0); (forvar829 < (3'h4)); forvar829 = (forvar829 + (1'h1)))
            begin
              reg830 = reg773;
              reg832 = (!({(&(reg843 ^ reg846)),
                  (!(reg764 ?
                      reg807 : reg683))} && $unsigned($signed(((7'h44) >> wire680)))));
              reg834 = $signed(((~|(reg735[(4'h8):(1'h1)] ?
                      $signed(reg753) : (~&wire776))) ?
                  (($unsigned(reg767) || reg753[(3'h6):(2'h2)]) ?
                      (~wire679[(3'h7):(3'h5)]) : reg728) : reg716[(1'h0):(1'h0)]));
              reg835 <= $unsigned((^{((!forvar842) ~^ {reg835}), (7'h48)}));
              reg836 <= reg838[(1'h0):(1'h0)];
            end
        end
      if ((^((wire736[(4'h8):(2'h2)] ?
          reg750[(3'h4):(1'h0)] : reg790) || $signed({$unsigned(reg800)}))))
        begin
          reg848 <= ({reg836} & reg708);
        end
      else
        begin
          if (reg831)
            begin
              reg848 <= ($signed(((+$signed(reg690)) ?
                      $signed(reg844[(2'h3):(2'h2)]) : (~^$unsigned(wire776)))) ?
                  ((|reg718[(2'h2):(1'h0)]) < ($signed((reg773 || reg831)) >>> {(reg838 << forvar842),
                      reg735})) : $signed($signed(reg830[(3'h7):(3'h5)])));
              reg849 <= ((!((+$unsigned(reg755)) > (8'hb4))) ?
                  forvar829[(1'h1):(1'h1)] : (($unsigned((reg844 ?
                              reg848 : reg697)) ?
                          reg698 : $unsigned($unsigned(reg735))) ?
                      $signed(wire681[(4'hb):(3'h6)]) : reg843));
              reg850 = reg699[(1'h1):(1'h1)];
            end
          else
            begin
              reg848 <= (((($unsigned(reg683) >> (reg848 ~^ reg733)) | (8'hb8)) << (reg826[(5'h11):(3'h5)] ?
                      reg821 : (~&$signed(wire681)))) ?
                  ((reg709[(1'h1):(1'h1)] * reg709[(1'h1):(1'h0)]) == (8'hb7)) : reg686[(1'h0):(1'h0)]);
              reg849 <= reg829;
              reg851 <= ($signed(reg740[(3'h7):(3'h5)]) >= (~|(^$signed((^reg786)))));
            end
          for (forvar852 = (1'h0); (forvar852 < (1'h0)); forvar852 = (forvar852 + (1'h1)))
            begin
              reg853 = (!$signed(reg716[(3'h4):(1'h1)]));
            end
          reg854 = $signed(reg808[(3'h4):(3'h4)]);
          reg855 = $signed((~|(($unsigned(reg707) ?
                  $signed((8'h9c)) : $signed(reg786)) ?
              (^reg767[(1'h0):(1'h0)]) : ((^~reg743) ?
                  (wire736 || reg768) : $signed((7'h45))))));
          if (reg692[(3'h4):(2'h2)])
            begin
              reg856 = (reg840 <<< {$signed((~$signed(reg844))),
                  $unsigned(wire680)});
              reg857 = (^$unsigned(reg851[(4'h9):(2'h3)]));
              reg858 = reg800;
            end
          else
            begin
              reg856 = {reg826[(1'h1):(1'h1)],
                  ({(reg741 ? $signed((8'ha1)) : (reg825 < reg764)),
                      (reg838 ?
                          (+reg742) : (&reg831))} >>> $signed($signed((reg683 ?
                      reg705 : reg718))))};
              reg857 = reg767[(4'hc):(1'h0)];
              reg858 = (reg849 >= (~|reg707[(4'h9):(3'h6)]));
              reg859 <= (^~reg761[(2'h2):(1'h0)]);
              reg860 <= reg757;
            end
        end
      for (forvar861 = (1'h0); (forvar861 < (1'h1)); forvar861 = (forvar861 + (1'h1)))
        begin
          reg862 = reg701[(5'h11):(3'h4)];
          for (forvar863 = (1'h0); (forvar863 < (2'h3)); forvar863 = (forvar863 + (1'h1)))
            begin
              reg864 <= {{reg742},
                  $unsigned(({reg837} <<< $unsigned((~&reg831))))};
              reg865 = reg753[(3'h7):(3'h7)];
              reg866 <= {$signed((!(reg762[(4'ha):(3'h6)] ?
                      {reg835, reg718} : $unsigned(reg837))))};
              reg867 <= reg840[(3'h5):(2'h2)];
              reg868 = ($unsigned(({{forvar842}} ?
                      ((reg772 ? reg746 : reg827) ?
                          {(8'ha1)} : (^~reg864)) : ((8'h9e) ?
                          $signed((8'h9c)) : {(8'ha3), (8'hac)}))) ?
                  reg740 : $signed(((!$signed(reg847)) ?
                      reg866[(4'hf):(3'h4)] : $unsigned($unsigned(reg761)))));
            end
          if (forvar861)
            begin
              reg869 <= (8'hb1);
            end
          else
            begin
              reg869 <= $signed({$unsigned(((~reg853) ?
                      (reg829 - reg851) : reg829[(1'h0):(1'h0)])),
                  (wire680[(4'h9):(3'h7)] >= (reg857 - (reg762 == (8'h9e))))});
              reg870 = {{wire736, (8'ha4)},
                  $unsigned(((8'h9f) > $unsigned(((7'h46) ?
                      reg725 : reg746))))};
            end
          if (reg834)
            begin
              reg871 = reg741[(4'ha):(3'h4)];
              reg872 = (reg860 != reg768[(2'h3):(1'h0)]);
              reg873 = (reg791 ?
                  {(((reg687 ~^ reg743) <= reg703[(3'h5):(3'h4)]) | $unsigned(reg790))} : reg853);
              reg874 = reg708[(3'h4):(2'h2)];
              reg875 = $signed($signed((|(~^wire776[(3'h5):(1'h0)]))));
            end
          else
            begin
              reg871 = {reg709[(2'h2):(1'h0)]};
              reg872 = (!($unsigned(reg844[(4'hf):(2'h3)]) ?
                  {($signed(reg832) & (&reg858)),
                      ($unsigned(reg707) ^ (reg697 && reg836))} : {$signed((reg855 - (8'hb4)))}));
            end
        end
      reg876 <= reg868[(4'h8):(2'h3)];
    end
  always
    @(posedge clk) begin
      for (forvar877 = (1'h0); (forvar877 < (2'h3)); forvar877 = (forvar877 + (1'h1)))
        begin
          reg878 = (^$signed((((reg821 ? reg707 : reg806) ?
                  (reg703 << reg692) : reg698[(3'h6):(1'h0)]) ?
              $unsigned((reg752 ?
                  reg792 : reg849)) : $unsigned($unsigned(reg735)))));
          reg879 = $signed((~&reg833));
        end
      if (($signed($unsigned($unsigned(reg794[(3'h7):(3'h5)]))) ?
          (~^(+($signed(reg878) ?
              $unsigned(reg725) : reg768))) : (~|(reg716[(2'h3):(1'h0)] != $signed((8'had))))))
        begin
          reg880 = $signed(wire679);
        end
      else
        begin
          for (forvar880 = (1'h0); (forvar880 < (2'h2)); forvar880 = (forvar880 + (1'h1)))
            begin
              reg881 = ($signed(forvar877) ?
                  reg743[(1'h1):(1'h1)] : {($unsigned($unsigned(reg794)) ?
                          reg683 : reg767),
                      {{((8'hbe) ? reg864 : reg741), $unsigned(reg859)},
                          reg848[(4'hb):(4'h9)]}});
              reg882 <= $signed((~&(reg752[(1'h0):(1'h0)] ?
                  {reg828[(1'h0):(1'h0)], $signed((8'haa))} : (&reg735))));
              reg883 <= $signed({$signed(reg757[(2'h3):(1'h1)]),
                  $unsigned(reg703)});
              reg884 <= (reg859[(2'h2):(1'h1)] ?
                  $unsigned($unsigned(reg836)) : reg687[(1'h1):(1'h0)]);
              reg885 = ((~&$unsigned(reg835[(4'hb):(4'ha)])) ?
                  reg882 : (reg750[(1'h0):(1'h0)] >= $signed($signed($unsigned((7'h43))))));
            end
          for (forvar886 = (1'h0); (forvar886 < (2'h3)); forvar886 = (forvar886 + (1'h1)))
            begin
              reg887 <= $signed((~&(-((reg786 ?
                  reg826 : reg791) >= (reg848 <<< reg752)))));
              reg888 = ($signed((reg876 * $unsigned(((8'ha1) ?
                      reg806 : reg733)))) ?
                  $signed(wire678) : ($signed($unsigned((!reg725))) ?
                      (reg882[(4'h8):(1'h0)] >>> {$unsigned(forvar877)}) : wire719));
            end
          for (forvar889 = (1'h0); (forvar889 < (2'h3)); forvar889 = (forvar889 + (1'h1)))
            begin
              reg890 <= $signed(reg825);
            end
          if ((~^$signed(reg884[(3'h6):(3'h4)])))
            begin
              reg891 <= $unsigned({(reg733[(1'h0):(1'h0)] ?
                      reg821 : (|(!(8'ha2))))});
              reg892 = reg716;
              reg893 = reg838;
              reg894 <= $signed(reg741);
              reg895 = (^~reg859[(4'h8):(3'h7)]);
            end
          else
            begin
              reg891 <= ((^~(((reg755 ? reg707 : reg750) << $unsigned(reg794)) ?
                  reg755[(4'h8):(1'h0)] : reg731[(3'h7):(2'h2)])) >>> reg820);
              reg894 <= reg762[(4'he):(3'h4)];
              reg895 = reg750;
              reg896 <= {reg821};
            end
        end
      for (forvar897 = (1'h0); (forvar897 < (2'h3)); forvar897 = (forvar897 + (1'h1)))
        begin
          reg898 <= ((~^reg887[(1'h1):(1'h0)]) <= {(8'hb6)});
        end
      for (forvar899 = (1'h0); (forvar899 < (1'h0)); forvar899 = (forvar899 + (1'h1)))
        begin
          reg900 = (reg741 ~^ (+((|{reg701, reg794}) ? reg892 : (~^(8'hb3)))));
          reg901 <= $unsigned((^~reg747));
          reg902 <= (^~(($unsigned($signed(reg750)) <= (^~reg900)) ?
              reg864 : (+{reg709})));
        end
      for (forvar903 = (1'h0); (forvar903 < (2'h3)); forvar903 = (forvar903 + (1'h1)))
        begin
          reg904 = wire799[(4'h8):(1'h0)];
          reg905 <= $signed($unsigned(wire682));
        end
    end
  always
    @(posedge clk) begin
      reg906 = reg786;
    end
  always
    @(posedge clk) begin
      reg907 <= reg755[(4'h8):(3'h5)];
      reg908 = reg883;
      reg909 <= (^{reg813, reg698[(1'h1):(1'h1)]});
    end
  always
    @(posedge clk) begin
      reg910 <= ((reg909[(3'h4):(3'h4)] ? reg695[(2'h2):(1'h0)] : wire776) ?
          {$unsigned(reg883)} : reg768);
      reg911 = $signed((&$unsigned(reg686)));
      reg912 <= (wire799 ?
          ({(8'hbf), reg859} + ((reg911 >= reg833[(4'h9):(4'h8)]) ?
              ($signed(wire776) ~^ {reg687, reg767}) : ((reg747 ?
                  wire680 : reg820) + (~|reg898)))) : reg746[(1'h0):(1'h0)]);
      reg913 <= reg848[(4'h9):(1'h0)];
      reg914 = $signed($signed({(&((7'h45) * reg753)), reg905}));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module385
#(parameter param654 = ((-((8'hbe) > (&((8'h9c) ? (8'hb3) : (8'ha6))))) ? {(((^(7'h49)) * (^~(8'h9e))) ? (&((8'ha6) ? (8'ha6) : (7'h48))) : ({(8'ha5), (8'haf)} ? ((8'ha5) ^ (7'h40)) : ((8'hac) && (8'ha1)))), {(((8'h9c) << (8'h9c)) ? (~|(8'hbf)) : ((8'haf) ? (8'ha5) : (8'ha6))), (~^(+(8'ha4)))}} : (({((8'haf) ? (8'h9c) : (8'h9d)), (~(8'hbd))} ? (^((7'h43) ? (7'h45) : (8'hb5))) : (((8'hb8) <<< (8'ha7)) ? (8'ha1) : (~(8'h9d)))) ? ((^((8'hb5) << (7'h44))) ? {((8'h9e) >= (8'ha7))} : (&((8'hb5) ? (7'h49) : (8'hb6)))) : ({((7'h44) ? (8'hb6) : (7'h41)), ((7'h46) ? (8'hbc) : (8'hb4))} ? ({(8'hbd), (8'ha6)} ^ (+(8'hbb))) : (((8'hb0) ? (8'hbb) : (8'hb4)) ? (+(8'h9d)) : (^(8'ha1)))))), 
parameter param655 = ((|{(^~{(7'h45), param654}), param654}) < (!(8'hae))))
(y, clk, wire389, wire388, wire387, wire386);
  output wire [(32'hd28):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire389;
  input wire [(5'h15):(1'h0)] wire388;
  input wire [(5'h12):(1'h0)] wire387;
  input wire signed [(4'h8):(1'h0)] wire386;
  wire [(5'h12):(1'h0)] wire587;
  wire signed [(5'h13):(1'h0)] wire562;
  wire [(5'h11):(1'h0)] wire561;
  wire [(3'h6):(1'h0)] wire545;
  wire signed [(5'h10):(1'h0)] wire544;
  wire [(4'hd):(1'h0)] wire516;
  wire signed [(4'ha):(1'h0)] wire515;
  wire [(5'h11):(1'h0)] wire514;
  wire signed [(5'h17):(1'h0)] wire470;
  wire signed [(2'h2):(1'h0)] wire400;
  wire [(2'h2):(1'h0)] wire399;
  reg [(3'h6):(1'h0)] reg650 = (1'h0);
  reg [(5'h17):(1'h0)] reg648 = (1'h0);
  reg [(4'hf):(1'h0)] reg644 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg643 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg642 = (1'h0);
  reg [(4'hd):(1'h0)] reg641 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg640 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg637 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg633 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg632 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg631 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg629 = (1'h0);
  reg [(5'h12):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg627 = (1'h0);
  reg [(3'h7):(1'h0)] reg626 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg625 = (1'h0);
  reg [(2'h2):(1'h0)] reg623 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg622 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg621 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg616 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg615 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg614 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg611 = (1'h0);
  reg [(3'h6):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg606 = (1'h0);
  reg [(4'hd):(1'h0)] reg605 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg602 = (1'h0);
  reg [(4'hc):(1'h0)] reg601 = (1'h0);
  reg [(4'h9):(1'h0)] reg594 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg598 = (1'h0);
  reg [(5'h11):(1'h0)] reg597 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg591 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg590 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg589 = (1'h0);
  reg [(5'h11):(1'h0)] reg584 = (1'h0);
  reg [(4'h8):(1'h0)] reg583 = (1'h0);
  reg [(5'h11):(1'h0)] reg580 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg575 = (1'h0);
  reg [(3'h7):(1'h0)] reg574 = (1'h0);
  reg [(5'h14):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg571 = (1'h0);
  reg [(5'h11):(1'h0)] reg567 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg565 = (1'h0);
  reg [(5'h17):(1'h0)] reg564 = (1'h0);
  reg [(3'h6):(1'h0)] reg563 = (1'h0);
  reg signed [(4'he):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg557 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg556 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg554 = (1'h0);
  reg [(4'h8):(1'h0)] reg551 = (1'h0);
  reg [(2'h3):(1'h0)] reg550 = (1'h0);
  reg [(4'he):(1'h0)] reg539 = (1'h0);
  reg [(5'h12):(1'h0)] reg538 = (1'h0);
  reg [(4'hf):(1'h0)] reg535 = (1'h0);
  reg [(5'h15):(1'h0)] reg529 = (1'h0);
  reg signed [(4'he):(1'h0)] reg527 = (1'h0);
  reg [(3'h7):(1'h0)] reg526 = (1'h0);
  reg [(5'h17):(1'h0)] reg525 = (1'h0);
  reg [(4'hb):(1'h0)] reg524 = (1'h0);
  reg [(5'h12):(1'h0)] reg523 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg520 = (1'h0);
  reg [(5'h16):(1'h0)] reg519 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg518 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg513 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg511 = (1'h0);
  reg [(5'h13):(1'h0)] reg509 = (1'h0);
  reg [(4'hf):(1'h0)] reg508 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg507 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg505 = (1'h0);
  reg [(4'h8):(1'h0)] reg504 = (1'h0);
  reg [(3'h6):(1'h0)] reg503 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg498 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg495 = (1'h0);
  reg [(5'h16):(1'h0)] reg494 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg489 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg486 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg485 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg483 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg481 = (1'h0);
  reg [(3'h6):(1'h0)] reg480 = (1'h0);
  reg [(4'hd):(1'h0)] reg479 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg478 = (1'h0);
  reg [(4'hc):(1'h0)] reg476 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg472 = (1'h0);
  reg [(5'h17):(1'h0)] reg471 = (1'h0);
  reg signed [(4'he):(1'h0)] reg467 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg466 = (1'h0);
  reg [(2'h3):(1'h0)] reg465 = (1'h0);
  reg [(2'h2):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg458 = (1'h0);
  reg [(3'h6):(1'h0)] reg457 = (1'h0);
  reg [(2'h2):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg451 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg449 = (1'h0);
  reg [(5'h10):(1'h0)] reg448 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg447 = (1'h0);
  reg [(4'hd):(1'h0)] reg446 = (1'h0);
  reg [(5'h13):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg441 = (1'h0);
  reg [(4'hb):(1'h0)] reg437 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg435 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg430 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg428 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg427 = (1'h0);
  reg [(4'he):(1'h0)] reg424 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg422 = (1'h0);
  reg [(4'he):(1'h0)] reg419 = (1'h0);
  reg [(3'h7):(1'h0)] reg417 = (1'h0);
  reg [(4'hc):(1'h0)] reg416 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg415 = (1'h0);
  reg [(4'hc):(1'h0)] reg413 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg412 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg410 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg408 = (1'h0);
  reg [(3'h7):(1'h0)] reg407 = (1'h0);
  reg [(5'h13):(1'h0)] reg404 = (1'h0);
  reg [(4'h8):(1'h0)] reg403 = (1'h0);
  reg [(5'h18):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg398 = (1'h0);
  reg [(2'h2):(1'h0)] reg397 = (1'h0);
  reg [(4'hd):(1'h0)] reg396 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg393 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg391 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg390 = (1'h0);
  reg [(3'h4):(1'h0)] reg653 = (1'h0);
  reg [(5'h12):(1'h0)] forvar652 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar649 = (1'h0);
  reg [(3'h4):(1'h0)] reg647 = (1'h0);
  reg [(5'h10):(1'h0)] reg646 = (1'h0);
  reg [(2'h2):(1'h0)] reg645 = (1'h0);
  reg [(4'hd):(1'h0)] reg639 = (1'h0);
  reg [(5'h13):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar636 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar635 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg634 = (1'h0);
  reg [(5'h12):(1'h0)] reg630 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar620 = (1'h0);
  reg [(4'hc):(1'h0)] reg619 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg618 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg617 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg613 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg612 = (1'h0);
  reg [(5'h16):(1'h0)] reg610 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar609 = (1'h0);
  reg [(2'h2):(1'h0)] reg607 = (1'h0);
  reg [(3'h5):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg603 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg600 = (1'h0);
  reg [(5'h14):(1'h0)] reg599 = (1'h0);
  reg [(3'h4):(1'h0)] forvar588 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg596 = (1'h0);
  reg [(4'hb):(1'h0)] reg595 = (1'h0);
  reg [(3'h4):(1'h0)] forvar594 = (1'h0);
  reg [(5'h13):(1'h0)] reg593 = (1'h0);
  reg [(5'h10):(1'h0)] reg592 = (1'h0);
  reg [(2'h3):(1'h0)] reg588 = (1'h0);
  reg [(5'h17):(1'h0)] reg586 = (1'h0);
  reg [(5'h16):(1'h0)] reg585 = (1'h0);
  reg [(5'h11):(1'h0)] reg582 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg581 = (1'h0);
  reg [(2'h3):(1'h0)] forvar579 = (1'h0);
  reg [(4'h8):(1'h0)] reg578 = (1'h0);
  reg [(5'h17):(1'h0)] reg577 = (1'h0);
  reg [(4'h9):(1'h0)] reg576 = (1'h0);
  reg [(5'h15):(1'h0)] reg572 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg569 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg568 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg566 = (1'h0);
  reg signed [(4'he):(1'h0)] reg560 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar558 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg555 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar551 = (1'h0);
  reg [(5'h15):(1'h0)] reg553 = (1'h0);
  reg [(4'h8):(1'h0)] reg552 = (1'h0);
  reg [(4'hf):(1'h0)] reg549 = (1'h0);
  reg [(3'h6):(1'h0)] reg548 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg547 = (1'h0);
  reg [(4'h9):(1'h0)] reg546 = (1'h0);
  reg [(2'h3):(1'h0)] reg543 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg542 = (1'h0);
  reg [(4'h9):(1'h0)] reg541 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg540 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar537 = (1'h0);
  reg [(4'hc):(1'h0)] reg536 = (1'h0);
  reg [(5'h11):(1'h0)] reg534 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg533 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar532 = (1'h0);
  reg [(5'h15):(1'h0)] forvar531 = (1'h0);
  reg [(2'h3):(1'h0)] reg530 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg522 = (1'h0);
  reg [(5'h17):(1'h0)] forvar521 = (1'h0);
  reg [(3'h5):(1'h0)] forvar517 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg512 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg510 = (1'h0);
  reg [(4'hd):(1'h0)] reg506 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg502 = (1'h0);
  reg [(5'h18):(1'h0)] reg501 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg500 = (1'h0);
  reg [(5'h13):(1'h0)] reg499 = (1'h0);
  reg [(5'h15):(1'h0)] forvar497 = (1'h0);
  reg [(3'h6):(1'h0)] reg496 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg493 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg492 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg490 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg488 = (1'h0);
  reg [(4'h8):(1'h0)] reg487 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg484 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg477 = (1'h0);
  reg [(3'h4):(1'h0)] reg475 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg474 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar473 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg455 = (1'h0);
  reg [(5'h17):(1'h0)] reg469 = (1'h0);
  reg [(3'h6):(1'h0)] reg468 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg464 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar463 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg462 = (1'h0);
  reg [(4'he):(1'h0)] reg460 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar455 = (1'h0);
  reg [(4'h9):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg452 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg450 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg444 = (1'h0);
  reg [(5'h13):(1'h0)] reg445 = (1'h0);
  reg [(4'hd):(1'h0)] forvar444 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg443 = (1'h0);
  reg [(5'h10):(1'h0)] reg440 = (1'h0);
  reg [(5'h15):(1'h0)] reg439 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg438 = (1'h0);
  reg [(5'h10):(1'h0)] forvar436 = (1'h0);
  reg [(4'hc):(1'h0)] reg434 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg433 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar432 = (1'h0);
  reg [(5'h17):(1'h0)] reg431 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg429 = (1'h0);
  reg [(4'hd):(1'h0)] forvar426 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg425 = (1'h0);
  reg signed [(4'he):(1'h0)] reg423 = (1'h0);
  reg [(3'h5):(1'h0)] forvar421 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg420 = (1'h0);
  reg signed [(4'he):(1'h0)] reg418 = (1'h0);
  reg [(3'h4):(1'h0)] forvar414 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg411 = (1'h0);
  reg [(5'h13):(1'h0)] reg409 = (1'h0);
  reg [(4'hf):(1'h0)] reg406 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg405 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar402 = (1'h0);
  reg [(4'ha):(1'h0)] reg395 = (1'h0);
  reg [(5'h11):(1'h0)] forvar394 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg392 = (1'h0);
  assign y = {wire587,
                 wire562,
                 wire561,
                 wire545,
                 wire544,
                 wire516,
                 wire515,
                 wire514,
                 wire470,
                 wire400,
                 wire399,
                 reg650,
                 reg648,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg640,
                 reg637,
                 reg633,
                 reg632,
                 reg631,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg625,
                 reg623,
                 reg622,
                 reg621,
                 reg616,
                 reg615,
                 reg614,
                 reg611,
                 reg608,
                 reg606,
                 reg605,
                 reg602,
                 reg601,
                 reg594,
                 reg598,
                 reg597,
                 reg591,
                 reg590,
                 reg589,
                 reg584,
                 reg583,
                 reg580,
                 reg575,
                 reg574,
                 reg573,
                 reg571,
                 reg567,
                 reg565,
                 reg564,
                 reg563,
                 reg559,
                 reg557,
                 reg556,
                 reg554,
                 reg551,
                 reg550,
                 reg539,
                 reg538,
                 reg535,
                 reg529,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg520,
                 reg519,
                 reg518,
                 reg513,
                 reg511,
                 reg509,
                 reg508,
                 reg507,
                 reg505,
                 reg504,
                 reg503,
                 reg498,
                 reg495,
                 reg494,
                 reg489,
                 reg486,
                 reg485,
                 reg483,
                 reg481,
                 reg480,
                 reg479,
                 reg478,
                 reg476,
                 reg472,
                 reg471,
                 reg467,
                 reg466,
                 reg465,
                 reg461,
                 reg458,
                 reg457,
                 reg453,
                 reg451,
                 reg449,
                 reg448,
                 reg447,
                 reg446,
                 reg442,
                 reg441,
                 reg437,
                 reg435,
                 reg430,
                 reg428,
                 reg427,
                 reg424,
                 reg422,
                 reg419,
                 reg417,
                 reg416,
                 reg415,
                 reg413,
                 reg412,
                 reg410,
                 reg408,
                 reg407,
                 reg404,
                 reg403,
                 reg401,
                 reg398,
                 reg397,
                 reg396,
                 reg393,
                 reg391,
                 reg390,
                 reg653,
                 forvar652,
                 reg651,
                 forvar649,
                 reg647,
                 reg646,
                 reg645,
                 reg639,
                 reg638,
                 forvar636,
                 forvar635,
                 reg634,
                 reg630,
                 reg624,
                 forvar620,
                 reg619,
                 reg618,
                 reg617,
                 reg613,
                 reg612,
                 reg610,
                 forvar609,
                 reg607,
                 reg604,
                 reg603,
                 reg600,
                 reg599,
                 forvar588,
                 reg596,
                 reg595,
                 forvar594,
                 reg593,
                 reg592,
                 reg588,
                 reg586,
                 reg585,
                 reg582,
                 reg581,
                 forvar579,
                 reg578,
                 reg577,
                 reg576,
                 reg572,
                 reg570,
                 reg569,
                 reg568,
                 reg566,
                 reg560,
                 forvar558,
                 reg555,
                 forvar551,
                 reg553,
                 reg552,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 reg543,
                 reg542,
                 reg541,
                 reg540,
                 forvar537,
                 reg536,
                 reg534,
                 reg533,
                 forvar532,
                 forvar531,
                 reg530,
                 reg528,
                 reg522,
                 forvar521,
                 forvar517,
                 reg512,
                 reg510,
                 reg506,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 forvar497,
                 reg496,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 reg488,
                 reg487,
                 reg484,
                 reg482,
                 reg477,
                 reg475,
                 reg474,
                 forvar473,
                 reg455,
                 reg469,
                 reg468,
                 reg464,
                 forvar463,
                 reg462,
                 reg460,
                 reg459,
                 reg456,
                 forvar455,
                 reg454,
                 reg452,
                 reg450,
                 reg444,
                 reg445,
                 forvar444,
                 reg443,
                 reg440,
                 reg439,
                 reg438,
                 forvar436,
                 reg434,
                 reg433,
                 forvar432,
                 reg431,
                 reg429,
                 forvar426,
                 reg425,
                 reg423,
                 forvar421,
                 reg420,
                 reg418,
                 forvar414,
                 reg411,
                 reg409,
                 reg406,
                 reg405,
                 forvar402,
                 reg395,
                 forvar394,
                 reg392,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire389[(5'h12):(5'h12)])
        begin
          reg390 <= $unsigned((~^wire389));
          reg391 <= ($signed($unsigned((-(-wire389)))) ?
              (^~$signed(((reg390 ?
                  wire386 : wire388) ^~ wire386))) : $unsigned(((&$unsigned(wire386)) << (wire388 && (wire386 ?
                  (8'hb6) : wire386)))));
        end
      else
        begin
          if (reg390)
            begin
              reg392 = (((reg390 ?
                      $signed(wire387[(4'he):(3'h4)]) : (~$signed(wire387))) ?
                  $signed($unsigned(wire386[(3'h7):(3'h7)])) : $signed(wire389[(1'h1):(1'h1)])) & $unsigned(wire386));
            end
          else
            begin
              reg392 = wire388;
            end
          reg393 <= wire387;
          for (forvar394 = (1'h0); (forvar394 < (3'h4)); forvar394 = (forvar394 + (1'h1)))
            begin
              reg395 = $unsigned((((wire386[(3'h5):(3'h5)] ?
                      $signed(wire389) : $unsigned(wire388)) * reg391) ?
                  ($unsigned(wire388[(5'h11):(4'hf)]) ~^ $unsigned((~&reg393))) : $signed(wire389[(4'h8):(3'h7)])));
              reg396 <= (wire388[(3'h7):(3'h4)] >>> $unsigned(($signed((reg392 ?
                  (7'h42) : (8'ha5))) | $unsigned(wire388[(4'h9):(3'h7)]))));
              reg397 <= reg390;
            end
          reg398 <= (~$unsigned(((!(&reg393)) * (-$signed(wire389)))));
        end
    end
  assign wire399 = $unsigned(($signed(reg390[(1'h1):(1'h1)]) ?
                       (~^(!wire388[(5'h13):(2'h3)])) : $signed(reg398[(4'hf):(3'h7)])));
  assign wire400 = ((~{((reg396 << wire386) - reg390[(2'h2):(2'h2)]),
                           $signed(reg396)}) ?
                       ($signed({((7'h48) | wire387)}) ?
                           (&{$signed(wire399),
                               $signed(reg398)}) : (8'hb4)) : (wire387 ?
                           (~($signed(reg397) ?
                               ((8'hbb) ? reg397 : reg393) : (reg391 ?
                                   reg393 : reg390))) : (!$signed((wire388 > reg390)))));
  always
    @(posedge clk) begin
      reg401 <= {(($unsigned((~&reg396)) ?
              (&$signed((8'ha1))) : $signed((wire388 ?
                  (8'hbe) : reg391))) <<< wire386[(4'h8):(1'h0)]),
          ({(^~(reg391 ~^ reg390)), reg397} ? {(7'h43)} : (8'hbe))};
      for (forvar402 = (1'h0); (forvar402 < (1'h1)); forvar402 = (forvar402 + (1'h1)))
        begin
          reg403 <= ((~^$unsigned((7'h49))) & $unsigned(($signed((reg401 ?
                  reg398 : (7'h40))) ?
              (^reg396[(4'ha):(3'h5)]) : wire387)));
          if (({reg403, $signed(($unsigned(reg396) ^ wire399[(1'h0):(1'h0)]))} ?
              $unsigned((((reg390 ? wire389 : wire389) ?
                  forvar402 : (!wire389)) >> reg397[(1'h1):(1'h1)])) : reg397[(2'h2):(1'h0)]))
            begin
              reg404 <= wire386;
              reg405 = $signed((~|(~^(&(!reg396)))));
              reg406 = (+reg397);
              reg407 <= wire399;
            end
          else
            begin
              reg405 = reg403[(1'h1):(1'h1)];
              reg407 <= ($unsigned(wire386) >= ((-(forvar402 ?
                  $unsigned(reg401) : (!reg397))) ^ ($signed(forvar402[(3'h6):(2'h3)]) ?
                  reg406[(4'h9):(2'h2)] : reg391)));
            end
        end
      reg408 <= (reg396 * $signed(reg393));
    end
  always
    @(posedge clk) begin
      if ((^wire399))
        begin
          reg409 = (((~{(~|reg407)}) ?
              ($unsigned($unsigned(reg398)) ?
                  reg407 : {$unsigned(wire386),
                      (~^reg396)}) : $unsigned((8'ha0))) ~^ {wire389[(5'h14):(5'h14)],
              ({$signed(reg407), (^~(8'hbe))} ?
                  (wire386 ^ (8'h9e)) : reg407[(2'h3):(2'h3)])});
        end
      else
        begin
          if (((-({(7'h48), (reg397 >>> reg401)} ?
                  $unsigned(wire388) : (~|(wire389 ? reg397 : wire389)))) ?
              {$signed((~|reg391)),
                  {(^~(!reg397)),
                      reg409[(4'he):(4'he)]}} : reg397[(1'h0):(1'h0)]))
            begin
              reg409 = wire386[(1'h1):(1'h1)];
              reg410 <= ({($signed((!reg408)) << ($signed(wire386) != $signed(reg391)))} ?
                  ((reg398 ?
                      $signed((~wire387)) : (((8'ha7) ?
                          reg390 : reg404) <<< (reg398 ?
                          wire389 : reg393))) > $unsigned((8'h9f))) : reg391[(4'ha):(1'h1)]);
              reg411 = (7'h47);
              reg412 <= reg411;
            end
          else
            begin
              reg410 <= (reg397 >= reg393);
              reg412 <= $signed(wire387);
              reg413 <= ($unsigned((&($signed(wire399) + (reg403 ?
                  (7'h40) : wire389)))) >>> $signed({$unsigned((reg408 ?
                      reg412 : reg412))}));
            end
          for (forvar414 = (1'h0); (forvar414 < (1'h0)); forvar414 = (forvar414 + (1'h1)))
            begin
              reg415 <= $signed(((+((8'h9d) ? $signed((8'hb7)) : {reg390})) ?
                  (reg391[(2'h2):(2'h2)] ^~ reg408) : ($unsigned((~&wire399)) >> $unsigned((wire399 ?
                      reg390 : forvar414)))));
            end
          if (reg415[(1'h1):(1'h1)])
            begin
              reg416 <= wire386;
              reg417 <= {wire387[(4'he):(1'h0)]};
            end
          else
            begin
              reg416 <= (reg410 ?
                  ({(reg413[(4'h8):(3'h6)] ?
                          (reg411 * reg416) : $unsigned(reg416)),
                      (wire388[(1'h1):(1'h0)] ?
                          (!(8'hae)) : (|reg398))} > {($signed((8'h9c)) ^ (reg410 ?
                          reg404 : reg417))}) : reg407);
              reg418 = (($signed(reg396) | (&(reg396 * reg404[(5'h10):(3'h6)]))) ^ wire389);
              reg419 <= reg413[(2'h2):(2'h2)];
              reg420 = reg419;
            end
          for (forvar421 = (1'h0); (forvar421 < (1'h0)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg422 <= (wire389 ?
                  reg393[(2'h3):(2'h3)] : ((|$unsigned(reg420)) ?
                      (|{(reg418 <= reg396),
                          $signed((8'h9f))}) : reg408[(2'h3):(2'h3)]));
              reg423 = (8'h9d);
              reg424 <= ((wire388[(5'h14):(2'h2)] != reg410[(4'ha):(4'ha)]) ?
                  (reg397[(2'h2):(1'h1)] ?
                      {((forvar414 ? reg397 : reg419) ?
                              reg412 : $signed(reg396))} : $signed(wire387[(4'he):(4'ha)])) : $signed($signed(((~reg411) ~^ (^(8'hba))))));
              reg425 = $signed((reg420 + $unsigned((!(reg418 << reg420)))));
            end
          for (forvar426 = (1'h0); (forvar426 < (1'h1)); forvar426 = (forvar426 + (1'h1)))
            begin
              reg427 <= $signed($signed(reg397));
              reg428 <= $unsigned(reg417[(3'h7):(3'h6)]);
              reg429 = $signed({(wire399 ?
                      (((8'haa) ~^ wire389) << (reg413 && (8'ha7))) : $signed(reg393[(1'h1):(1'h0)])),
                  (-$unsigned((reg411 ? (8'haf) : reg410)))});
              reg430 <= {(reg416 & reg415[(3'h4):(2'h3)]),
                  $unsigned($signed((~|(reg420 || reg396))))};
              reg431 = $signed(({(((8'hba) ? wire400 : reg410) ?
                          ((8'hba) ? reg409 : reg403) : ((7'h45) ^ reg417))} ?
                  reg403[(1'h0):(1'h0)] : (($unsigned(reg429) ?
                      reg416 : reg398[(4'hb):(3'h6)]) | $unsigned($unsigned((8'hbf))))));
            end
        end
      for (forvar432 = (1'h0); (forvar432 < (1'h0)); forvar432 = (forvar432 + (1'h1)))
        begin
          reg433 = {$unsigned((($signed(reg401) >= reg418) | $unsigned($unsigned(reg430))))};
          reg434 = (&reg408[(1'h0):(1'h0)]);
          reg435 <= wire387;
          for (forvar436 = (1'h0); (forvar436 < (3'h4)); forvar436 = (forvar436 + (1'h1)))
            begin
              reg437 <= (-reg396[(4'ha):(1'h0)]);
              reg438 = {(!reg419)};
              reg439 = $unsigned(($unsigned(((reg438 ? reg438 : (8'ha8)) ?
                      $unsigned(reg416) : reg408)) ?
                  ((7'h40) ?
                      $signed(((8'hbc) ?
                          reg409 : reg427)) : reg420) : $unsigned(({forvar432} ?
                      (7'h44) : forvar426))));
            end
          if (($signed(reg428[(5'h10):(5'h10)]) < $unsigned(reg398)))
            begin
              reg440 = forvar414[(3'h4):(2'h2)];
            end
          else
            begin
              reg441 <= $signed(reg434);
              reg442 <= (^forvar421[(3'h4):(2'h2)]);
            end
        end
      reg443 = $signed({$unsigned($signed($unsigned(reg442)))});
      if (((+(reg434 ? reg441[(5'h16):(3'h6)] : reg434)) ?
          (((~^$signed(wire388)) < ((^~reg418) >= wire388)) != reg403[(3'h4):(2'h2)]) : ($unsigned((reg403[(4'h8):(3'h4)] < forvar421[(2'h2):(1'h0)])) ?
              (&reg390[(1'h0):(1'h0)]) : ((reg403 | (&reg403)) <<< (~^$unsigned(reg440))))))
        begin
          for (forvar444 = (1'h0); (forvar444 < (2'h2)); forvar444 = (forvar444 + (1'h1)))
            begin
              reg445 = (reg407[(1'h1):(1'h0)] ?
                  (&reg390) : (forvar444[(1'h1):(1'h1)] ?
                      ((reg430[(2'h2):(2'h2)] ^~ (forvar436 ?
                              reg428 : reg434)) ?
                          (reg440[(4'h8):(3'h7)] ?
                              forvar414 : reg419[(2'h2):(2'h2)]) : $signed($unsigned(reg434))) : (reg440 && reg417[(2'h2):(1'h0)])));
            end
          reg446 <= (($unsigned($signed((&reg442))) * $unsigned($signed($signed(reg412)))) != reg390);
          reg447 <= (reg435 << $signed(wire388[(3'h7):(2'h2)]));
          reg448 <= reg428;
          reg449 <= ($signed(reg393[(3'h4):(3'h4)]) ?
              {forvar432[(5'h13):(4'h9)]} : ((|(reg397 >= reg401)) ?
                  (-$signed(wire388[(3'h5):(3'h5)])) : $unsigned($signed(reg420))));
        end
      else
        begin
          reg444 = (-reg440);
          if (($signed((~$unsigned((~|reg447)))) >= $signed({((+forvar421) ?
                  (reg437 >>> reg404) : $signed(reg403)),
              (7'h43)})))
            begin
              reg445 = reg409;
              reg446 <= wire386;
              reg450 = (($signed(reg425) ^~ (reg446[(3'h6):(2'h2)] != ($signed(reg417) == $unsigned(reg397)))) ?
                  (reg430 ?
                      (reg403 ?
                          $unsigned(reg430[(3'h6):(2'h3)]) : ((reg416 ?
                                  wire386 : reg446) ?
                              {forvar444,
                                  reg433} : $unsigned((8'ha9)))) : reg415[(2'h2):(1'h0)]) : ((+($unsigned(forvar414) + (reg423 >= wire400))) >>> reg393));
              reg451 <= reg396[(4'hc):(4'hb)];
              reg452 = $unsigned($unsigned(reg450[(3'h6):(3'h4)]));
            end
          else
            begin
              reg445 = ((reg411[(5'h14):(5'h11)] ?
                      (~&$signed($unsigned((8'hb1)))) : $signed((reg424[(3'h4):(2'h3)] || (reg427 ?
                          reg448 : reg413)))) ?
                  ($signed((-reg401)) == $unsigned($unsigned($unsigned((8'hab))))) : reg428);
              reg446 <= (8'hbd);
            end
          reg453 <= $signed($unsigned($unsigned(((reg439 >> reg434) ~^ ((7'h41) == reg452)))));
          reg454 = $unsigned($unsigned((reg428 ?
              ((~&reg431) == $unsigned(wire386)) : $unsigned(reg438[(2'h3):(2'h3)]))));
        end
      if ((($unsigned((reg442 & $signed(reg431))) <= (($signed(reg451) <= (reg452 != forvar426)) ?
          (|(^~forvar436)) : (~{reg430}))) * ($signed($signed((~reg437))) ?
          reg437[(4'h8):(1'h1)] : (($signed(wire387) || (reg437 ?
              reg413 : reg416)) && $unsigned(reg403[(4'h8):(2'h3)])))))
        begin
          for (forvar455 = (1'h0); (forvar455 < (1'h1)); forvar455 = (forvar455 + (1'h1)))
            begin
              reg456 = $unsigned($unsigned((~|wire399[(2'h2):(1'h0)])));
              reg457 <= {($unsigned(reg413) | {{(reg428 ? reg452 : reg451),
                          reg451[(3'h5):(2'h3)]}})};
            end
          reg458 <= ((^$signed(((8'ha6) || (~&reg404)))) ?
              {(^{$signed(reg446)})} : ((!reg427) ?
                  $unsigned(reg454[(2'h2):(1'h1)]) : (~|($signed(reg434) ?
                      forvar414 : {forvar444, reg409}))));
          if ({reg419, {reg454[(3'h6):(3'h4)], wire386}})
            begin
              reg459 = ({(((7'h45) * ((7'h46) + forvar444)) ?
                      reg427 : (+{reg411, reg411})),
                  $unsigned((reg396[(1'h1):(1'h0)] ?
                      reg456 : forvar421[(3'h5):(1'h0)]))} < reg443);
              reg460 = {($signed(reg409) > reg442)};
              reg461 <= (forvar436 ?
                  {{($unsigned(reg460) ? $unsigned(reg449) : forvar436)},
                      $signed(((reg446 << forvar421) ?
                          (reg457 ?
                              reg445 : (8'h9f)) : reg404[(4'ha):(4'h9)]))} : ((-((8'hbe) ?
                          reg419[(1'h1):(1'h0)] : (|reg447))) ?
                      (-({reg437, reg425} < {reg412,
                          reg438})) : $unsigned(reg448[(4'hf):(3'h6)])));
            end
          else
            begin
              reg459 = (8'ha9);
              reg461 <= (forvar414 ?
                  (wire387 - ((^(reg396 - reg411)) <<< {(reg444 ?
                          reg396 : reg437)})) : {reg430,
                      (((reg420 ? reg418 : reg428) & (^~(8'hb7))) ?
                          $unsigned({reg418}) : $signed(reg433))});
              reg462 = ({((^~(reg398 ? reg420 : reg445)) > ((forvar414 ?
                              reg401 : wire387) ?
                          (8'hac) : {forvar426, reg452})),
                      (((reg458 || (7'h43)) ?
                          reg444 : (!reg390)) << $signed(reg420[(4'h9):(3'h7)]))} ?
                  reg431 : reg390[(2'h2):(1'h1)]);
            end
          for (forvar463 = (1'h0); (forvar463 < (2'h3)); forvar463 = (forvar463 + (1'h1)))
            begin
              reg464 = reg454;
              reg465 <= (~|reg416[(3'h5):(2'h2)]);
              reg466 <= ($unsigned($unsigned(reg407)) ?
                  ((((~|reg401) ? reg460 : reg453) ?
                          (~&(wire399 <<< reg409)) : ((7'h40) ~^ $unsigned(reg412))) ?
                      ($unsigned($unsigned(reg415)) ?
                          ((reg398 && reg461) ?
                              {reg428,
                                  reg419} : $signed(reg445)) : ((~reg456) <= (reg460 || reg418))) : $signed($unsigned(reg461))) : reg397);
              reg467 <= ({(&reg411[(5'h17):(5'h10)])} ?
                  ((^($unsigned(reg403) ?
                      {reg419} : (forvar414 | reg450))) != wire387[(4'h8):(4'h8)]) : (((^((8'ha7) ?
                              wire400 : (7'h48))) ?
                          (reg453 >> (wire388 >>> reg424)) : reg408) ?
                      reg429 : forvar436));
              reg468 = reg435[(1'h1):(1'h0)];
            end
          reg469 = ((&$signed(reg415[(3'h6):(2'h3)])) > $unsigned({reg453[(1'h1):(1'h0)],
              $signed((reg409 ? reg451 : (8'h9d)))}));
        end
      else
        begin
          reg455 = $signed($signed(forvar455));
        end
    end
  assign wire470 = (($signed(reg448) ~^ $signed(({wire389,
                       reg458} ^~ $unsigned(reg457)))) ^~ {$signed({(8'h9f)}),
                       wire399});
  always
    @(posedge clk) begin
      reg471 <= reg417[(3'h7):(2'h2)];
      reg472 <= reg446[(1'h0):(1'h0)];
      if ($signed(($unsigned((^(wire387 + wire399))) ?
          $signed({reg391[(4'ha):(2'h2)],
              (!reg437)}) : $unsigned(reg407[(2'h3):(2'h3)]))))
        begin
          for (forvar473 = (1'h0); (forvar473 < (2'h3)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 = reg422;
              reg475 = ((reg453 ?
                  reg398[(3'h7):(3'h6)] : forvar473[(4'hc):(4'hc)]) * $signed($signed(reg466[(3'h4):(1'h1)])));
              reg476 <= wire386[(3'h7):(2'h3)];
            end
        end
      else
        begin
          for (forvar473 = (1'h0); (forvar473 < (2'h2)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg476 <= {(reg403 + $signed((reg417[(2'h2):(2'h2)] <= $unsigned(reg416)))),
                  (8'hb0)};
              reg477 = (reg437[(2'h3):(1'h0)] ? (!{(&(8'hb0))}) : (8'hba));
              reg478 <= $unsigned((^$signed(({(8'ha6), (8'hbd)} ?
                  reg448[(4'hb):(2'h3)] : {reg475}))));
              reg479 <= reg448[(5'h10):(4'h9)];
            end
          reg480 <= ($signed({((~&(8'had)) > $unsigned((8'hb3)))}) ?
              ({$unsigned((forvar473 >> wire387))} ?
                  (|reg416[(3'h6):(3'h5)]) : {$signed(reg476),
                      ($unsigned((8'hba)) ?
                          {reg396, wire400} : {reg442,
                              reg398})}) : $signed(reg461[(1'h1):(1'h1)]));
          reg481 <= $signed(($unsigned($signed($signed(reg408))) ?
              (~^{(reg465 != reg422)}) : reg396[(3'h6):(1'h1)]));
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned(reg448))
        begin
          if ($unsigned(((((~|reg398) >> wire470) && $signed(reg398[(5'h13):(4'h8)])) ?
              $signed(reg424[(1'h0):(1'h0)]) : $signed(reg437[(2'h2):(1'h0)]))))
            begin
              reg482 = $signed($signed((~^((reg466 ? reg451 : reg471) ?
                  $signed(reg428) : (reg466 ? reg472 : reg441)))));
            end
          else
            begin
              reg483 <= ($unsigned(reg422) < $unsigned((reg442 ~^ ((~|reg424) ^ $signed(reg480)))));
              reg484 = $unsigned($signed((7'h41)));
              reg485 <= reg401[(5'h12):(1'h1)];
              reg486 <= ($signed(reg417) == (+(^~($signed(reg437) ?
                  reg427 : (+(8'hb9))))));
              reg487 = $unsigned((~({reg427, $signed(reg391)} ?
                  ($signed(reg412) ?
                      reg428 : $signed(reg401)) : reg419[(4'hc):(3'h5)])));
            end
          reg488 = reg458;
        end
      else
        begin
          reg482 = $signed($signed(reg461[(2'h2):(1'h0)]));
          if ($signed($signed($signed((+(reg437 ? (8'hae) : wire388))))))
            begin
              reg484 = (!($unsigned((((7'h4a) == (8'h9f)) ?
                  $unsigned(reg482) : (reg453 == reg480))) >>> reg484));
              reg487 = ($signed((+($signed(reg391) ^ (~|reg488)))) ?
                  $signed({(8'hb1)}) : $signed((^~((~|wire386) <<< reg410[(3'h4):(3'h4)]))));
              reg489 <= $signed((-($signed((8'hbe)) != ((!reg458) + (^reg476)))));
            end
          else
            begin
              reg483 <= reg397;
              reg484 = reg488;
              reg487 = (-$unsigned(reg404[(1'h1):(1'h1)]));
              reg489 <= (reg447[(3'h7):(3'h6)] | (&wire470[(4'hf):(4'ha)]));
            end
          reg490 = (+$signed($unsigned(wire399[(1'h0):(1'h0)])));
          if ($unsigned(reg457[(2'h2):(1'h0)]))
            begin
              reg491 = ({$signed(((reg471 ? reg441 : reg398) ?
                          $unsigned((8'hbc)) : (reg416 ? reg465 : reg412))),
                      reg471[(5'h12):(5'h11)]} ?
                  (reg422[(1'h0):(1'h0)] ?
                      $signed($signed(reg482)) : reg403) : ($signed(wire400[(2'h2):(1'h0)]) ?
                      ($signed(reg466[(3'h4):(3'h4)]) || ((reg422 ?
                          reg415 : reg485) - (reg448 != reg447))) : reg446));
            end
          else
            begin
              reg491 = $unsigned((|($unsigned(reg461) ?
                  ((reg489 >= reg482) >= {reg458, reg466}) : (|{reg424,
                      reg404}))));
              reg492 = (({$unsigned((wire399 ? reg435 : reg476))} ?
                      (reg412 < ((8'ha6) ?
                          reg416[(2'h2):(1'h1)] : $signed(reg424))) : $signed($unsigned((~^(8'ha7))))) ?
                  (wire388[(1'h0):(1'h0)] == $signed({(wire400 ?
                          (8'hbe) : reg430)})) : $signed(reg407));
              reg493 = (reg415[(3'h4):(3'h4)] ?
                  $signed(wire400[(1'h1):(1'h0)]) : (7'h48));
            end
          reg494 <= $signed($unsigned(((^(reg485 ? (7'h46) : reg407)) ?
              reg489[(5'h14):(2'h3)] : {$signed(wire386)})));
        end
      reg495 <= ((8'hae) - (({$signed((8'hb6)),
              (wire470 ? reg403 : reg390)} | $unsigned((reg397 ?
              reg407 : reg472))) ?
          $unsigned((reg447 ?
              (reg483 ? wire388 : reg390) : (&reg417))) : reg484));
      reg496 = (&($signed((8'hbc)) ?
          (($unsigned((8'hb0)) ? (|reg487) : $unsigned(reg419)) ?
              (reg453 || ((8'hbe) ?
                  reg458 : reg398)) : wire400[(2'h2):(1'h0)]) : reg404));
    end
  always
    @(posedge clk) begin
      for (forvar497 = (1'h0); (forvar497 < (3'h4)); forvar497 = (forvar497 + (1'h1)))
        begin
          reg498 <= (~^reg396[(4'hc):(4'hb)]);
          if ((~&$unsigned((|((^reg404) ? reg428 : reg437)))))
            begin
              reg499 = $signed(reg398);
              reg500 = $signed(((((wire388 ? wire386 : wire389) ?
                      (reg430 + (8'hab)) : {reg430, reg447}) ?
                  {(reg479 >>> wire400),
                      $signed((8'ha8))} : {(~^reg481)}) == ($unsigned($signed(reg435)) | {reg415[(2'h2):(1'h0)],
                  $unsigned(reg412)})));
              reg501 = (((reg471 == reg410[(1'h1):(1'h0)]) ?
                  ((^~wire470[(3'h4):(1'h1)]) ?
                      $signed($unsigned(reg427)) : reg465) : (reg467 != ($unsigned(reg391) || reg498[(2'h3):(2'h3)]))) >> {reg390});
              reg502 = reg451;
            end
          else
            begin
              reg503 <= ($unsigned(($signed($signed(reg467)) ^ ($unsigned(reg457) ^~ reg500))) ?
                  reg415[(3'h6):(1'h1)] : (reg416[(4'hb):(1'h1)] ?
                      $unsigned(reg416) : ($unsigned($signed(wire389)) == (reg422 ?
                          wire400[(1'h1):(1'h1)] : (reg467 + reg500)))));
              reg504 <= reg415[(2'h2):(1'h1)];
              reg505 <= (~|(((reg458 ? reg419 : (^reg501)) ?
                      $unsigned((reg413 ?
                          (8'had) : wire387)) : ($unsigned(reg398) ?
                          (~^(7'h4a)) : (8'hbe))) ?
                  reg393 : $signed(reg407)));
              reg506 = {$signed(wire399),
                  $signed((reg401[(3'h6):(2'h2)] ~^ reg397[(1'h1):(1'h0)]))};
              reg507 <= {({(reg413[(3'h4):(1'h0)] * (8'hb1))} != reg502),
                  $unsigned(wire387)};
            end
          reg508 <= wire389;
          reg509 <= (reg415 ?
              $unsigned((7'h41)) : (reg472[(4'ha):(1'h0)] >> reg504));
          if (({$signed(wire470[(3'h7):(2'h2)]),
                  $signed($signed(reg508[(1'h0):(1'h0)]))} ?
              wire389[(2'h2):(2'h2)] : $signed(({(&reg465),
                  reg486} && (^(reg461 ? reg441 : reg427))))))
            begin
              reg510 = reg424[(4'hc):(3'h4)];
            end
          else
            begin
              reg511 <= reg506;
            end
        end
      reg512 = $unsigned((~|reg465[(1'h0):(1'h0)]));
      reg513 <= {{($unsigned(reg446[(3'h5):(2'h3)]) ?
                  {(!(7'h46)), reg419[(3'h6):(3'h5)]} : {(~reg419)}),
              $unsigned((((7'h41) ? reg509 : (8'hbb)) == (reg419 | reg481)))}};
    end
  assign wire514 = {reg461[(1'h1):(1'h0)]};
  assign wire515 = ((&(^~(7'h44))) < (&((8'hbf) ^~ $unsigned(reg498))));
  assign wire516 = {($unsigned(reg481[(2'h2):(1'h1)]) == ((reg508 & $unsigned((8'hb1))) ?
                           ($unsigned(reg508) ?
                               reg509[(4'hd):(3'h6)] : (8'hac)) : ((&(8'ha2)) ?
                               (reg413 ^ reg478) : $signed(reg413)))),
                       reg448[(4'h9):(4'h9)]};
  always
    @(posedge clk) begin
      for (forvar517 = (1'h0); (forvar517 < (2'h3)); forvar517 = (forvar517 + (1'h1)))
        begin
          if (reg466)
            begin
              reg518 <= wire386[(1'h1):(1'h0)];
              reg519 <= (($unsigned((&(^reg485))) ^~ $unsigned(($unsigned(reg472) >> ((8'ha1) ^~ wire515)))) ?
                  (reg472[(1'h0):(1'h0)] <<< ($signed((reg422 ?
                      reg507 : reg483)) + reg480)) : (!(reg503[(1'h1):(1'h0)] >= (8'h9d))));
              reg520 <= (reg396[(2'h2):(1'h0)] ?
                  {$signed((~reg410[(2'h2):(1'h1)]))} : forvar517);
            end
          else
            begin
              reg518 <= $unsigned($unsigned((+reg393[(2'h3):(1'h1)])));
            end
          for (forvar521 = (1'h0); (forvar521 < (1'h0)); forvar521 = (forvar521 + (1'h1)))
            begin
              reg522 = ((~(!$signed((wire386 << (7'h47))))) - $unsigned(reg403));
              reg523 <= (~^(|$unsigned(($unsigned(reg448) ?
                  (reg404 >= reg393) : reg416))));
            end
          reg524 <= reg410;
          reg525 <= $signed($unsigned(forvar521));
          if ((~$signed($signed((~{reg435, reg505})))))
            begin
              reg526 <= wire399;
              reg527 <= (~|(reg448 & ($unsigned((reg483 < reg518)) ?
                  $signed((wire386 << reg447)) : $unsigned((wire388 << (8'h9f))))));
              reg528 = reg441;
              reg529 <= (~&$signed(($unsigned($signed(wire470)) ?
                  {wire515} : (&(reg415 ? reg407 : (8'ha4))))));
              reg530 = reg478[(4'hc):(4'ha)];
            end
          else
            begin
              reg526 <= (&reg417);
              reg528 = reg401[(3'h5):(3'h4)];
            end
        end
      for (forvar531 = (1'h0); (forvar531 < (3'h4)); forvar531 = (forvar531 + (1'h1)))
        begin
          for (forvar532 = (1'h0); (forvar532 < (1'h1)); forvar532 = (forvar532 + (1'h1)))
            begin
              reg533 = (~reg401[(3'h7):(3'h5)]);
              reg534 = reg498;
              reg535 <= ({(~reg520)} ~^ reg505[(2'h2):(2'h2)]);
              reg536 = ($unsigned(($unsigned({reg404, reg505}) ?
                  $signed($unsigned(reg498)) : (~{reg483}))) != $unsigned((((~reg485) + reg495[(3'h7):(2'h2)]) <<< reg466[(3'h4):(1'h0)])));
            end
          for (forvar537 = (1'h0); (forvar537 < (1'h1)); forvar537 = (forvar537 + (1'h1)))
            begin
              reg538 <= reg480[(3'h4):(3'h4)];
              reg539 <= $signed((^~reg407[(3'h4):(2'h3)]));
              reg540 = (reg430 ?
                  $signed((!$signed((reg419 ? reg449 : (8'hb2))))) : (8'hbb));
            end
          reg541 = ($signed({wire386, ($signed(reg538) ^~ $signed(wire387))}) ?
              (((-(reg410 ?
                  reg446 : (7'h42))) ~^ $signed((!reg503))) ~^ reg422[(1'h1):(1'h0)]) : ((^reg430[(4'ha):(2'h2)]) & reg527));
          reg542 = ((!($unsigned(reg505[(3'h4):(2'h3)]) ?
              reg508[(3'h4):(2'h3)] : (8'hb2))) * (~&({reg466[(1'h0):(1'h0)],
                  $signed(reg508)} ?
              $unsigned(((7'h42) ? reg539 : reg442)) : $unsigned({reg541,
                  (8'hba)}))));
        end
    end
  always
    @(posedge clk) begin
      reg543 = (wire399[(1'h0):(1'h0)] ^ reg478);
    end
  assign wire544 = reg527[(3'h4):(1'h0)];
  assign wire545 = reg476;
  always
    @(posedge clk) begin
      reg546 = (~$unsigned((((reg453 & reg472) + reg413[(3'h7):(1'h1)]) ?
          reg448 : ($unsigned(reg525) ^~ $signed(reg539)))));
      if (((8'hae) ? reg524[(4'h8):(3'h7)] : $signed(reg485[(2'h2):(1'h0)])))
        begin
          reg547 = (reg401 ?
              ((reg523[(1'h0):(1'h0)] - (&$unsigned(reg498))) <<< (^$unsigned(reg508[(4'h9):(2'h2)]))) : reg407[(1'h1):(1'h1)]);
          if ((|reg447[(1'h1):(1'h1)]))
            begin
              reg548 = $signed(((~^$signed($unsigned(reg472))) + reg494));
              reg549 = reg430[(2'h2):(1'h1)];
              reg550 <= ((^(+$unsigned((|reg509)))) ?
                  $unsigned({((~|reg476) ? reg529 : (|reg422)),
                      (8'had)}) : (((^(reg391 ?
                      reg503 : reg508)) >> $signed(reg549)) ^ (&((~reg457) && $unsigned(reg539)))));
              reg551 <= (8'hae);
            end
          else
            begin
              reg548 = $unsigned(($signed((~|(reg539 - (8'ha5)))) ?
                  (&reg412[(1'h0):(1'h0)]) : (-{(^~(7'h42)), (^~reg413)})));
              reg549 = reg525[(3'h7):(3'h5)];
              reg552 = wire470;
              reg553 = (({(~^$signed(reg437))} << (!($unsigned(reg476) ?
                      $signed(reg481) : $signed((8'hb3))))) ?
                  (reg472[(3'h5):(2'h2)] ?
                      (|{reg489[(4'hb):(4'h9)]}) : ({{reg408}} <= wire515[(2'h3):(2'h3)])) : $signed((wire388[(4'h8):(3'h7)] & $unsigned(reg396[(1'h1):(1'h1)]))));
            end
          reg554 <= reg430;
        end
      else
        begin
          reg547 = $signed($unsigned($unsigned($signed({reg428}))));
          reg550 <= (reg448 ?
              (8'hb6) : (reg524 >= ((7'h49) != reg509[(4'ha):(3'h5)])));
          for (forvar551 = (1'h0); (forvar551 < (2'h2)); forvar551 = (forvar551 + (1'h1)))
            begin
              reg554 <= reg505[(2'h3):(1'h0)];
              reg555 = (reg509[(4'hc):(3'h6)] != reg478);
              reg556 <= reg408[(3'h4):(3'h4)];
              reg557 <= reg527;
            end
          for (forvar558 = (1'h0); (forvar558 < (2'h2)); forvar558 = (forvar558 + (1'h1)))
            begin
              reg559 <= $signed($unsigned((8'hae)));
            end
        end
      reg560 = (((^~$unsigned((reg546 ?
              reg403 : (8'hbb)))) > (~&(~^wire516[(4'h8):(3'h7)]))) ?
          $signed(reg559[(4'hb):(4'h9)]) : reg449[(2'h3):(1'h0)]);
    end
  assign wire561 = reg505[(1'h0):(1'h0)];
  assign wire562 = {reg397,
                       $signed(({(reg408 >>> reg526)} ?
                           $unsigned(wire544[(4'hf):(4'hb)]) : $signed((7'h40))))};
  always
    @(posedge clk) begin
      if ((~&wire388))
        begin
          if ($signed(reg451[(4'hc):(3'h5)]))
            begin
              reg563 <= (~&$unsigned((((reg550 >> reg397) ?
                  $unsigned(reg551) : reg498[(4'h8):(1'h1)]) >> ((^reg505) != (reg519 ?
                  (7'h48) : reg412)))));
              reg564 <= {((^~reg390) ?
                      $unsigned((8'hb5)) : $signed($unsigned($unsigned(reg529))))};
              reg565 <= $unsigned($unsigned(($signed(reg518) <= (~|(reg427 <= reg424)))));
              reg566 = ($unsigned(({reg486, $signed(reg480)} ?
                      (~|reg457[(2'h2):(1'h0)]) : ($unsigned(reg524) << (wire516 != reg520)))) ?
                  (($signed((~(8'hb4))) ^~ ((~^(8'hb4)) & $signed(reg479))) || ((~&(reg441 ?
                      wire561 : reg437)) * (reg447 >> reg412))) : {$signed($signed((reg391 <= reg513))),
                      (+reg563)});
              reg567 <= $signed(($signed(reg486[(2'h3):(2'h3)]) ?
                  reg403 : (~wire399[(1'h0):(1'h0)])));
            end
          else
            begin
              reg563 <= $unsigned($signed(reg461));
              reg566 = ((reg525[(1'h1):(1'h0)] ?
                  (~&{reg507}) : $unsigned(reg489)) ~^ reg467[(3'h7):(3'h6)]);
              reg568 = reg563[(2'h3):(2'h3)];
            end
        end
      else
        begin
          reg563 <= (({($signed(reg483) == reg504[(3'h5):(3'h4)]), reg523} ?
              {(~^(&(8'ha7))),
                  $unsigned((^(8'hb1)))} : ($unsigned(wire386[(3'h7):(3'h7)]) | reg403[(2'h2):(1'h0)])) <<< $unsigned((&((reg567 == reg483) ~^ $unsigned(reg557)))));
        end
      if (reg554[(3'h4):(2'h3)])
        begin
          reg569 = $signed((&({{(8'hbb), reg416}} ?
              (~^wire388[(4'ha):(4'ha)]) : $signed(reg483))));
          reg570 = $unsigned(reg441);
        end
      else
        begin
          if (((8'hbe) & ({reg478[(4'he):(3'h6)]} ?
              ((wire544[(1'h1):(1'h1)] ? reg554 : $unsigned(reg570)) ?
                  ((~reg509) & $unsigned(reg551)) : reg507[(4'h8):(2'h3)]) : (~&(~&$signed(reg559))))))
            begin
              reg569 = $unsigned((+reg461));
              reg571 <= $unsigned((~((~&$unsigned(reg419)) >= reg494)));
              reg572 = (^$signed(reg504[(3'h6):(1'h1)]));
            end
          else
            begin
              reg571 <= ($signed(((|(reg476 <<< wire388)) ?
                      $unsigned((wire399 & wire386)) : reg408[(3'h7):(3'h4)])) ?
                  reg563[(3'h6):(3'h4)] : (reg486[(4'h8):(2'h3)] ?
                      $unsigned($unsigned({(7'h44)})) : (reg466 ?
                          ((8'hb9) ?
                              $signed((8'hb9)) : $signed(wire516)) : (~&((8'ha4) ?
                              reg446 : reg485)))));
              reg573 <= ((&reg489[(3'h5):(2'h2)]) > $signed(reg480[(2'h3):(2'h2)]));
              reg574 <= (|$signed($unsigned(((8'hbb) << ((8'hae) ?
                  (8'had) : reg467)))));
              reg575 <= reg571;
              reg576 = reg503;
            end
          reg577 = reg401[(5'h17):(5'h12)];
          reg578 = $signed(reg437[(3'h6):(1'h0)]);
        end
      for (forvar579 = (1'h0); (forvar579 < (1'h0)); forvar579 = (forvar579 + (1'h1)))
        begin
          reg580 <= reg465[(2'h3):(1'h0)];
          if ((~|({(&(reg461 == reg538))} + (~|$unsigned($unsigned(reg571))))))
            begin
              reg581 = ($signed((({(8'hb3), reg416} <= {reg416,
                  reg524}) >>> {(~&reg573),
                  (reg479 - reg430)})) + ((-wire386[(2'h2):(1'h0)]) ?
                  (|(reg427[(1'h0):(1'h0)] | reg519)) : $signed(reg556)));
              reg582 = reg413[(2'h3):(1'h1)];
              reg583 <= {((~|(|wire562)) + reg410[(3'h4):(2'h3)]), reg576};
              reg584 <= (8'h9e);
              reg585 = reg401;
            end
          else
            begin
              reg581 = (reg523 | (($signed($unsigned(reg442)) << $signed(reg508)) < reg403[(1'h0):(1'h0)]));
            end
          reg586 = (reg393[(3'h5):(3'h4)] ?
              {(^~(~&$unsigned((8'hab)))),
                  $signed({reg538[(5'h10):(2'h3)],
                      reg503})} : (~&(~(reg441[(5'h11):(5'h11)] >>> (reg407 || reg580)))));
        end
    end
  assign wire587 = $unsigned($signed(($unsigned(wire389[(2'h2):(1'h0)]) >> ({reg565,
                       reg580} < (wire388 != reg574)))));
  always
    @(posedge clk) begin
      if ($unsigned($signed($unsigned(((~(8'h9f)) && (reg573 < reg401))))))
        begin
          reg588 = reg458;
          if ((((^~$unsigned(reg574[(3'h4):(2'h2)])) ?
              (~^{reg422[(3'h7):(1'h0)]}) : reg588) >> (|$unsigned((&$signed(reg495))))))
            begin
              reg589 <= ($unsigned(reg483) < {reg575});
              reg590 <= reg563[(3'h6):(3'h6)];
              reg591 <= {$unsigned((reg575[(3'h4):(1'h0)] && $unsigned($signed(reg504)))),
                  reg505};
              reg592 = reg503[(2'h3):(1'h0)];
              reg593 = {(^{(wire516 & (reg461 ? reg461 : reg390))}),
                  reg435[(1'h0):(1'h0)]};
            end
          else
            begin
              reg589 <= reg483;
            end
          for (forvar594 = (1'h0); (forvar594 < (2'h2)); forvar594 = (forvar594 + (1'h1)))
            begin
              reg595 = $unsigned($unsigned((reg412[(3'h4):(2'h2)] >> wire388)));
              reg596 = ($unsigned({$unsigned((reg451 ? (8'hbc) : reg476)),
                      reg442[(3'h7):(1'h0)]}) ?
                  (~^$signed(reg465[(1'h0):(1'h0)])) : {(-$unsigned(reg467))});
              reg597 <= ($unsigned((((reg485 ? reg415 : (7'h44)) + (-(8'hb3))) ?
                      $unsigned({reg573}) : reg494)) ?
                  $unsigned(reg494) : reg465[(1'h1):(1'h1)]);
              reg598 <= (^~$signed(({$signed(reg559), $signed(reg467)} ?
                  {(reg588 && wire562),
                      {reg417, wire516}} : reg509[(5'h10):(3'h4)])));
            end
        end
      else
        begin
          for (forvar588 = (1'h0); (forvar588 < (2'h3)); forvar588 = (forvar588 + (1'h1)))
            begin
              reg592 = (reg479 != {reg396});
              reg593 = reg571[(5'h13):(3'h5)];
            end
          reg594 <= ((8'hba) << $signed(({(reg390 ? wire470 : reg575),
                  reg593[(4'he):(1'h0)]} ?
              (reg449[(3'h6):(1'h0)] ^ (~|reg412)) : {reg393})));
          reg595 = reg485;
          if (reg446[(1'h0):(1'h0)])
            begin
              reg597 <= $signed(reg523[(4'h9):(1'h0)]);
              reg598 <= ((reg556[(2'h2):(2'h2)] ?
                  ((~reg589[(2'h2):(1'h0)]) ?
                      reg430 : reg494[(4'h9):(4'h9)]) : (8'haf)) <<< (reg539[(2'h2):(1'h1)] <= $signed($unsigned($signed(reg520)))));
              reg599 = (~($signed($unsigned($unsigned(reg525))) ?
                  ($unsigned((reg518 & reg589)) ?
                      $signed((reg513 ?
                          reg527 : reg435)) : (-(reg592 >> reg483))) : $unsigned($unsigned({reg404,
                      (8'ha3)}))));
            end
          else
            begin
              reg597 <= reg390[(1'h0):(1'h0)];
              reg598 <= ($signed((((reg599 | reg430) ? (|reg580) : {reg593}) ?
                  $unsigned($signed(reg503)) : $signed($unsigned(reg523)))) >>> $signed(((!reg554[(2'h3):(1'h1)]) << {reg598,
                  reg442[(4'ha):(3'h5)]})));
              reg599 = {wire545[(2'h3):(2'h3)],
                  $unsigned(reg592[(1'h1):(1'h1)])};
              reg600 = ($signed(reg518[(4'hf):(4'h9)]) ?
                  ({{reg538}, ({wire545} + (reg457 & reg504))} ?
                      reg458 : ((-(reg556 ? reg398 : reg465)) ?
                          $unsigned((reg538 + reg523)) : {reg594})) : $unsigned((reg523 ?
                      reg556 : $signed((8'ha6)))));
            end
          if ({wire544[(4'hf):(2'h3)],
              (((8'haa) != reg458) ?
                  (((forvar588 <= reg508) != reg494[(5'h14):(4'he)]) >> $signed({(8'hb2)})) : (reg448 * reg486[(3'h7):(1'h0)]))})
            begin
              reg601 <= reg449[(3'h4):(2'h3)];
              reg602 <= $unsigned((7'h48));
              reg603 = reg575;
              reg604 = (reg453 <= ((wire386[(4'h8):(4'h8)] * (-reg508)) || reg539));
              reg605 <= (~^(7'h42));
            end
          else
            begin
              reg601 <= $signed(reg415[(2'h3):(2'h3)]);
              reg602 <= ($signed($unsigned((|(reg481 ? reg428 : reg393)))) ?
                  (8'ha9) : reg591[(3'h5):(1'h1)]);
            end
        end
      if (reg556)
        begin
          reg606 <= {$unsigned((reg557 * $signed(reg424)))};
          reg607 = reg419;
          reg608 <= $signed($unsigned(wire388[(4'hf):(4'hb)]));
        end
      else
        begin
          reg607 = reg393[(3'h6):(1'h1)];
        end
      for (forvar609 = (1'h0); (forvar609 < (3'h4)); forvar609 = (forvar609 + (1'h1)))
        begin
          reg610 = $unsigned($signed(reg551[(2'h2):(1'h0)]));
        end
      if ($signed((&reg404)))
        begin
          if (({reg397} * ($signed(reg595[(2'h2):(2'h2)]) > $signed(reg550[(2'h2):(1'h0)]))))
            begin
              reg611 <= (~^reg495[(1'h0):(1'h0)]);
              reg612 = (|(((reg601 ?
                      (reg513 != reg481) : reg466[(2'h2):(2'h2)]) || $unsigned($signed(reg407))) ?
                  reg594[(3'h6):(3'h6)] : $signed(reg563)));
              reg613 = reg404;
            end
          else
            begin
              reg612 = (-$unsigned((|$unsigned((reg505 >> reg412)))));
              reg614 <= $unsigned((-$unsigned((~&((8'h9e) ?
                  reg613 : reg593)))));
              reg615 <= ((($signed(reg396[(4'hc):(4'hb)]) > $signed($unsigned(reg518))) ?
                  ({$signed(reg593)} >> (8'ha1)) : forvar594) && {reg580});
              reg616 <= ($unsigned($signed(reg458[(4'hf):(3'h5)])) ?
                  reg435[(2'h2):(1'h1)] : wire544[(1'h1):(1'h1)]);
            end
          reg617 = reg605;
        end
      else
        begin
          reg612 = reg457;
          if (reg396)
            begin
              reg614 <= (reg476[(3'h6):(3'h5)] * $unsigned(($unsigned(reg617) ?
                  reg485 : (^$unsigned(reg424)))));
              reg617 = $signed($signed((($signed(reg554) == $signed(wire561)) != $unsigned((wire587 & wire387)))));
              reg618 = reg447[(1'h1):(1'h0)];
              reg619 = ((((^~(-reg610)) != (((8'hb7) + (7'h46)) & wire545[(2'h2):(1'h0)])) ?
                  forvar588 : $signed({$unsigned(reg453),
                      (reg505 >>> (8'h9d))})) || (reg594 ^~ ($unsigned(reg618) >= $signed((~reg580)))));
            end
          else
            begin
              reg614 <= (8'hbb);
              reg617 = $unsigned($unsigned((reg604 ?
                  $unsigned((~^reg606)) : ($signed(reg527) ~^ (reg607 ?
                      (8'ha5) : reg526)))));
            end
          for (forvar620 = (1'h0); (forvar620 < (3'h4)); forvar620 = (forvar620 + (1'h1)))
            begin
              reg621 <= reg595[(2'h3):(1'h1)];
              reg622 <= {(wire544 == (^reg404[(3'h4):(1'h1)])),
                  ($unsigned(reg403[(1'h1):(1'h1)]) ?
                      {(forvar609 != reg494[(5'h10):(4'hf)]),
                          reg486[(1'h0):(1'h0)]} : ($unsigned(reg527) ~^ $signed($signed(reg599))))};
              reg623 <= $unsigned({(8'hb9),
                  $signed(((!reg559) - (reg415 > reg605)))});
              reg624 = $unsigned(reg461);
              reg625 <= $unsigned(reg471);
            end
          if ($signed((~|($signed($signed(reg397)) ^ reg413[(2'h2):(2'h2)]))))
            begin
              reg626 <= (reg498[(4'h9):(3'h4)] ?
                  $signed({$signed({reg580, reg419})}) : reg550);
              reg627 <= ($signed(reg422) ?
                  reg538 : ({(+(reg588 >> (8'hb3)))} ^ (7'h46)));
              reg628 <= (|(!reg626[(3'h6):(2'h3)]));
              reg629 <= ((reg413[(3'h4):(2'h3)] ?
                      ((~|$unsigned(reg625)) && $signed($unsigned((8'ha7)))) : (reg422 < {(reg476 || reg428)})) ?
                  $unsigned($signed(($unsigned(reg503) | {reg419,
                      reg427}))) : (~((~&reg580[(1'h0):(1'h0)]) ?
                      ({reg615, (8'hbd)} | (-wire470)) : reg498)));
            end
          else
            begin
              reg630 = reg616;
              reg631 <= (reg614 ?
                  (reg519[(5'h15):(5'h14)] ^~ $signed($signed(reg538))) : reg457[(3'h5):(1'h1)]);
              reg632 <= $unsigned($unsigned({(reg498[(1'h1):(1'h0)] > $signed(reg424)),
                  $signed(reg476[(3'h4):(2'h2)])}));
              reg633 <= $unsigned(reg574[(2'h3):(2'h2)]);
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed({reg446}))
        begin
          reg634 = (wire387[(3'h5):(2'h2)] || ((((reg621 ?
                  (8'hbc) : (8'hac)) + $signed(reg507)) > ((~^(8'haf)) | $unsigned(reg504))) ?
              reg584[(3'h4):(3'h4)] : (((reg551 >> (7'h47)) ?
                      reg574 : reg511[(2'h3):(2'h2)]) ?
                  $unsigned((wire515 ?
                      (7'h44) : reg498)) : ($unsigned(wire516) >> reg631[(4'h8):(1'h1)]))));
        end
      else
        begin
          reg634 = (|$signed((($unsigned(wire399) + $signed(reg554)) ?
              (&{reg461, (8'ha5)}) : $signed($signed(reg397)))));
        end
      for (forvar635 = (1'h0); (forvar635 < (1'h1)); forvar635 = (forvar635 + (1'h1)))
        begin
          for (forvar636 = (1'h0); (forvar636 < (3'h4)); forvar636 = (forvar636 + (1'h1)))
            begin
              reg637 <= ((wire389[(4'hc):(1'h0)] ?
                      $unsigned(reg538[(4'h8):(3'h4)]) : $unsigned(reg451)) ?
                  reg526 : $unsigned($unsigned(($unsigned(reg494) ?
                      reg435[(1'h0):(1'h0)] : (reg495 ? reg466 : reg526)))));
              reg638 = (!(~|$signed((reg611[(3'h4):(1'h0)] ^ ((8'ha5) ?
                  reg401 : reg511)))));
              reg639 = $signed({(~|$unsigned($unsigned(reg594))),
                  reg415[(3'h6):(2'h2)]});
              reg640 <= $signed((~|(8'hbd)));
              reg641 <= $unsigned($unsigned($signed((-$unsigned(reg480)))));
            end
          reg642 <= ((+$unsigned(({reg614} ?
              (reg471 ?
                  (8'hac) : (7'h43)) : $unsigned(reg626)))) | $unsigned((7'h48)));
          reg643 <= reg608;
          if (reg641[(3'h7):(3'h5)])
            begin
              reg644 <= reg527[(4'h9):(3'h7)];
              reg645 = reg605;
              reg646 = $signed($unsigned(reg594[(3'h7):(3'h5)]));
            end
          else
            begin
              reg645 = (reg638 >>> (((8'hac) - ((reg393 ?
                      reg614 : reg507) | $signed(reg550))) ?
                  {$unsigned(reg646)} : $unsigned((8'haf))));
              reg646 = reg448[(1'h1):(1'h0)];
              reg647 = reg614[(2'h2):(1'h0)];
              reg648 <= reg638;
            end
          for (forvar649 = (1'h0); (forvar649 < (2'h3)); forvar649 = (forvar649 + (1'h1)))
            begin
              reg650 <= reg503;
            end
        end
      reg651 = reg623[(1'h0):(1'h0)];
      for (forvar652 = (1'h0); (forvar652 < (2'h2)); forvar652 = (forvar652 + (1'h1)))
        begin
          reg653 = (reg645[(2'h2):(1'h0)] * (^$signed(wire400[(1'h1):(1'h1)])));
        end
    end
endmodule