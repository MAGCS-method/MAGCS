(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param264 = (!{{(((8'hb8) ? (8'hbd) : (8'h9f)) ? ((8'hae) <<< (8'hb2)) : (^(8'ha7)))}, (-({(8'ha1)} ? ((8'ha2) || (8'hba)) : ((8'had) <= (8'hb3))))}), 
parameter param265 = (8'hac))
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h342):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire4;
  input wire [(4'hb):(1'h0)] wire3;
  input wire signed [(4'h9):(1'h0)] wire2;
  input wire [(4'hc):(1'h0)] wire1;
  input wire [(2'h3):(1'h0)] wire0;
  wire signed [(3'h4):(1'h0)] wire263;
  wire [(4'he):(1'h0)] wire262;
  wire signed [(4'ha):(1'h0)] wire261;
  wire [(5'h12):(1'h0)] wire246;
  wire [(4'hc):(1'h0)] wire230;
  wire [(4'hd):(1'h0)] wire229;
  wire [(5'h15):(1'h0)] wire227;
  wire signed [(3'h7):(1'h0)] wire226;
  wire signed [(5'h15):(1'h0)] wire225;
  wire signed [(5'h13):(1'h0)] wire224;
  wire [(4'hc):(1'h0)] wire223;
  wire [(4'h9):(1'h0)] wire222;
  wire signed [(5'h14):(1'h0)] wire220;
  wire signed [(4'h8):(1'h0)] wire26;
  wire [(4'h9):(1'h0)] wire25;
  wire [(4'hb):(1'h0)] wire6;
  wire signed [(5'h11):(1'h0)] wire5;
  reg [(4'hc):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg259 = (1'h0);
  reg [(5'h13):(1'h0)] reg258 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg255 = (1'h0);
  reg [(4'hf):(1'h0)] reg253 = (1'h0);
  reg signed [(4'he):(1'h0)] reg251 = (1'h0);
  reg [(4'hc):(1'h0)] reg244 = (1'h0);
  reg [(4'hc):(1'h0)] reg240 = (1'h0);
  reg [(4'ha):(1'h0)] reg238 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg236 = (1'h0);
  reg [(5'h12):(1'h0)] reg233 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg232 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg231 = (1'h0);
  reg [(5'h12):(1'h0)] reg10 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg13 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg14 = (1'h0);
  reg [(5'h11):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg17 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg18 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg21 = (1'h0);
  reg [(3'h6):(1'h0)] reg24 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg [(4'he):(1'h0)] reg256 = (1'h0);
  reg [(4'hc):(1'h0)] reg254 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg252 = (1'h0);
  reg [(2'h3):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg249 = (1'h0);
  reg [(2'h3):(1'h0)] reg248 = (1'h0);
  reg [(5'h10):(1'h0)] reg247 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg245 = (1'h0);
  reg [(4'hb):(1'h0)] reg243 = (1'h0);
  reg [(5'h15):(1'h0)] reg242 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg241 = (1'h0);
  reg signed [(4'he):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg239 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg237 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar234 = (1'h0);
  reg [(3'h7):(1'h0)] reg7 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg23 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg19 = (1'h0);
  reg [(4'ha):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg9 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg8 = (1'h0);
  reg [(5'h14):(1'h0)] forvar7 = (1'h0);
  assign y = {wire263,
                 wire262,
                 wire261,
                 wire246,
                 wire230,
                 wire229,
                 wire227,
                 wire226,
                 wire225,
                 wire224,
                 wire223,
                 wire222,
                 wire220,
                 wire26,
                 wire25,
                 wire6,
                 wire5,
                 reg260,
                 reg259,
                 reg258,
                 reg255,
                 reg253,
                 reg251,
                 reg244,
                 reg240,
                 reg238,
                 reg236,
                 reg233,
                 reg232,
                 reg231,
                 reg10,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg21,
                 reg24,
                 reg257,
                 reg256,
                 reg254,
                 reg252,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg245,
                 reg243,
                 reg242,
                 reg241,
                 reg234,
                 reg239,
                 reg237,
                 reg235,
                 forvar234,
                 reg7,
                 reg23,
                 reg22,
                 reg20,
                 reg19,
                 reg11,
                 reg9,
                 reg8,
                 forvar7,
                 (1'h0)};
  assign wire5 = wire0;
  assign wire6 = {(((wire3[(3'h5):(3'h5)] == wire5[(4'ha):(3'h6)]) <<< ((wire4 ?
                             wire1 : wire4) == $unsigned((8'had)))) ?
                         (((wire4 ? wire2 : wire3) - wire5[(4'hd):(2'h2)]) ?
                             wire3[(3'h7):(1'h0)] : $signed((-wire0))) : ((~|wire0) ?
                             $unsigned(wire0[(1'h0):(1'h0)]) : $unsigned($signed((8'hba))))),
                     ($unsigned($signed($signed(wire4))) || wire5)};
  always
    @(posedge clk) begin
      if ($signed(wire3[(4'h8):(2'h3)]))
        begin
          for (forvar7 = (1'h0); (forvar7 < (3'h4)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg8 = wire6;
              reg9 = $signed(reg8[(1'h1):(1'h0)]);
              reg10 <= $signed(((((wire4 ? wire2 : (8'hb3)) ?
                      (wire0 != reg9) : {(8'hb8), reg8}) ?
                  wire2 : wire5[(4'hd):(1'h1)]) != wire0));
              reg11 = $signed((wire1 >= wire6[(1'h1):(1'h0)]));
            end
          if (reg9[(3'h5):(1'h1)])
            begin
              reg12 <= ((8'hb7) ^~ {((reg8 ? wire5 : (^reg9)) ?
                      (!$signed((8'ha0))) : $signed(wire2[(4'h9):(4'h9)])),
                  (wire0[(2'h2):(1'h1)] == wire2)});
              reg13 <= (forvar7 ? reg9 : {forvar7});
            end
          else
            begin
              reg12 <= reg8[(2'h2):(2'h2)];
              reg13 <= (&((&($unsigned(reg10) || (wire5 - wire5))) < $signed(((reg8 ?
                      wire0 : forvar7) ?
                  reg13[(1'h0):(1'h0)] : $unsigned(reg12)))));
            end
          reg14 <= $signed({$unsigned(($unsigned((8'ha2)) > $unsigned((7'h41))))});
          if (reg12)
            begin
              reg15 <= wire3;
              reg16 <= $signed($signed(((((7'h40) ? reg9 : wire4) ?
                      reg8 : (~&wire0)) ?
                  $unsigned({wire1}) : ($signed(wire4) ?
                      $unsigned(reg14) : (wire0 <= reg8)))));
              reg17 <= (wire1 ? $unsigned(forvar7[(5'h12):(3'h5)]) : reg10);
              reg18 <= $signed((reg17[(4'h9):(4'h9)] ?
                  $signed($unsigned((&reg12))) : (&reg11[(2'h2):(1'h0)])));
            end
          else
            begin
              reg19 = (~^(wire2 ? reg17[(1'h1):(1'h1)] : reg15));
              reg20 = $signed((($signed($unsigned(reg19)) ?
                      (reg17[(4'hd):(4'ha)] != {reg18}) : ((8'ha5) && reg8[(2'h3):(2'h3)])) ?
                  reg8 : $signed((reg8[(2'h2):(1'h1)] ?
                      $unsigned(forvar7) : $unsigned((8'hbb))))));
              reg21 <= ((reg20[(4'ha):(1'h1)] ?
                  (reg17 & $unsigned({reg9,
                      reg19})) : (~^(reg12[(2'h2):(1'h1)] ?
                      reg18[(3'h7):(3'h7)] : (wire3 ~^ wire5)))) >= reg17[(4'hf):(4'ha)]);
              reg22 = {wire0[(2'h2):(1'h1)]};
            end
          reg23 = reg10;
        end
      else
        begin
          reg7 = $unsigned($signed({(~|(7'h44)),
              {wire0[(1'h0):(1'h0)], {forvar7}}}));
        end
      reg24 <= ($unsigned((^~wire0[(1'h1):(1'h1)])) ?
          wire1 : wire5[(3'h6):(3'h6)]);
    end
  assign wire25 = ((wire6 ?
                      ($signed(reg10) ?
                          ((wire3 ? (7'h43) : wire2) ?
                              reg15[(3'h6):(3'h6)] : $signed(reg13)) : $signed((+(8'ha7)))) : reg12) < wire0);
  assign wire26 = reg17[(1'h1):(1'h1)];
  module27 #() modinst221 (.y(wire220), .wire32(reg16), .wire28(reg14), .clk(clk), .wire29(wire1), .wire30(reg21), .wire31(wire5));
  assign wire222 = $signed((^~wire0));
  assign wire223 = wire26;
  assign wire224 = (wire1[(3'h5):(1'h1)] ?
                       (~|(-wire0[(1'h1):(1'h0)])) : $signed({reg17,
                           $unsigned(wire6)}));
  assign wire225 = (reg12 <= reg21);
  assign wire226 = (wire223[(2'h2):(1'h1)] ^ ((reg17[(1'h0):(1'h0)] ?
                           $signed((wire1 ? wire220 : wire26)) : reg10) ?
                       wire222[(3'h6):(2'h2)] : $signed((^((8'h9e) <<< wire5)))));
  module56 #() modinst228 (.wire59(reg13), .wire60(reg16), .wire58(reg17), .wire57(reg14), .clk(clk), .y(wire227));
  assign wire229 = (reg21 >= $unsigned((+($signed(wire220) >>> reg15[(3'h4):(1'h0)]))));
  assign wire230 = $unsigned((($unsigned((reg24 ? reg16 : reg18)) ?
                           reg24[(2'h3):(1'h1)] : wire0[(2'h2):(1'h0)]) ?
                       ($signed((wire26 >= wire1)) - reg12) : wire223));
  always
    @(posedge clk) begin
      if ($signed(reg17))
        begin
          if ($unsigned(($unsigned(((~&(8'hbc)) && wire229)) & reg18)))
            begin
              reg231 <= (($signed($unsigned({reg21, wire0})) ?
                      $signed($signed(reg21)) : ($signed(wire2) || wire229)) ?
                  wire6[(4'h8):(1'h0)] : (wire0[(1'h0):(1'h0)] ?
                      $signed({$signed(reg16)}) : {((reg16 >>> reg13) >= (reg14 >= reg24)),
                          {(^(8'h9f)), reg14[(3'h5):(1'h1)]}}));
              reg232 <= wire26[(3'h5):(2'h2)];
              reg233 <= $signed($signed($signed($unsigned((wire226 != wire223)))));
            end
          else
            begin
              reg231 <= reg233[(4'hd):(4'h9)];
            end
          for (forvar234 = (1'h0); (forvar234 < (1'h0)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 = reg231;
              reg236 <= (reg18 && $unsigned((wire6[(4'ha):(1'h0)] ?
                  $unsigned((~^reg14)) : $unsigned($unsigned(wire26)))));
              reg237 = wire3[(4'hb):(3'h5)];
              reg238 <= $unsigned((((reg10 << (-(8'ha2))) <= (wire225 - (wire227 << reg237))) == ((8'haa) ?
                  (!$signed((8'hba))) : ($signed(wire229) < reg236[(1'h1):(1'h1)]))));
              reg239 = reg233;
            end
          reg240 <= {{wire3[(4'h9):(3'h6)], wire220}};
        end
      else
        begin
          reg234 = $unsigned(wire4);
          reg235 = reg10[(4'ha):(3'h4)];
          reg237 = $signed($unsigned({$unsigned(reg16[(5'h12):(4'hf)]),
              ($unsigned(reg12) ? $signed(wire25) : wire2)}));
          if (reg16)
            begin
              reg239 = ($signed(reg24[(2'h2):(2'h2)]) - (8'ha2));
              reg240 <= reg233[(3'h7):(3'h5)];
            end
          else
            begin
              reg239 = {wire4[(1'h1):(1'h1)]};
            end
        end
      if (reg237)
        begin
          reg241 = $unsigned(($unsigned((|reg16)) ?
              ($signed($signed(reg15)) >> wire227) : (-(8'haf))));
          reg242 = (~|reg234);
          reg243 = (8'hb5);
          reg244 <= (+(8'h9c));
        end
      else
        begin
          reg244 <= $unsigned(($unsigned((+$signed(wire25))) ?
              reg15[(4'hc):(3'h6)] : (~^$signed($signed(reg24)))));
          reg245 = (+wire227[(5'h11):(3'h7)]);
        end
    end
  assign wire246 = $unsigned(wire222);
  always
    @(posedge clk) begin
      if (reg17[(4'hc):(3'h6)])
        begin
          reg247 = (-reg18[(4'h9):(2'h3)]);
          reg248 = (&reg247[(1'h0):(1'h0)]);
          if (reg15[(4'hd):(3'h5)])
            begin
              reg249 = (|wire2);
              reg250 = ($signed($signed(reg233)) - ((!((reg18 == wire224) <<< {reg18})) || (wire229[(4'ha):(2'h3)] || reg232)));
            end
          else
            begin
              reg249 = wire0[(2'h3):(1'h1)];
              reg251 <= ((|{((^reg238) * $unsigned(reg248))}) != $signed((($signed(wire246) + (wire222 ^~ wire246)) ?
                  wire246[(2'h3):(1'h0)] : $unsigned($unsigned(reg240)))));
            end
          if ((reg236[(1'h0):(1'h0)] ~^ $unsigned((8'ha2))))
            begin
              reg252 = $signed((8'hba));
            end
          else
            begin
              reg253 <= wire5[(4'h9):(3'h4)];
              reg254 = (+$signed({reg249[(4'hb):(3'h6)]}));
              reg255 <= $unsigned(wire5[(1'h0):(1'h0)]);
            end
        end
      else
        begin
          if ((~^(!$signed({$signed(reg231), (reg252 & wire229)}))))
            begin
              reg251 <= wire225[(3'h6):(2'h3)];
            end
          else
            begin
              reg251 <= $unsigned($unsigned((8'hbc)));
              reg252 = $signed(reg247[(4'hc):(2'h3)]);
            end
          reg253 <= (|(reg244 ?
              ($signed((^~wire4)) ?
                  {reg248} : $signed((reg231 | reg24))) : reg10[(1'h1):(1'h0)]));
          if ($signed((+(&(-$signed(wire25))))))
            begin
              reg255 <= $signed(reg12[(4'h8):(3'h6)]);
              reg256 = wire2;
              reg257 = reg253;
            end
          else
            begin
              reg255 <= (~^$signed((+((~&reg14) ? reg10 : reg252))));
            end
        end
      reg258 <= (($signed((+$unsigned(wire226))) ?
          wire4 : {$signed($signed(reg18))}) * $unsigned(($unsigned(reg24[(1'h1):(1'h0)]) >> (!wire6))));
      reg259 <= ($unsigned(wire220) && wire246[(4'h9):(3'h4)]);
      reg260 <= ({(~|$signed((wire226 < reg15))),
          (~|$signed(reg231[(1'h1):(1'h0)]))} << (~^({$unsigned(wire1)} << $unsigned((reg15 ?
          reg231 : reg255)))));
    end
  assign wire261 = (~&reg12);
  assign wire262 = $unsigned($signed({wire220[(3'h4):(1'h0)]}));
  assign wire263 = {reg24,
                       {(($signed(wire224) ?
                               (reg18 >> reg16) : (reg13 ?
                                   reg233 : reg259)) | reg259),
                           {$unsigned({wire220}), {$unsigned(wire227)}}}};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module27
#(parameter param218 = ((((!((8'hac) <<< (8'ha8))) ? ((+(8'hab)) ~^ ((8'hab) | (7'h41))) : (^(^~(8'ha1)))) != ((~&((8'ha8) ? (8'ha4) : (8'h9e))) ? (((8'hb6) && (7'h41)) << {(8'h9f), (8'hb5)}) : ((8'h9e) || ((8'ha1) ^ (7'h40))))) >= (({((8'h9d) && (7'h41)), ((8'hb4) ? (8'ha0) : (8'ha6))} ? (~{(8'ha2)}) : (((8'ha7) != (8'hbe)) ~^ (~|(8'ha4)))) ? ((+((8'hb6) ^ (8'hb4))) ? ((~&(8'hb3)) ~^ (~^(8'hb7))) : (((8'hab) ? (8'hb2) : (8'hb2)) > (^(8'hb6)))) : {(((8'hbb) && (8'hbd)) ~^ ((8'hbb) ? (8'h9c) : (8'hb0))), (-((8'hb3) || (8'ha9)))})), 
parameter param219 = param218)
(y, clk, wire28, wire29, wire30, wire31, wire32);
  output wire [(32'h1c8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire28;
  input wire [(4'hc):(1'h0)] wire29;
  input wire [(3'h7):(1'h0)] wire30;
  input wire signed [(5'h10):(1'h0)] wire31;
  input wire signed [(5'h15):(1'h0)] wire32;
  wire [(3'h6):(1'h0)] wire216;
  wire [(2'h3):(1'h0)] wire215;
  wire signed [(5'h13):(1'h0)] wire214;
  wire signed [(3'h5):(1'h0)] wire213;
  wire [(4'ha):(1'h0)] wire212;
  wire [(5'h11):(1'h0)] wire211;
  wire signed [(2'h3):(1'h0)] wire210;
  wire signed [(3'h6):(1'h0)] wire209;
  wire signed [(4'hf):(1'h0)] wire208;
  wire signed [(2'h3):(1'h0)] wire207;
  wire [(5'h12):(1'h0)] wire206;
  wire signed [(4'hf):(1'h0)] wire205;
  wire [(2'h2):(1'h0)] wire204;
  wire [(4'hd):(1'h0)] wire203;
  wire [(3'h5):(1'h0)] wire201;
  reg [(5'h15):(1'h0)] reg217 = (1'h0);
  reg [(4'hf):(1'h0)] reg34 = (1'h0);
  reg [(4'hd):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg36 = (1'h0);
  reg [(4'hb):(1'h0)] reg37 = (1'h0);
  reg [(4'hc):(1'h0)] reg38 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg41 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg49 = (1'h0);
  reg [(5'h15):(1'h0)] reg51 = (1'h0);
  reg [(4'he):(1'h0)] reg53 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg54 = (1'h0);
  reg [(3'h7):(1'h0)] reg55 = (1'h0);
  reg [(4'hf):(1'h0)] reg52 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg50 = (1'h0);
  reg [(4'h9):(1'h0)] reg48 = (1'h0);
  reg [(5'h12):(1'h0)] reg47 = (1'h0);
  reg [(4'ha):(1'h0)] reg45 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg44 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar43 = (1'h0);
  reg [(4'he):(1'h0)] reg40 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg39 = (1'h0);
  reg [(5'h15):(1'h0)] forvar33 = (1'h0);
  assign y = {wire216,
                 wire215,
                 wire214,
                 wire213,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 wire208,
                 wire207,
                 wire206,
                 wire205,
                 wire204,
                 wire203,
                 wire201,
                 reg217,
                 reg34,
                 reg35,
                 reg36,
                 reg37,
                 reg38,
                 reg41,
                 reg42,
                 reg46,
                 reg49,
                 reg51,
                 reg53,
                 reg54,
                 reg55,
                 reg52,
                 reg50,
                 reg48,
                 reg47,
                 reg45,
                 reg44,
                 forvar43,
                 reg40,
                 reg39,
                 forvar33,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar33 = (1'h0); (forvar33 < (2'h3)); forvar33 = (forvar33 + (1'h1)))
        begin
          reg34 <= wire29[(2'h2):(1'h0)];
          if (wire28[(2'h2):(2'h2)])
            begin
              reg35 <= $unsigned(wire30[(3'h7):(2'h3)]);
              reg36 <= {($signed(({wire32, wire30} || {reg34,
                      (8'hab)})) * wire29),
                  (wire30 >= ($signed((~&reg34)) ?
                      ($unsigned(wire32) <= (~&wire31)) : (~^((8'ha6) ^ wire28))))};
              reg37 <= wire31;
              reg38 <= $signed(forvar33[(5'h14):(3'h6)]);
            end
          else
            begin
              reg39 = reg37[(4'h8):(3'h4)];
              reg40 = (-((!wire29) ^~ $signed(forvar33)));
              reg41 <= {(~|wire28)};
              reg42 <= {(8'hbc), wire28};
            end
          for (forvar43 = (1'h0); (forvar43 < (3'h4)); forvar43 = (forvar43 + (1'h1)))
            begin
              reg44 = (|($unsigned((8'hbb)) >= $unsigned($unsigned((~^wire30)))));
              reg45 = ((~^$unsigned($unsigned((forvar43 ?
                  reg39 : wire30)))) || (&$signed(wire30[(2'h3):(1'h1)])));
              reg46 <= (reg40 ?
                  $signed(wire32) : (wire31[(4'hd):(1'h0)] && (reg40 ?
                      (~^(8'hb1)) : $unsigned((reg39 ? reg35 : forvar43)))));
              reg47 = (wire31[(3'h7):(3'h5)] ?
                  (8'hba) : {reg34[(4'h9):(4'h8)]});
              reg48 = wire28;
            end
          if ((($unsigned({$unsigned(reg46), $signed(reg37)}) ?
              (($signed(reg48) ? (|reg40) : wire31[(1'h1):(1'h1)]) ?
                  ((^~reg35) & (reg38 >= (8'ha3))) : (-(reg36 || forvar43))) : (reg46 << (^wire28[(1'h1):(1'h1)]))) ^ ((wire30[(1'h1):(1'h0)] ?
                  ($signed(reg35) <<< $signed((8'ha2))) : $unsigned((~^wire31))) ?
              ((wire29 ?
                  (wire31 & reg47) : reg46) >>> {$unsigned((8'ha6))}) : $unsigned((~^$signed((8'hab)))))))
            begin
              reg49 <= reg47[(5'h12):(4'hf)];
              reg50 = (reg36[(1'h1):(1'h0)] != $signed(wire32[(5'h15):(3'h4)]));
              reg51 <= wire28;
              reg52 = ({$signed((&$unsigned(reg39))),
                  $unsigned({{reg49, (8'hba)}})} ^~ (reg42 ?
                  $signed(reg49[(1'h0):(1'h0)]) : (~|(reg40[(3'h5):(3'h4)] >= (reg45 ?
                      reg51 : (8'hb9))))));
              reg53 <= (-reg49);
            end
          else
            begin
              reg50 = $signed(wire31[(3'h7):(3'h4)]);
              reg52 = (~|(~|$signed(reg42[(2'h2):(1'h1)])));
              reg53 <= $signed((~^reg41[(4'hc):(1'h1)]));
              reg54 <= $signed(reg38[(4'hc):(4'h8)]);
            end
        end
      reg55 <= (!$unsigned((-(~|reg37[(4'ha):(4'h8)]))));
    end
  module56 #() modinst202 (wire201, clk, reg49, wire31, reg34, reg51);
  assign wire203 = ((wire28 ?
                           ($unsigned($unsigned(reg36)) ?
                               (^$signed(reg53)) : (+(wire30 >>> (8'haa)))) : (wire201[(2'h2):(2'h2)] ?
                               $unsigned((8'h9c)) : ((~|wire28) ?
                                   $signed(reg37) : $signed(wire201)))) ?
                       $unsigned(($unsigned((reg36 ?
                           wire201 : (8'hae))) + reg49[(3'h4):(2'h2)])) : ((((wire31 ~^ reg37) != $unsigned((8'ha6))) ?
                           wire29 : reg42[(3'h7):(3'h5)]) | $signed($unsigned($signed(wire201)))));
  assign wire204 = reg55;
  assign wire205 = (wire30 ? (!$signed({(~&reg53)})) : reg42[(2'h2):(2'h2)]);
  assign wire206 = {(8'hb8), reg46};
  assign wire207 = reg53[(4'hc):(4'h8)];
  assign wire208 = $unsigned(wire31);
  assign wire209 = reg34[(3'h6):(1'h0)];
  assign wire210 = (reg46[(3'h7):(2'h2)] ?
                       $unsigned($unsigned($signed(wire207[(1'h1):(1'h1)]))) : wire28[(1'h0):(1'h0)]);
  assign wire211 = $signed($signed((reg55[(3'h4):(2'h2)] ?
                       ((wire204 ? reg34 : wire207) ?
                           {wire29,
                               reg35} : $unsigned(reg36)) : reg55[(2'h3):(1'h0)])));
  assign wire212 = reg54[(3'h5):(3'h4)];
  assign wire213 = $signed((!wire205[(4'hc):(4'ha)]));
  assign wire214 = $signed(reg55[(3'h5):(3'h4)]);
  assign wire215 = (~($signed((((8'hb3) ? wire28 : reg38) ?
                           (wire211 && reg55) : $unsigned(reg38))) ?
                       $unsigned((reg35[(4'ha):(4'h9)] <= reg51)) : $signed(reg49[(2'h3):(1'h1)])));
  assign wire216 = (((($signed(wire211) >>> $signed(reg35)) ?
                           wire208 : $signed(reg34[(2'h3):(2'h2)])) > ((wire207 >>> reg35) ~^ (~|reg34))) ?
                       $unsigned((^$signed((|reg54)))) : wire201[(2'h3):(2'h2)]);
  always
    @(posedge clk) begin
      reg217 <= (wire213[(1'h0):(1'h0)] - $signed($unsigned($signed(wire201[(2'h2):(1'h0)]))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module56
#(parameter param199 = {(8'haa)}, 
parameter param200 = ((~|{{(~param199), param199}}) - (~&(((param199 || param199) ? (param199 || param199) : param199) >= param199))))
(y, clk, wire60, wire59, wire58, wire57);
  output wire [(32'h167):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire60;
  input wire signed [(5'h10):(1'h0)] wire59;
  input wire signed [(4'hc):(1'h0)] wire58;
  input wire [(4'ha):(1'h0)] wire57;
  wire signed [(3'h4):(1'h0)] wire198;
  wire [(5'h14):(1'h0)] wire196;
  wire signed [(5'h10):(1'h0)] wire107;
  wire signed [(4'hd):(1'h0)] wire106;
  wire [(5'h11):(1'h0)] wire104;
  wire signed [(5'h15):(1'h0)] wire81;
  wire signed [(3'h6):(1'h0)] wire80;
  wire [(4'h8):(1'h0)] wire79;
  wire signed [(2'h3):(1'h0)] wire78;
  wire signed [(5'h13):(1'h0)] wire77;
  wire signed [(4'he):(1'h0)] wire76;
  wire signed [(5'h13):(1'h0)] wire75;
  wire signed [(5'h11):(1'h0)] wire74;
  reg signed [(5'h13):(1'h0)] reg62 = (1'h0);
  reg [(5'h11):(1'h0)] reg63 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg66 = (1'h0);
  reg [(4'hc):(1'h0)] reg68 = (1'h0);
  reg [(3'h7):(1'h0)] reg71 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg67 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg70 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar67 = (1'h0);
  reg [(5'h12):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg61 = (1'h0);
  assign y = {wire198,
                 wire196,
                 wire107,
                 wire106,
                 wire104,
                 wire81,
                 wire80,
                 wire79,
                 wire78,
                 wire77,
                 wire76,
                 wire75,
                 wire74,
                 reg62,
                 reg63,
                 reg64,
                 reg66,
                 reg68,
                 reg71,
                 reg67,
                 reg72,
                 reg73,
                 reg70,
                 reg69,
                 forvar67,
                 reg65,
                 reg61,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg61 = (~(8'hb7));
      if ({(wire60[(5'h10):(3'h5)] ?
              ((8'hb6) ?
                  (-$unsigned(wire60)) : $signed(wire57[(3'h5):(2'h2)])) : {$signed((reg61 & wire57))})})
        begin
          if ($signed(wire60))
            begin
              reg62 <= {(-wire60)};
              reg63 <= reg61;
              reg64 <= (({((reg61 ? wire57 : (8'haa)) || (^~reg62)),
                      (-$signed(reg63))} <<< $signed($unsigned(wire60))) ?
                  $signed({(~wire59), wire57}) : (~|(^reg61[(4'he):(3'h6)])));
            end
          else
            begin
              reg62 <= ($signed(((~(|reg62)) - $signed(reg64[(4'h8):(3'h5)]))) & ($signed($signed(reg64[(3'h7):(2'h3)])) ?
                  $unsigned($unsigned($unsigned(reg62))) : (+reg64[(3'h7):(3'h7)])));
              reg65 = {reg61};
              reg66 <= (!(|$unsigned((~^(reg65 >>> (8'hbd))))));
            end
          for (forvar67 = (1'h0); (forvar67 < (2'h3)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 <= (((|$unsigned($signed(wire57))) >>> reg61[(1'h1):(1'h1)]) * wire59);
            end
          if (((reg68 ?
              $signed($signed((^wire59))) : ((reg65[(3'h5):(1'h1)] ?
                  reg63[(4'hd):(4'hb)] : $signed(wire59)) || wire57)) == $unsigned(wire58[(3'h7):(2'h2)])))
            begin
              reg69 = reg64[(3'h7):(3'h6)];
              reg70 = ((~$signed(({wire60, reg69} ? wire58 : (~&reg61)))) ?
                  $signed(((reg64[(2'h3):(2'h2)] ?
                          reg63[(1'h1):(1'h1)] : forvar67) ?
                      $signed((reg62 ^~ reg63)) : reg61)) : wire59[(2'h2):(1'h0)]);
            end
          else
            begin
              reg71 <= reg70;
            end
        end
      else
        begin
          if (reg62)
            begin
              reg62 <= ((-($unsigned((|reg68)) ?
                  reg63[(4'hc):(4'hc)] : reg63)) <<< (!$signed(((reg68 ?
                  wire60 : reg66) >= $unsigned((8'hbf))))));
              reg65 = $signed($unsigned(reg62));
              reg66 <= {({reg62, $unsigned(reg63[(3'h5):(2'h3)])} ?
                      (^(~|{reg61, reg61})) : (&(+(reg62 ? reg69 : reg66)))),
                  ($unsigned($unsigned({wire59, reg64})) ?
                      $unsigned(reg61[(5'h11):(3'h5)]) : wire59[(3'h5):(3'h5)])};
              reg67 <= (&((($unsigned(reg71) >>> reg70[(5'h11):(3'h6)]) ?
                  (reg71 ?
                      (reg68 ^~ reg62) : {(8'h9e),
                          reg66}) : reg65) || $signed((8'ha5))));
            end
          else
            begin
              reg62 <= (~^(reg71 ? (|reg71[(3'h7):(1'h0)]) : reg70));
            end
          if ((wire58 ?
              $unsigned((~reg63[(3'h4):(2'h2)])) : $signed($unsigned({(wire57 || (8'ha5)),
                  $signed(reg65)}))))
            begin
              reg69 = (reg61 > $unsigned((($unsigned(reg68) > (~forvar67)) * reg65)));
              reg70 = (~|$signed((((7'h44) ~^ {reg65, reg65}) ?
                  ((&(8'ha8)) | reg68[(4'h8):(4'h8)]) : (+(!reg63)))));
              reg71 <= reg71;
              reg72 <= wire60;
              reg73 <= (8'hb6);
            end
          else
            begin
              reg69 = $unsigned($unsigned($signed((((8'ha4) ? wire60 : wire59) ?
                  $signed(reg69) : $unsigned(reg71)))));
              reg71 <= (((~&reg68[(3'h5):(3'h5)]) << {$signed(forvar67[(4'h9):(3'h5)]),
                      (|(wire57 ? wire60 : reg70))}) ?
                  (~wire60) : wire60);
            end
        end
    end
  assign wire74 = $unsigned(((|reg71) * reg72[(4'hd):(2'h2)]));
  assign wire75 = (((reg62[(3'h5):(3'h4)] ? (~^reg71) : reg62) ?
                      (wire57[(4'ha):(3'h7)] >>> $unsigned(wire58[(3'h6):(3'h6)])) : wire60) << reg73[(1'h0):(1'h0)]);
  assign wire76 = (((~&wire60[(4'hf):(2'h3)]) - $unsigned((-$signed(reg67)))) ?
                      reg72[(3'h5):(1'h0)] : reg62[(3'h4):(1'h1)]);
  assign wire77 = {wire76};
  assign wire78 = (~&{$signed($signed($signed(wire77)))});
  assign wire79 = (~(~{((reg73 ? reg73 : wire77) ?
                          reg66[(4'hc):(4'h8)] : wire77[(5'h10):(3'h4)]),
                      reg63}));
  assign wire80 = reg62;
  assign wire81 = wire57;
  module82 #() modinst105 (.wire86(wire76), .wire85(wire60), .y(wire104), .clk(clk), .wire83(wire74), .wire84(wire58));
  assign wire106 = (-reg67[(2'h3):(2'h2)]);
  assign wire107 = ($signed(wire75) ? (7'h44) : reg71[(3'h7):(3'h6)]);
  module108 #() modinst197 (.wire109(wire81), .wire113(wire74), .y(wire196), .wire110(wire75), .clk(clk), .wire112(wire76), .wire111(reg72));
  assign wire198 = (+(~|(((wire59 ? wire81 : wire74) ?
                       (~reg73) : $signed(wire77)) < $signed($signed(wire107)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module108
#(parameter param195 = (~^(&((((8'h9c) ? (8'hb8) : (7'h43)) || {(8'hbb), (8'hb7)}) ? ({(8'ha8), (8'hb0)} ? (-(8'ha6)) : {(7'h40)}) : (8'ha8)))))
(y, clk, wire113, wire112, wire111, wire110, wire109);
  output wire [(32'h3c5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire113;
  input wire [(3'h7):(1'h0)] wire112;
  input wire [(3'h6):(1'h0)] wire111;
  input wire signed [(5'h13):(1'h0)] wire110;
  input wire [(5'h15):(1'h0)] wire109;
  wire [(5'h10):(1'h0)] wire192;
  wire signed [(5'h15):(1'h0)] wire191;
  wire signed [(5'h15):(1'h0)] wire190;
  wire signed [(4'hf):(1'h0)] wire189;
  wire [(3'h7):(1'h0)] wire188;
  wire [(4'h8):(1'h0)] wire187;
  wire [(3'h5):(1'h0)] wire147;
  wire signed [(5'h14):(1'h0)] wire146;
  wire [(3'h7):(1'h0)] wire145;
  wire signed [(4'hf):(1'h0)] wire144;
  wire signed [(2'h3):(1'h0)] wire143;
  wire signed [(3'h4):(1'h0)] wire142;
  wire signed [(4'hc):(1'h0)] wire141;
  wire signed [(3'h4):(1'h0)] wire140;
  wire signed [(4'ha):(1'h0)] wire139;
  wire [(5'h15):(1'h0)] wire138;
  wire signed [(5'h10):(1'h0)] wire137;
  wire [(4'hf):(1'h0)] wire136;
  wire [(5'h15):(1'h0)] wire135;
  wire [(5'h12):(1'h0)] wire134;
  reg signed [(2'h3):(1'h0)] reg186 = (1'h0);
  reg [(5'h11):(1'h0)] reg185 = (1'h0);
  reg [(4'h9):(1'h0)] reg183 = (1'h0);
  reg [(5'h10):(1'h0)] reg182 = (1'h0);
  reg [(3'h7):(1'h0)] reg179 = (1'h0);
  reg [(4'hd):(1'h0)] reg175 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg174 = (1'h0);
  reg signed [(4'he):(1'h0)] reg173 = (1'h0);
  reg [(5'h11):(1'h0)] reg171 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg163 = (1'h0);
  reg [(4'hc):(1'h0)] reg161 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg157 = (1'h0);
  reg [(2'h3):(1'h0)] reg155 = (1'h0);
  reg [(4'ha):(1'h0)] reg153 = (1'h0);
  reg [(4'hd):(1'h0)] reg150 = (1'h0);
  reg [(5'h14):(1'h0)] reg148 = (1'h0);
  reg [(4'hc):(1'h0)] reg131 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg130 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg126 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg118 = (1'h0);
  reg [(5'h12):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg194 = (1'h0);
  reg [(2'h3):(1'h0)] reg193 = (1'h0);
  reg [(4'h8):(1'h0)] reg184 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg181 = (1'h0);
  reg [(5'h13):(1'h0)] reg180 = (1'h0);
  reg [(4'hc):(1'h0)] reg178 = (1'h0);
  reg [(3'h4):(1'h0)] reg177 = (1'h0);
  reg [(4'hd):(1'h0)] reg176 = (1'h0);
  reg [(4'hf):(1'h0)] reg172 = (1'h0);
  reg [(4'h8):(1'h0)] reg170 = (1'h0);
  reg [(4'hd):(1'h0)] reg169 = (1'h0);
  reg [(5'h10):(1'h0)] reg168 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar165 = (1'h0);
  reg [(2'h2):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg162 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar160 = (1'h0);
  reg [(4'hb):(1'h0)] reg159 = (1'h0);
  reg [(2'h3):(1'h0)] reg158 = (1'h0);
  reg [(4'he):(1'h0)] reg156 = (1'h0);
  reg [(4'h9):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg151 = (1'h0);
  reg [(2'h3):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg132 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg129 = (1'h0);
  reg [(3'h5):(1'h0)] reg127 = (1'h0);
  reg [(4'h9):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg123 = (1'h0);
  reg [(5'h11):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg121 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg119 = (1'h0);
  reg [(3'h5):(1'h0)] reg117 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg116 = (1'h0);
  reg [(5'h14):(1'h0)] reg114 = (1'h0);
  assign y = {wire192,
                 wire191,
                 wire190,
                 wire189,
                 wire188,
                 wire187,
                 wire147,
                 wire146,
                 wire145,
                 wire144,
                 wire143,
                 wire142,
                 wire141,
                 wire140,
                 wire139,
                 wire138,
                 wire137,
                 wire136,
                 wire135,
                 wire134,
                 reg186,
                 reg185,
                 reg183,
                 reg182,
                 reg179,
                 reg175,
                 reg174,
                 reg173,
                 reg171,
                 reg167,
                 reg163,
                 reg161,
                 reg157,
                 reg155,
                 reg153,
                 reg150,
                 reg148,
                 reg131,
                 reg130,
                 reg128,
                 reg126,
                 reg124,
                 reg120,
                 reg118,
                 reg115,
                 reg194,
                 reg193,
                 reg184,
                 reg181,
                 reg180,
                 reg178,
                 reg177,
                 reg176,
                 reg172,
                 reg170,
                 reg169,
                 reg168,
                 reg166,
                 forvar165,
                 reg164,
                 reg162,
                 forvar160,
                 reg159,
                 reg158,
                 reg156,
                 reg154,
                 reg152,
                 reg151,
                 reg149,
                 reg133,
                 reg132,
                 reg129,
                 reg127,
                 reg125,
                 reg123,
                 reg122,
                 reg121,
                 reg119,
                 reg117,
                 reg116,
                 reg114,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned(wire110))
        begin
          if ((~$unsigned((wire113[(4'h8):(1'h0)] ?
              (^~((8'ha3) == wire109)) : ($signed(wire109) != (~&wire113))))))
            begin
              reg114 = (^~((^~$signed(wire109)) ?
                  wire112 : (~$unsigned((&wire109)))));
              reg115 <= wire109;
              reg116 = wire109;
              reg117 = wire112;
              reg118 <= wire113[(1'h1):(1'h1)];
            end
          else
            begin
              reg114 = ({wire110} && $unsigned((^~$unsigned($signed(reg115)))));
              reg116 = reg116[(1'h0):(1'h0)];
              reg118 <= ($unsigned((reg114 & (&(-reg117)))) < wire110);
            end
          if (($signed($signed({(-reg117)})) ^~ $signed(reg115)))
            begin
              reg119 = $signed(wire110[(4'hb):(4'h9)]);
              reg120 <= reg119[(2'h2):(1'h1)];
              reg121 = {{($signed($signed(reg116)) ?
                          ($signed(wire111) == reg117) : wire113)},
                  ($signed($signed((reg115 << wire112))) ?
                      $unsigned(((8'hbe) - wire109[(4'he):(2'h3)])) : $unsigned($unsigned(reg115[(5'h12):(4'ha)])))};
              reg122 = (+(&(((wire110 > wire113) ?
                      (-(8'ha3)) : reg119[(2'h2):(1'h1)]) ?
                  $unsigned((reg114 ?
                      reg115 : wire113)) : reg120[(2'h2):(1'h1)])));
              reg123 = $unsigned(reg114);
            end
          else
            begin
              reg120 <= (^~reg118);
              reg121 = ($signed((((~^reg123) <= $signed(reg114)) ?
                  reg122[(4'hf):(3'h7)] : $unsigned(((8'h9c) <<< (8'hbd))))) <<< $unsigned({((8'hb6) > $unsigned(reg121)),
                  ((reg117 ? wire111 : (8'ha6)) != wire109)}));
            end
          if (reg121[(4'ha):(3'h5)])
            begin
              reg124 <= wire111;
            end
          else
            begin
              reg125 = $signed({reg124, $signed(reg120)});
              reg126 <= wire111;
              reg127 = ($signed($signed(((reg118 == reg124) > ((8'hbb) << wire113)))) - reg122[(2'h3):(2'h3)]);
              reg128 <= $unsigned(((-{reg122[(4'h9):(1'h0)],
                  $signed(reg127)}) * reg124));
              reg129 = reg123[(4'h8):(2'h2)];
            end
          reg130 <= (~^$unsigned(reg128[(2'h3):(1'h1)]));
          if ((reg121 ?
              reg114[(4'hc):(4'ha)] : (reg129[(4'h9):(3'h7)] ?
                  (8'h9f) : reg124)))
            begin
              reg131 <= reg130;
              reg132 = (reg120 ?
                  ((reg120[(3'h5):(3'h5)] ?
                      $unsigned(reg128[(1'h1):(1'h0)]) : $unsigned((reg124 || (8'h9d)))) - (reg115 ?
                      $signed(reg119) : $signed((-reg131)))) : reg122[(5'h11):(4'hb)]);
              reg133 = (($signed((&(reg132 << (8'ha2)))) != (((~&reg125) >= $signed(reg130)) ^~ ($signed(reg132) >>> reg124[(4'hf):(3'h7)]))) >>> $unsigned(reg122[(3'h5):(3'h5)]));
            end
          else
            begin
              reg131 <= reg124;
            end
        end
      else
        begin
          if (reg125[(2'h3):(2'h2)])
            begin
              reg115 <= $signed(reg118[(2'h3):(1'h1)]);
              reg116 = ($unsigned(($unsigned((reg116 == wire112)) ?
                  $unsigned((~&(8'h9e))) : ((~^reg115) ^ (reg126 ?
                      (8'hab) : reg133)))) ^ (reg132 ?
                  $signed((&(reg132 || reg122))) : reg114));
              reg117 = {$unsigned(($signed($unsigned(reg123)) ?
                      {reg122, reg132[(3'h4):(1'h1)]} : reg129))};
              reg118 <= (!$signed($signed(reg122)));
            end
          else
            begin
              reg114 = $unsigned((^(~|reg114[(3'h5):(3'h5)])));
              reg115 <= wire111;
              reg118 <= ($unsigned(($signed(reg132) ?
                  (-(reg120 ?
                      reg133 : reg122)) : ((reg118 && reg116) << $signed(reg120)))) <<< $signed((reg132[(3'h4):(2'h2)] ^~ reg118[(3'h4):(1'h1)])));
              reg119 = reg131;
              reg120 <= reg122;
            end
          reg121 = $unsigned(reg120);
          reg124 <= (+reg121[(1'h0):(1'h0)]);
        end
    end
  assign wire134 = ($signed($signed(((^~(8'ha7)) ?
                       (^reg130) : (reg131 ? reg131 : wire109)))) ^ (7'h42));
  assign wire135 = ((((reg115 * (reg124 & reg128)) ?
                               (reg131[(3'h7):(2'h2)] ~^ $unsigned((8'hac))) : (|$signed(reg130))) ?
                           (8'hb7) : ((!$unsigned(reg115)) ?
                               wire111[(3'h6):(2'h2)] : reg130)) ?
                       (({$signed(reg128),
                               reg120[(2'h2):(1'h1)]} == $unsigned(wire109[(5'h14):(2'h2)])) ?
                           (wire111 + wire112) : wire109) : wire113[(2'h2):(1'h1)]);
  assign wire136 = ((((8'h9c) ?
                           wire134 : ((reg130 < wire112) ?
                               $signed(wire134) : {(8'ha1)})) ^~ ($signed($signed(reg126)) || (~^(+wire110)))) ?
                       reg130[(3'h4):(2'h3)] : (!(wire112 ?
                           ($signed(reg130) <<< (reg120 ?
                               reg118 : wire110)) : $signed(reg131[(4'h8):(2'h2)]))));
  assign wire137 = $signed((wire136[(4'hc):(4'ha)] || wire110));
  assign wire138 = (({$unsigned(wire109[(4'h8):(2'h2)])} ?
                           {reg130[(4'h9):(3'h6)],
                               $unsigned((&(8'hac)))} : wire113) ?
                       (^({(wire137 << wire136), (reg120 ? (8'hb4) : reg128)} ?
                           ((wire134 ?
                               (8'ha0) : (8'hb7)) + ((8'hae) >>> reg131)) : (-{reg120,
                               (8'hb0)}))) : reg128[(1'h1):(1'h1)]);
  assign wire139 = $unsigned({(^~(~&$signed(reg118))),
                       (^$signed($signed(wire138)))});
  assign wire140 = ({$signed(wire137)} ?
                       $signed((($unsigned(wire135) ?
                               $signed((8'hb3)) : {wire139, wire134}) ?
                           wire113 : $signed(((8'haf) - reg130)))) : (&((~(^~reg115)) ?
                           ($unsigned((8'hb5)) ?
                               (wire139 ?
                                   wire111 : wire111) : wire109[(3'h4):(2'h2)]) : wire139)));
  assign wire141 = (8'ha8);
  assign wire142 = (wire113[(3'h7):(2'h3)] || ($signed(wire134[(2'h3):(2'h2)]) ?
                       $signed((|$signed(reg130))) : $unsigned((+$unsigned(wire113)))));
  assign wire143 = (!$unsigned(($signed(((8'ha8) ?
                       reg124 : reg115)) & wire140[(1'h0):(1'h0)])));
  assign wire144 = $signed({(reg131[(3'h5):(2'h3)] ?
                           ($unsigned(reg118) ?
                               ((8'h9c) <= (8'hbf)) : wire136) : ((wire134 ?
                                   wire137 : (8'hb2)) ?
                               (wire143 ?
                                   reg124 : wire142) : (wire141 >>> reg124))),
                       $signed((|$unsigned(wire143)))});
  assign wire145 = $unsigned(wire144);
  assign wire146 = $signed((~|reg126[(4'hc):(3'h6)]));
  assign wire147 = ($unsigned(wire144[(3'h7):(3'h4)]) ?
                       ((!(~|(~&reg115))) ?
                           $signed(((wire111 ?
                               wire134 : wire140) * $signed(wire111))) : $signed(({(8'hb4)} ?
                               (wire135 & reg126) : (reg120 ^ reg131)))) : $unsigned((7'h42)));
  always
    @(posedge clk) begin
      if ((8'h9e))
        begin
          if (wire145[(3'h7):(2'h2)])
            begin
              reg148 <= wire113;
              reg149 = ($signed(($unsigned((reg131 << wire135)) ?
                  $unsigned((wire139 * wire146)) : (wire147[(3'h4):(1'h1)] ?
                      ((8'hb8) ?
                          wire109 : wire139) : $signed(reg124)))) + {reg126,
                  wire113[(4'h8):(3'h5)]});
              reg150 <= (8'hbe);
              reg151 = reg115;
            end
          else
            begin
              reg149 = wire143[(1'h0):(1'h0)];
            end
          if ($unsigned(($unsigned({wire112[(3'h4):(3'h4)]}) ^~ $signed((reg124[(4'hb):(4'h8)] < wire110)))))
            begin
              reg152 = $unsigned(reg124[(3'h5):(3'h5)]);
              reg153 <= wire138;
            end
          else
            begin
              reg152 = reg131[(2'h3):(2'h2)];
              reg154 = {(^$unsigned((!$unsigned(wire141))))};
            end
          if ({$unsigned((~^(wire145 ?
                  wire138[(4'hd):(3'h4)] : ((8'ha8) >>> (8'ha0))))),
              (-wire140[(3'h4):(1'h0)])})
            begin
              reg155 <= ((+((&(8'haf)) | $signed({wire112}))) ?
                  wire142[(2'h2):(1'h0)] : (wire109 ?
                      $unsigned(wire135[(2'h3):(2'h2)]) : (wire144[(2'h3):(1'h1)] ?
                          $unsigned(wire111) : reg153)));
              reg156 = $signed((^$unsigned($signed((reg153 ?
                  wire110 : wire139)))));
            end
          else
            begin
              reg155 <= $signed(reg149[(1'h1):(1'h0)]);
              reg157 <= $signed((^~(~$signed($signed(wire138)))));
              reg158 = reg149[(2'h3):(1'h1)];
            end
          reg159 = reg131;
          for (forvar160 = (1'h0); (forvar160 < (1'h1)); forvar160 = (forvar160 + (1'h1)))
            begin
              reg161 <= (~reg124);
              reg162 = wire144;
              reg163 <= $unsigned({reg120[(1'h1):(1'h0)],
                  $signed(((reg158 ? wire144 : wire110) ?
                      {(8'ha5)} : $signed(reg148)))});
              reg164 = (^{reg155[(2'h2):(2'h2)]});
            end
        end
      else
        begin
          reg148 <= reg151[(1'h1):(1'h1)];
        end
      for (forvar165 = (1'h0); (forvar165 < (2'h2)); forvar165 = (forvar165 + (1'h1)))
        begin
          if ({wire142[(3'h4):(2'h3)]})
            begin
              reg166 = (-forvar165[(4'h9):(3'h5)]);
              reg167 <= {((^~wire145) + ($signed((wire147 >= reg130)) ?
                      {reg150[(4'h8):(3'h6)],
                          (^wire144)} : $signed({reg148})))};
              reg168 = (-($signed($signed($unsigned(wire138))) >> reg156));
              reg169 = reg157;
              reg170 = ($unsigned(wire139[(3'h4):(3'h4)]) ?
                  reg166 : $unsigned({$unsigned($signed((8'ha0)))}));
            end
          else
            begin
              reg166 = (((^~(^~wire113)) ?
                      $unsigned((reg161[(1'h1):(1'h0)] ?
                          $unsigned(reg153) : (reg158 ^~ wire113))) : {reg152[(3'h7):(2'h2)],
                          (8'ha4)}) ?
                  {$unsigned((!(8'ha8))),
                      (-reg158[(2'h2):(1'h0)])} : reg150[(2'h3):(2'h2)]);
            end
        end
      if ({(($unsigned($unsigned(wire145)) < ((reg159 | wire110) ?
                  wire135[(1'h0):(1'h0)] : $signed((8'ha1)))) ?
              reg166[(3'h4):(2'h3)] : reg151)})
        begin
          reg171 <= $signed(($signed(((wire138 ?
                  reg120 : wire138) < $signed(reg166))) ?
              (((reg124 ? forvar160 : reg168) ~^ reg151) ?
                  reg159 : $unsigned($unsigned(reg163))) : $signed(reg159[(1'h1):(1'h0)])));
        end
      else
        begin
          if (($unsigned(reg148[(4'hd):(3'h6)]) ? reg167 : wire143))
            begin
              reg172 = reg149[(1'h0):(1'h0)];
              reg173 <= $unsigned((+$unsigned($signed({wire138}))));
              reg174 <= reg161[(1'h1):(1'h1)];
            end
          else
            begin
              reg172 = (reg118 ? reg170[(3'h7):(2'h3)] : $signed((8'hae)));
              reg173 <= ((((+(wire146 ? wire144 : reg156)) << (~&(!(8'hbd)))) ?
                  reg120[(2'h3):(1'h0)] : {(^$signed(wire140))}) - (!(!{$signed(reg153),
                  $signed(reg151)})));
              reg174 <= $signed((8'ha9));
            end
          if ($signed($unsigned($unsigned((~^$signed((8'hb1)))))))
            begin
              reg175 <= $unsigned(((($unsigned(reg171) != (!wire141)) << (8'ha7)) ^ $unsigned(reg120[(3'h5):(1'h1)])));
              reg176 = (8'ha1);
              reg177 = wire144[(4'hb):(3'h5)];
            end
          else
            begin
              reg175 <= wire145[(2'h2):(1'h0)];
              reg176 = (((&{reg164[(1'h1):(1'h0)]}) ?
                      reg171[(4'he):(4'hc)] : (+reg148[(2'h3):(1'h0)])) ?
                  (~^{$signed((~&reg150))}) : (!forvar165));
              reg177 = reg157;
              reg178 = $signed((~|wire145));
            end
          if ((reg115[(2'h2):(1'h0)] | ($signed(wire139[(1'h0):(1'h0)]) ?
              $signed((^reg176[(4'hb):(3'h6)])) : $unsigned({$unsigned((8'haf)),
                  reg124[(4'ha):(2'h2)]}))))
            begin
              reg179 <= wire134;
              reg180 = wire111[(2'h2):(1'h0)];
              reg181 = ((~|$signed((^~$unsigned(wire134)))) ?
                  $unsigned(reg153[(3'h5):(3'h5)]) : {((&$unsigned(reg177)) ?
                          reg118[(4'h8):(3'h6)] : $signed(wire142)),
                      $signed($signed((|reg172)))});
            end
          else
            begin
              reg179 <= (((reg150[(4'hd):(4'ha)] & ($signed(reg176) || (~&(8'ha9)))) ?
                  $unsigned($unsigned(wire109)) : $signed({{wire111}})) >= reg179);
              reg182 <= $unsigned(reg181);
              reg183 <= ({(+$signed((~^wire146))),
                  (&{((8'hbe) ?
                          (8'ha1) : wire109)})} << $signed(((~&$signed(wire139)) <<< (-reg118))));
              reg184 = $signed($signed((~^($signed(reg148) ?
                  reg167[(4'h9):(3'h5)] : $unsigned((8'ha0))))));
            end
          reg185 <= (~^$unsigned((~(((8'haf) ?
              wire134 : reg158) >>> $unsigned(wire145)))));
          reg186 <= (wire112 || {wire141, (~&(+(reg183 ~^ reg118)))});
        end
    end
  assign wire187 = $signed(reg150[(3'h5):(2'h3)]);
  assign wire188 = (+({($unsigned(wire135) ? {reg157} : (reg182 > reg128))} ?
                       {wire137,
                           $signed((reg161 * reg126))} : $unsigned(((~&reg179) <<< {(8'ha3)}))));
  assign wire189 = $unsigned({(((!wire138) ?
                               reg173[(2'h2):(1'h1)] : (reg175 <<< reg163)) ?
                           {wire137[(1'h1):(1'h1)],
                               (8'ha2)} : wire147[(1'h1):(1'h1)]),
                       $signed((((8'hba) && reg183) ?
                           (^~reg183) : wire134[(3'h4):(1'h1)]))});
  assign wire190 = reg115[(5'h12):(4'hb)];
  assign wire191 = (wire109[(1'h0):(1'h0)] ?
                       ((($unsigned(reg128) ^~ {reg183, reg118}) ?
                               $unsigned((~&reg150)) : ($signed(wire137) * $signed(wire146))) ?
                           $unsigned(wire143[(2'h2):(1'h0)]) : (~|($signed(reg186) ~^ (^~reg183)))) : ((wire134[(4'hb):(4'h8)] ?
                           ((wire140 ?
                               wire112 : (8'h9d)) <<< (wire110 != wire135)) : $unsigned({reg186,
                               wire110})) && (!$signed((reg150 <<< reg115)))));
  assign wire192 = ($unsigned($signed(reg155[(1'h0):(1'h0)])) + reg185);
  always
    @(posedge clk) begin
      reg193 = $signed((&$signed(wire190)));
      reg194 = (reg175 & (~&reg171));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module82  (y, clk, wire86, wire85, wire84, wire83);
  output wire [(32'hed):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire86;
  input wire signed [(2'h3):(1'h0)] wire85;
  input wire [(4'hc):(1'h0)] wire84;
  input wire [(5'h11):(1'h0)] wire83;
  wire [(4'hd):(1'h0)] wire103;
  wire signed [(4'ha):(1'h0)] wire102;
  wire signed [(5'h10):(1'h0)] wire101;
  wire [(4'hd):(1'h0)] wire100;
  wire [(5'h15):(1'h0)] wire99;
  wire [(4'hf):(1'h0)] wire98;
  wire [(3'h7):(1'h0)] wire97;
  wire [(4'hc):(1'h0)] wire96;
  wire [(5'h13):(1'h0)] wire89;
  wire [(5'h14):(1'h0)] wire88;
  wire [(4'h9):(1'h0)] wire87;
  reg [(5'h11):(1'h0)] reg94 = (1'h0);
  reg [(5'h15):(1'h0)] reg93 = (1'h0);
  reg [(4'ha):(1'h0)] reg91 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg95 = (1'h0);
  reg [(3'h6):(1'h0)] reg92 = (1'h0);
  reg [(4'hf):(1'h0)] reg90 = (1'h0);
  assign y = {wire103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 wire97,
                 wire96,
                 wire89,
                 wire88,
                 wire87,
                 reg94,
                 reg93,
                 reg91,
                 reg95,
                 reg92,
                 reg90,
                 (1'h0)};
  assign wire87 = wire84[(4'hc):(3'h7)];
  assign wire88 = {($signed($unsigned(wire86)) ?
                          {$signed((wire86 <<< (8'hb3)))} : wire86[(1'h0):(1'h0)]),
                      wire85};
  assign wire89 = $unsigned(((~{wire84}) ^ ((~((8'ha3) + wire83)) & $unsigned({wire88}))));
  always
    @(posedge clk) begin
      if (wire85)
        begin
          reg90 = $unsigned(wire84[(3'h7):(3'h4)]);
        end
      else
        begin
          if ($unsigned(wire83))
            begin
              reg90 = ({$signed(({wire84} >> (reg90 ?
                      (8'ha8) : wire88)))} & (((&$unsigned((8'ha4))) - $signed($signed(reg90))) == ((|$unsigned(reg90)) >> ((~&(7'h41)) ?
                  (|wire86) : {reg90, reg90}))));
            end
          else
            begin
              reg91 <= $unsigned(wire84[(1'h0):(1'h0)]);
              reg92 = ($signed((~($unsigned((8'hb8)) ?
                      (8'h9e) : $unsigned(wire87)))) ?
                  wire84 : (~&(wire83[(5'h11):(4'he)] ?
                      ((reg90 >>> wire83) ?
                          wire88 : $unsigned(reg90)) : (wire89[(5'h11):(2'h3)] ^ (+(8'hb2))))));
              reg93 <= ($signed((($signed(wire83) << (^wire84)) ?
                      (~&wire84) : wire85[(2'h2):(2'h2)])) ?
                  (^~reg90) : reg90[(4'hd):(4'h9)]);
              reg94 <= $unsigned($unsigned($signed({{reg91, wire87}})));
              reg95 = (wire89 >> reg94[(5'h10):(3'h4)]);
            end
        end
    end
  assign wire96 = $signed($unsigned(((^reg91) ?
                      (wire89 ? wire86 : reg91[(2'h2):(1'h1)]) : wire89)));
  assign wire97 = $signed(wire96);
  assign wire98 = $signed(($unsigned(wire88) < reg91));
  assign wire99 = reg91;
  assign wire100 = (8'hb3);
  assign wire101 = (($unsigned((~$signed(wire100))) ?
                       {$unsigned(reg93)} : {$signed((reg93 >> (8'ha6)))}) << {(&$unsigned(((8'ha7) ?
                           wire100 : wire86)))});
  assign wire102 = ($signed((!wire88[(4'h8):(3'h4)])) >>> {reg94[(4'hb):(4'h9)],
                       ($signed((wire101 ? reg91 : reg94)) - (|wire85))});
  assign wire103 = $signed(($unsigned((8'ha7)) <= $unsigned(((wire85 ?
                       wire83 : reg91) < (reg94 <= wire98)))));
endmodule