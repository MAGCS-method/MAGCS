(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param265 = {{(^((|(8'h9e)) ? ((8'hb3) ? (7'h43) : (8'ha2)) : (^(8'hb2)))), {(8'h9f)}}, ((-(^~(^~(8'ha7)))) * (~&(!(^(8'ha2)))))}, 
parameter param266 = (((~&((param265 ? param265 : (8'h9d)) <<< (^param265))) ? (8'hba) : (&({param265, param265} ? (param265 ? param265 : param265) : (param265 >>> (8'h9d))))) + ((8'hbb) ? {(((8'ha2) && (8'ha0)) ? (param265 || param265) : param265), param265} : {((!param265) - {param265, param265})})))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h285):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire0;
  input wire signed [(4'hb):(1'h0)] wire1;
  input wire signed [(4'ha):(1'h0)] wire2;
  input wire [(5'h10):(1'h0)] wire3;
  wire signed [(5'h10):(1'h0)] wire264;
  wire signed [(3'h5):(1'h0)] wire262;
  wire signed [(5'h15):(1'h0)] wire244;
  wire signed [(5'h14):(1'h0)] wire243;
  wire signed [(4'hb):(1'h0)] wire242;
  wire signed [(5'h14):(1'h0)] wire240;
  wire signed [(2'h2):(1'h0)] wire239;
  wire [(5'h13):(1'h0)] wire238;
  wire signed [(3'h7):(1'h0)] wire236;
  reg [(5'h14):(1'h0)] reg6 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7 = (1'h0);
  reg [(4'hd):(1'h0)] reg8 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg9 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg11 = (1'h0);
  reg [(4'hc):(1'h0)] reg12 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg15 = (1'h0);
  reg [(5'h14):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg17 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg18 = (1'h0);
  reg [(3'h5):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg20 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg21 = (1'h0);
  reg [(5'h11):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg23 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg246 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg247 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg249 = (1'h0);
  reg [(4'ha):(1'h0)] reg251 = (1'h0);
  reg [(3'h6):(1'h0)] reg253 = (1'h0);
  reg [(4'ha):(1'h0)] reg245 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg255 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg258 = (1'h0);
  reg [(2'h3):(1'h0)] reg259 = (1'h0);
  reg [(5'h13):(1'h0)] reg260 = (1'h0);
  reg [(5'h12):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg256 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg254 = (1'h0);
  reg [(4'ha):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg250 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar245 = (1'h0);
  reg [(5'h12):(1'h0)] forvar19 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg14 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar10 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar4 = (1'h0);
  assign y = {wire264,
                 wire262,
                 wire244,
                 wire243,
                 wire242,
                 wire240,
                 wire239,
                 wire238,
                 wire236,
                 reg6,
                 reg7,
                 reg8,
                 reg9,
                 reg11,
                 reg12,
                 reg13,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg241,
                 reg246,
                 reg247,
                 reg248,
                 reg249,
                 reg251,
                 reg253,
                 reg245,
                 reg255,
                 reg258,
                 reg259,
                 reg260,
                 reg261,
                 reg257,
                 reg256,
                 reg254,
                 reg252,
                 reg250,
                 forvar245,
                 forvar19,
                 reg14,
                 forvar10,
                 forvar5,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (2'h3)); forvar4 = (forvar4 + (1'h1)))
        begin
          for (forvar5 = (1'h0); (forvar5 < (3'h4)); forvar5 = (forvar5 + (1'h1)))
            begin
              reg6 <= $unsigned(wire1);
              reg7 <= ($unsigned({$unsigned((wire2 ? forvar5 : wire2))}) ?
                  $unsigned(wire2) : $unsigned(forvar5));
            end
          reg8 <= ((|$unsigned($unsigned(forvar4))) ?
              (|$signed((wire1[(1'h1):(1'h1)] ?
                  forvar5[(1'h1):(1'h1)] : (reg6 & wire1)))) : $unsigned(wire0[(1'h1):(1'h1)]));
          reg9 <= $unsigned((wire0 ?
              ($signed(forvar5) < ($unsigned((8'ha6)) ^~ wire0)) : (!((reg7 ?
                      reg6 : reg7) ?
                  (^wire3) : {forvar5, wire3}))));
          for (forvar10 = (1'h0); (forvar10 < (1'h1)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg11 <= $unsigned(forvar4[(5'h15):(5'h10)]);
              reg12 <= reg9[(2'h3):(2'h3)];
              reg13 <= (((~{$signed((8'hb7)),
                      (wire3 ? forvar4 : wire1)}) && (~(wire0 ?
                      (reg11 ? reg12 : reg9) : (reg6 ? forvar5 : reg12)))) ?
                  ($signed(wire2) ^ forvar10[(1'h0):(1'h0)]) : (^~$unsigned($signed({wire3,
                      forvar10}))));
            end
          reg14 = (~|(~|$unsigned((&wire1[(2'h2):(1'h1)]))));
        end
      reg15 <= $signed(wire3);
    end
  always
    @(posedge clk) begin
      reg16 <= $signed((^~reg6[(4'hb):(3'h4)]));
      reg17 <= ($signed($unsigned($unsigned((|(8'hb8))))) && (($unsigned((reg6 << (7'h40))) ?
          reg16[(1'h1):(1'h1)] : $unsigned({reg13})) ~^ wire2));
      if ($unsigned(((((reg13 * reg6) || reg13[(1'h0):(1'h0)]) & $unsigned((reg12 <<< wire3))) >>> reg13[(2'h2):(1'h1)])))
        begin
          reg18 <= $signed(((wire3[(4'ha):(3'h7)] ?
                  (^reg16) : (^~(reg13 != wire1))) ?
              {wire3} : (~|{$unsigned(reg15)})));
          reg19 <= reg18[(4'hb):(3'h7)];
          reg20 <= $signed(reg6[(3'h7):(3'h4)]);
          reg21 <= ($signed(((!$unsigned(wire1)) - $signed(reg20))) ?
              $unsigned(reg17[(3'h7):(3'h6)]) : ((~&reg13[(1'h0):(1'h0)]) ?
                  {(~(wire3 ? reg19 : reg8)),
                      ((|wire0) ?
                          {reg13,
                              reg18} : reg19)} : (reg16[(1'h1):(1'h0)] ^ ($unsigned(reg20) ?
                      (~|reg16) : (reg7 < reg8)))));
        end
      else
        begin
          reg18 <= (reg6 + ($signed(($signed(reg7) & $signed(wire1))) ?
              ((((8'haf) ? reg17 : reg6) ?
                  $unsigned((8'hb9)) : (wire2 ?
                      reg13 : reg8)) ^~ wire3) : reg11));
          for (forvar19 = (1'h0); (forvar19 < (2'h3)); forvar19 = (forvar19 + (1'h1)))
            begin
              reg20 <= {(reg7 ? wire1[(2'h2):(2'h2)] : reg20),
                  $unsigned(forvar19)};
            end
        end
      reg22 <= $unsigned($signed($unsigned(reg20)));
      reg23 <= reg16[(1'h1):(1'h0)];
    end
  module24 #() modinst237 (.wire27(reg6), .wire26(wire0), .y(wire236), .wire29(reg17), .clk(clk), .wire25(reg16), .wire28(reg9));
  assign wire238 = reg11[(5'h11):(4'hb)];
  assign wire239 = ($signed(wire3) ?
                       ($unsigned($signed((reg15 ?
                           reg22 : (8'ha2)))) >= reg20) : {reg22});
  assign wire240 = $signed((reg15 != (-($unsigned(reg7) ?
                       reg6[(4'ha):(2'h3)] : $signed(reg17)))));
  always
    @(posedge clk) begin
      reg241 <= reg7[(3'h4):(2'h2)];
    end
  assign wire242 = (-$unsigned(wire239));
  assign wire243 = ($unsigned($signed(((reg7 | reg9) & (~(8'haf))))) + reg16[(5'h13):(3'h4)]);
  assign wire244 = $signed(reg6);
  always
    @(posedge clk) begin
      if ((wire236[(3'h6):(2'h3)] ?
          ((wire2 ?
                  ({reg12, wire236} ?
                      reg9 : (reg20 ?
                          reg19 : wire240)) : wire1[(4'h8):(1'h0)]) ?
              (8'hbb) : (^~((+wire2) ^ $signed(wire239)))) : (~&$signed($signed(wire2[(2'h2):(1'h0)])))))
        begin
          for (forvar245 = (1'h0); (forvar245 < (1'h1)); forvar245 = (forvar245 + (1'h1)))
            begin
              reg246 <= ($signed($unsigned(((~^wire243) ?
                  reg15[(4'hd):(4'hc)] : $signed((8'hb2))))) >= ((({reg6} ?
                          reg16[(5'h14):(4'hc)] : wire239) ?
                      (^$unsigned(wire242)) : $unsigned((reg9 ?
                          wire242 : wire238))) ?
                  (~^reg6) : {wire238}));
              reg247 <= $unsigned((^~$signed(((|(8'hb0)) ?
                  $signed(reg7) : reg20[(5'h10):(2'h2)]))));
              reg248 <= {$unsigned((!((reg17 ? (8'ha8) : wire243) ?
                      $unsigned(reg12) : {wire2, reg15}))),
                  (reg6 ?
                      (8'hbe) : (((~^wire1) ?
                              reg247[(3'h5):(2'h3)] : reg15[(4'h9):(3'h7)]) ?
                          ($unsigned(wire3) ?
                              wire1[(3'h5):(1'h0)] : $signed(reg7)) : (((8'ha8) >= (8'ha8)) != $signed(wire238))))};
              reg249 <= (~reg23[(2'h2):(1'h0)]);
              reg250 = {reg20,
                  (wire236 ? $signed(reg246[(4'h9):(1'h0)]) : {reg15})};
            end
          reg251 <= wire0;
          reg252 = {(reg246 ?
                  $signed(reg248[(3'h5):(1'h1)]) : reg23[(2'h2):(1'h1)])};
          reg253 <= (~|((~^(!$unsigned(wire243))) ? (8'hba) : wire242));
          reg254 = $unsigned($unsigned(reg7));
        end
      else
        begin
          reg245 <= (({reg12[(1'h1):(1'h1)],
              $signed((reg22 ? wire236 : reg18))} ~^ ((~&(&(8'hbf))) ?
              reg20 : (reg250[(3'h4):(1'h1)] ?
                  $signed(reg12) : {wire239,
                      reg18}))) + (($unsigned(reg17[(5'h12):(4'hc)]) && {$signed(forvar245),
              (^wire0)}) || wire1[(4'hb):(3'h7)]));
          reg246 <= (($unsigned($signed(wire240[(2'h2):(1'h1)])) ?
              reg16 : reg247[(1'h0):(1'h0)]) >> $signed((^~wire239)));
          reg250 = wire3;
          reg251 <= reg15;
        end
      reg255 <= $unsigned($signed($signed((8'hb5))));
      reg256 = (8'hbe);
      if ((reg19[(2'h3):(1'h1)] ? (8'hac) : (|(^reg20))))
        begin
          reg257 = {reg252[(2'h2):(1'h1)],
              (~((^~$signed(reg13)) ?
                  $unsigned(((8'ha1) ? wire240 : (8'ha1))) : (~wire243)))};
          reg258 <= wire3[(2'h2):(1'h1)];
          reg259 <= (($unsigned(reg250) ?
              reg11[(3'h7):(3'h5)] : (!(reg241[(2'h3):(1'h0)] == (reg7 * (8'hb5))))) >> ((~|((reg257 ?
                      reg13 : reg20) ?
                  $unsigned(reg22) : reg241)) ?
              ($unsigned((wire242 ? reg248 : reg23)) * {wire239[(2'h2):(1'h1)],
                  reg246[(2'h2):(1'h0)]}) : $unsigned((^~{reg7, wire2}))));
          reg260 <= {reg12, reg245};
          reg261 <= ($signed(wire0[(2'h2):(1'h0)]) << ((!(~&(wire239 * reg252))) <= (reg248[(3'h4):(1'h1)] ?
              reg245 : $signed(wire244))));
        end
      else
        begin
          reg258 <= $unsigned(reg11[(5'h10):(1'h0)]);
          reg259 <= (~&$unsigned(((~&$signed(reg256)) ?
              (forvar245[(2'h2):(2'h2)] >= reg251) : $unsigned({(8'hba),
                  reg11}))));
        end
    end
  module24 #() modinst263 (.wire28(reg16), .wire29(wire0), .y(wire262), .wire26(reg23), .clk(clk), .wire25(wire240), .wire27(reg249));
  assign wire264 = reg258;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module24
#(parameter param235 = ((~|{((^(8'ha9)) ? ((8'ha5) ? (8'hbf) : (8'hb3)) : ((8'hb4) >= (7'h42))), (^((8'hac) ~^ (8'ha8)))}) | ({(((8'hbb) ? (8'ha1) : (8'ha6)) >= ((8'hb4) == (8'hbe)))} | ({(-(8'hb4))} + ({(8'ha6), (8'hba)} ? (~|(8'hbe)) : ((8'hb9) != (8'haf)))))))
(y, clk, wire25, wire26, wire27, wire28, wire29);
  output wire [(32'h196):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire25;
  input wire [(5'h15):(1'h0)] wire26;
  input wire [(5'h14):(1'h0)] wire27;
  input wire signed [(4'h9):(1'h0)] wire28;
  input wire signed [(5'h14):(1'h0)] wire29;
  wire signed [(2'h3):(1'h0)] wire234;
  wire signed [(4'he):(1'h0)] wire233;
  wire [(4'he):(1'h0)] wire227;
  wire [(3'h4):(1'h0)] wire226;
  wire [(4'h9):(1'h0)] wire225;
  wire signed [(4'hc):(1'h0)] wire224;
  wire signed [(5'h15):(1'h0)] wire223;
  wire [(4'hb):(1'h0)] wire221;
  wire signed [(4'hf):(1'h0)] wire172;
  wire signed [(5'h11):(1'h0)] wire171;
  wire [(5'h14):(1'h0)] wire170;
  wire [(5'h14):(1'h0)] wire169;
  wire [(4'he):(1'h0)] wire155;
  wire [(2'h3):(1'h0)] wire153;
  wire signed [(5'h12):(1'h0)] wire119;
  wire [(5'h11):(1'h0)] wire118;
  wire [(5'h13):(1'h0)] wire116;
  wire [(4'hb):(1'h0)] wire51;
  reg signed [(4'hd):(1'h0)] reg232 = (1'h0);
  reg signed [(4'he):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg229 = (1'h0);
  reg [(2'h3):(1'h0)] reg228 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg166 = (1'h0);
  reg [(3'h4):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg164 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg161 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg159 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg157 = (1'h0);
  reg [(2'h2):(1'h0)] reg156 = (1'h0);
  reg [(2'h2):(1'h0)] reg231 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg168 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar163 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg160 = (1'h0);
  reg [(4'he):(1'h0)] forvar158 = (1'h0);
  assign y = {wire234,
                 wire233,
                 wire227,
                 wire226,
                 wire225,
                 wire224,
                 wire223,
                 wire221,
                 wire172,
                 wire171,
                 wire170,
                 wire169,
                 wire155,
                 wire153,
                 wire119,
                 wire118,
                 wire116,
                 wire51,
                 reg232,
                 reg230,
                 reg229,
                 reg228,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg162,
                 reg161,
                 reg159,
                 reg157,
                 reg156,
                 reg231,
                 reg168,
                 forvar163,
                 reg160,
                 forvar158,
                 (1'h0)};
  assign wire118 = wire51[(2'h3):(1'h0)];
  assign wire119 = wire28[(1'h1):(1'h0)];
  assign wire155 = wire26[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg156 <= (wire29[(4'h8):(3'h7)] ?
          $signed(wire51[(2'h3):(1'h1)]) : wire26[(2'h2):(2'h2)]);
      reg157 <= $unsigned($signed(wire25[(4'hb):(4'h8)]));
      for (forvar158 = (1'h0); (forvar158 < (1'h0)); forvar158 = (forvar158 + (1'h1)))
        begin
          reg159 <= wire27[(5'h14):(3'h4)];
          reg160 = wire27;
          reg161 <= (($unsigned({(wire25 ? reg157 : wire155),
                  $signed(wire153)}) ^ wire28[(4'h8):(2'h3)]) ?
              (wire116 ?
                  ($signed({wire26, wire29}) ?
                      $signed(reg160[(1'h0):(1'h0)]) : ($signed(wire25) ?
                          wire28[(4'h8):(1'h1)] : (&wire155))) : forvar158[(1'h1):(1'h1)]) : reg159[(1'h0):(1'h0)]);
          reg162 <= wire27;
          for (forvar163 = (1'h0); (forvar163 < (2'h3)); forvar163 = (forvar163 + (1'h1)))
            begin
              reg164 <= ((-($signed($signed(wire51)) <<< forvar163)) && $signed((forvar163 ?
                  (8'hac) : $unsigned(wire27))));
              reg165 <= ($signed((wire116[(2'h3):(1'h1)] >>> wire51)) ^ ((^~(~^reg161[(3'h7):(1'h0)])) ?
                  (!(((8'hac) ?
                      wire153 : reg160) << $unsigned(forvar163))) : (((~|(8'hb8)) ~^ $unsigned(reg161)) <<< wire28[(2'h2):(1'h1)])));
              reg166 <= wire153[(1'h0):(1'h0)];
              reg167 <= wire153[(1'h0):(1'h0)];
            end
        end
      reg168 = wire28[(1'h0):(1'h0)];
    end
  assign wire169 = $signed((^~($signed(wire155) < $signed((wire25 ?
                       (7'h41) : wire116)))));
  assign wire170 = wire29[(5'h10):(4'he)];
  assign wire171 = wire169;
  assign wire172 = (({wire153[(2'h2):(1'h0)]} ?
                           $unsigned(reg166[(1'h0):(1'h0)]) : reg164[(5'h11):(4'hc)]) ?
                       reg165 : $signed(wire153[(2'h2):(2'h2)]));
  assign wire223 = {wire172[(3'h6):(1'h0)]};
  assign wire224 = $signed(wire223);
  assign wire225 = wire27;
  assign wire226 = ({wire153, wire223} > wire51[(2'h3):(1'h1)]);
  assign wire227 = (($signed(wire118) ?
                       $unsigned({$signed((8'h9e))}) : {(8'ha7),
                           ((reg157 ? wire224 : reg161) ?
                               $unsigned(wire29) : {reg162})}) * ($unsigned(wire225) & reg167));
  always
    @(posedge clk) begin
      reg228 <= wire51[(3'h6):(3'h4)];
      reg229 <= $signed({wire119[(4'hd):(3'h7)], wire226[(1'h0):(1'h0)]});
      reg230 <= reg162[(1'h0):(1'h0)];
      reg231 = ((({(wire26 ? wire29 : wire172), (wire172 | wire29)} ?
              reg166 : ({wire223, wire155} ^~ wire118[(4'ha):(2'h2)])) ?
          wire26[(3'h6):(3'h6)] : {{reg229[(5'h13):(4'hf)],
                  $signed(wire170)}}) != (+(((reg228 & wire26) ^ $signed(wire227)) | (&(reg157 & wire223)))));
      reg232 <= $signed(wire171[(5'h11):(4'hf)]);
    end
  assign wire233 = $signed(wire223[(3'h7):(2'h2)]);
  assign wire234 = wire233;
endmodule
