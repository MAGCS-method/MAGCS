(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param3358 = ((8'h9f) || {{((!(8'hae)) << ((8'hb2) >>> (8'hb2)))}}))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h13eb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h1a):(1'h0)] wire0;
  input wire signed [(5'h13):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire2;
  input wire [(5'h18):(1'h0)] wire3;
  wire signed [(4'h9):(1'h0)] wire3216;
  wire [(5'h1b):(1'h0)] wire3211;
  wire [(5'h17):(1'h0)] wire3210;
  wire signed [(4'hf):(1'h0)] wire3209;
  wire [(3'h7):(1'h0)] wire3198;
  wire [(5'h1b):(1'h0)] wire3197;
  wire [(3'h5):(1'h0)] wire3196;
  wire [(5'h1a):(1'h0)] wire3076;
  wire signed [(4'he):(1'h0)] wire4;
  wire [(5'h13):(1'h0)] wire5;
  wire [(5'h15):(1'h0)] wire3071;
  wire [(5'h13):(1'h0)] wire3073;
  wire signed [(5'h18):(1'h0)] wire3074;
  wire [(5'h16):(1'h0)] wire3078;
  wire [(5'h1b):(1'h0)] wire3079;
  wire [(5'h13):(1'h0)] wire3105;
  wire [(5'h1f):(1'h0)] wire3193;
  wire [(4'he):(1'h0)] wire3194;
  wire [(5'h19):(1'h0)] wire3218;
  wire signed [(4'hc):(1'h0)] wire3219;
  wire signed [(5'h14):(1'h0)] wire3353;
  wire signed [(4'h8):(1'h0)] wire3356;
  reg signed [(5'h18):(1'h0)] reg3080 = (1'h0);
  reg [(5'h15):(1'h0)] reg3081 = (1'h0);
  reg [(5'h12):(1'h0)] reg3085 = (1'h0);
  reg [(3'h7):(1'h0)] reg3087 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3090 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3091 = (1'h0);
  reg [(4'h8):(1'h0)] reg3094 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3095 = (1'h0);
  reg [(5'h14):(1'h0)] reg3099 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3100 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3101 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3103 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3104 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3108 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3109 = (1'h0);
  reg [(2'h3):(1'h0)] reg3110 = (1'h0);
  reg [(4'ha):(1'h0)] reg3115 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3119 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3122 = (1'h0);
  reg [(3'h4):(1'h0)] reg3126 = (1'h0);
  reg [(5'h16):(1'h0)] reg3128 = (1'h0);
  reg [(5'h13):(1'h0)] reg3129 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3131 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3133 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3134 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3135 = (1'h0);
  reg [(5'h15):(1'h0)] reg3136 = (1'h0);
  reg [(4'hc):(1'h0)] reg3140 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3141 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3142 = (1'h0);
  reg [(4'h8):(1'h0)] reg3144 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3146 = (1'h0);
  reg [(5'h10):(1'h0)] reg3148 = (1'h0);
  reg [(3'h4):(1'h0)] reg3149 = (1'h0);
  reg [(3'h6):(1'h0)] reg3150 = (1'h0);
  reg [(4'hc):(1'h0)] reg3151 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3153 = (1'h0);
  reg [(4'ha):(1'h0)] reg3155 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3156 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3157 = (1'h0);
  reg [(5'h13):(1'h0)] reg3162 = (1'h0);
  reg [(4'hf):(1'h0)] reg3163 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3165 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3167 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3168 = (1'h0);
  reg [(4'hb):(1'h0)] reg3170 = (1'h0);
  reg [(4'hb):(1'h0)] reg3171 = (1'h0);
  reg [(5'h11):(1'h0)] reg3173 = (1'h0);
  reg [(5'h13):(1'h0)] reg3176 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3177 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3179 = (1'h0);
  reg [(4'hf):(1'h0)] reg3181 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3183 = (1'h0);
  reg [(5'h13):(1'h0)] reg3184 = (1'h0);
  reg [(5'h11):(1'h0)] reg3186 = (1'h0);
  reg [(4'hb):(1'h0)] reg3188 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3191 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3203 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3204 = (1'h0);
  reg [(5'h15):(1'h0)] reg3206 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3207 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3208 = (1'h0);
  reg [(5'h10):(1'h0)] reg3212 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3213 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3224 = (1'h0);
  reg [(3'h7):(1'h0)] reg3225 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3229 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3231 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3232 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3234 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3237 = (1'h0);
  reg [(3'h4):(1'h0)] reg3243 = (1'h0);
  reg [(4'hf):(1'h0)] reg3244 = (1'h0);
  reg [(4'hc):(1'h0)] reg3246 = (1'h0);
  reg [(5'h13):(1'h0)] reg3247 = (1'h0);
  reg [(4'hb):(1'h0)] reg3249 = (1'h0);
  reg [(5'h16):(1'h0)] reg3250 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3257 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3259 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3264 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3265 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3266 = (1'h0);
  reg [(2'h3):(1'h0)] reg3268 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3269 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3272 = (1'h0);
  reg [(4'hc):(1'h0)] reg3275 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3277 = (1'h0);
  reg [(5'h13):(1'h0)] reg3280 = (1'h0);
  reg [(5'h11):(1'h0)] reg3282 = (1'h0);
  reg [(5'h14):(1'h0)] reg3283 = (1'h0);
  reg [(2'h3):(1'h0)] reg3284 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3286 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3289 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3290 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3291 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3292 = (1'h0);
  reg [(5'h10):(1'h0)] reg3295 = (1'h0);
  reg [(5'h16):(1'h0)] reg3296 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3297 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3299 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3300 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3301 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3302 = (1'h0);
  reg [(5'h10):(1'h0)] reg3303 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3305 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3308 = (1'h0);
  reg [(3'h7):(1'h0)] reg3312 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3313 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3315 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3316 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3319 = (1'h0);
  reg [(5'h18):(1'h0)] reg3323 = (1'h0);
  reg [(3'h7):(1'h0)] reg3325 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3328 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3332 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3321 = (1'h0);
  reg [(4'hf):(1'h0)] reg3334 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3335 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3338 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3340 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3341 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3342 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3343 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3345 = (1'h0);
  reg [(5'h13):(1'h0)] reg3346 = (1'h0);
  reg [(4'hc):(1'h0)] reg3349 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3352 = (1'h0);
  reg [(5'h15):(1'h0)] reg3355 = (1'h0);
  reg [(5'h13):(1'h0)] reg3351 = (1'h0);
  reg [(4'hc):(1'h0)] reg3350 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3348 = (1'h0);
  reg [(4'h8):(1'h0)] reg3347 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3344 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3339 = (1'h0);
  reg [(5'h19):(1'h0)] reg3337 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3336 = (1'h0);
  reg [(5'h16):(1'h0)] reg3333 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar3330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3326 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3318 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3331 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3330 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3329 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3327 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3326 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3324 = (1'h0);
  reg [(5'h16):(1'h0)] reg3322 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3321 = (1'h0);
  reg [(5'h13):(1'h0)] reg3320 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3318 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3317 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3314 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3311 = (1'h0);
  reg [(4'he):(1'h0)] reg3310 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3309 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3307 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3306 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3304 = (1'h0);
  reg [(3'h5):(1'h0)] reg3298 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3296 = (1'h0);
  reg [(4'h9):(1'h0)] reg3293 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3294 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3293 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3288 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3287 = (1'h0);
  reg [(4'hc):(1'h0)] reg3285 = (1'h0);
  reg [(5'h19):(1'h0)] reg3276 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3281 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3279 = (1'h0);
  reg [(2'h2):(1'h0)] reg3278 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3276 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3273 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3269 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3274 = (1'h0);
  reg [(5'h13):(1'h0)] forvar3273 = (1'h0);
  reg [(5'h19):(1'h0)] reg3271 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3270 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3267 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3263 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3262 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3261 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3260 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3258 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3256 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3255 = (1'h0);
  reg [(4'he):(1'h0)] reg3254 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3253 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3252 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3251 = (1'h0);
  reg [(5'h16):(1'h0)] reg3248 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3245 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3242 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3241 = (1'h0);
  reg [(2'h3):(1'h0)] reg3240 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3239 = (1'h0);
  reg [(4'hd):(1'h0)] reg3238 = (1'h0);
  reg [(5'h14):(1'h0)] reg3236 = (1'h0);
  reg [(2'h3):(1'h0)] reg3235 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3233 = (1'h0);
  reg [(5'h10):(1'h0)] reg3230 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3228 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3227 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3226 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3223 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3222 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar3221 = (1'h0);
  reg [(5'h16):(1'h0)] forvar3220 = (1'h0);
  reg [(4'h8):(1'h0)] reg3215 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3214 = (1'h0);
  reg [(3'h4):(1'h0)] reg3205 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3202 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar3201 = (1'h0);
  reg [(5'h18):(1'h0)] forvar3200 = (1'h0);
  reg [(4'h8):(1'h0)] reg3192 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3190 = (1'h0);
  reg [(3'h7):(1'h0)] reg3189 = (1'h0);
  reg [(4'hf):(1'h0)] reg3187 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar3185 = (1'h0);
  reg [(3'h7):(1'h0)] reg3182 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3180 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3178 = (1'h0);
  reg [(5'h10):(1'h0)] reg3175 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3174 = (1'h0);
  reg [(5'h17):(1'h0)] reg3172 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3169 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3166 = (1'h0);
  reg [(5'h19):(1'h0)] reg3159 = (1'h0);
  reg [(4'hf):(1'h0)] reg3152 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3149 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3145 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3139 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar3131 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3164 = (1'h0);
  reg [(4'h8):(1'h0)] reg3161 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3160 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3159 = (1'h0);
  reg [(4'hd):(1'h0)] reg3158 = (1'h0);
  reg [(4'hb):(1'h0)] reg3154 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar3152 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3147 = (1'h0);
  reg [(5'h16):(1'h0)] forvar3145 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3143 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3139 = (1'h0);
  reg [(5'h17):(1'h0)] reg3138 = (1'h0);
  reg [(4'hf):(1'h0)] reg3137 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3132 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3130 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3127 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3125 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3124 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3123 = (1'h0);
  reg [(5'h18):(1'h0)] reg3121 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3120 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3118 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar3117 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3116 = (1'h0);
  reg [(2'h3):(1'h0)] reg3114 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3113 = (1'h0);
  reg [(4'hb):(1'h0)] reg3112 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3111 = (1'h0);
  reg [(4'he):(1'h0)] forvar3107 = (1'h0);
  reg [(4'he):(1'h0)] forvar3106 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3102 = (1'h0);
  reg [(4'hb):(1'h0)] reg3098 = (1'h0);
  reg [(4'hf):(1'h0)] reg3097 = (1'h0);
  reg [(5'h19):(1'h0)] reg3096 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3093 = (1'h0);
  reg [(4'h9):(1'h0)] reg3092 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3089 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3088 = (1'h0);
  reg [(4'hf):(1'h0)] reg3086 = (1'h0);
  reg [(5'h13):(1'h0)] reg3084 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3083 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3082 = (1'h0);
  assign y = {wire3216,
                 wire3211,
                 wire3210,
                 wire3209,
                 wire3198,
                 wire3197,
                 wire3196,
                 wire3076,
                 wire4,
                 wire5,
                 wire3071,
                 wire3073,
                 wire3074,
                 wire3078,
                 wire3079,
                 wire3105,
                 wire3193,
                 wire3194,
                 wire3218,
                 wire3219,
                 wire3353,
                 wire3356,
                 reg3080,
                 reg3081,
                 reg3085,
                 reg3087,
                 reg3090,
                 reg3091,
                 reg3094,
                 reg3095,
                 reg3099,
                 reg3100,
                 reg3101,
                 reg3103,
                 reg3104,
                 reg3108,
                 reg3109,
                 reg3110,
                 reg3115,
                 reg3119,
                 reg3122,
                 reg3126,
                 reg3128,
                 reg3129,
                 reg3131,
                 reg3133,
                 reg3134,
                 reg3135,
                 reg3136,
                 reg3140,
                 reg3141,
                 reg3142,
                 reg3144,
                 reg3146,
                 reg3148,
                 reg3149,
                 reg3150,
                 reg3151,
                 reg3153,
                 reg3155,
                 reg3156,
                 reg3157,
                 reg3162,
                 reg3163,
                 reg3165,
                 reg3167,
                 reg3168,
                 reg3170,
                 reg3171,
                 reg3173,
                 reg3176,
                 reg3177,
                 reg3179,
                 reg3181,
                 reg3183,
                 reg3184,
                 reg3186,
                 reg3188,
                 reg3191,
                 reg3203,
                 reg3204,
                 reg3206,
                 reg3207,
                 reg3208,
                 reg3212,
                 reg3213,
                 reg3224,
                 reg3225,
                 reg3229,
                 reg3231,
                 reg3232,
                 reg3234,
                 reg3237,
                 reg3243,
                 reg3244,
                 reg3246,
                 reg3247,
                 reg3249,
                 reg3250,
                 reg3257,
                 reg3259,
                 reg3264,
                 reg3265,
                 reg3266,
                 reg3268,
                 reg3269,
                 reg3272,
                 reg3275,
                 reg3277,
                 reg3280,
                 reg3282,
                 reg3283,
                 reg3284,
                 reg3286,
                 reg3289,
                 reg3290,
                 reg3291,
                 reg3292,
                 reg3295,
                 reg3296,
                 reg3297,
                 reg3299,
                 reg3300,
                 reg3301,
                 reg3302,
                 reg3303,
                 reg3305,
                 reg3308,
                 reg3312,
                 reg3313,
                 reg3315,
                 reg3316,
                 reg3319,
                 reg3323,
                 reg3325,
                 reg3328,
                 reg3332,
                 reg3321,
                 reg3334,
                 reg3335,
                 reg3338,
                 reg3340,
                 reg3341,
                 reg3342,
                 reg3343,
                 reg3345,
                 reg3346,
                 reg3349,
                 reg3352,
                 reg3355,
                 reg3351,
                 reg3350,
                 reg3348,
                 reg3347,
                 reg3344,
                 reg3339,
                 reg3337,
                 reg3336,
                 reg3333,
                 forvar3330,
                 reg3326,
                 forvar3318,
                 reg3331,
                 reg3330,
                 reg3329,
                 reg3327,
                 forvar3326,
                 reg3324,
                 reg3322,
                 forvar3321,
                 reg3320,
                 reg3318,
                 reg3317,
                 reg3314,
                 reg3311,
                 reg3310,
                 reg3309,
                 forvar3307,
                 reg3306,
                 reg3304,
                 reg3298,
                 forvar3296,
                 reg3293,
                 reg3294,
                 forvar3293,
                 reg3288,
                 reg3287,
                 reg3285,
                 reg3276,
                 reg3281,
                 reg3279,
                 reg3278,
                 forvar3276,
                 reg3273,
                 forvar3269,
                 reg3274,
                 forvar3273,
                 reg3271,
                 reg3270,
                 reg3267,
                 reg3263,
                 reg3262,
                 forvar3261,
                 reg3260,
                 reg3258,
                 forvar3256,
                 reg3255,
                 reg3254,
                 reg3253,
                 forvar3252,
                 reg3251,
                 reg3248,
                 forvar3245,
                 forvar3242,
                 reg3241,
                 reg3240,
                 reg3239,
                 reg3238,
                 reg3236,
                 reg3235,
                 reg3233,
                 reg3230,
                 reg3228,
                 reg3227,
                 reg3226,
                 forvar3223,
                 reg3222,
                 forvar3221,
                 forvar3220,
                 reg3215,
                 reg3214,
                 reg3205,
                 reg3202,
                 forvar3201,
                 forvar3200,
                 reg3192,
                 reg3190,
                 reg3189,
                 reg3187,
                 forvar3185,
                 reg3182,
                 reg3180,
                 reg3178,
                 reg3175,
                 reg3174,
                 reg3172,
                 reg3169,
                 reg3166,
                 reg3159,
                 reg3152,
                 forvar3149,
                 reg3145,
                 forvar3139,
                 forvar3131,
                 reg3164,
                 reg3161,
                 reg3160,
                 forvar3159,
                 reg3158,
                 reg3154,
                 forvar3152,
                 reg3147,
                 forvar3145,
                 reg3143,
                 reg3139,
                 reg3138,
                 reg3137,
                 reg3132,
                 reg3130,
                 reg3127,
                 reg3125,
                 reg3124,
                 reg3123,
                 reg3121,
                 forvar3120,
                 forvar3118,
                 forvar3117,
                 reg3116,
                 reg3114,
                 reg3113,
                 reg3112,
                 reg3111,
                 forvar3107,
                 forvar3106,
                 reg3102,
                 reg3098,
                 reg3097,
                 reg3096,
                 reg3093,
                 reg3092,
                 forvar3089,
                 reg3088,
                 reg3086,
                 reg3084,
                 forvar3083,
                 reg3082,
                 (1'h0)};
  assign wire4 = ($signed($unsigned(wire0[(1'h1):(1'h1)])) ? (7'h40) : wire3);
  assign wire5 = (wire4 ?
                     (&$unsigned(($signed(wire0) >> (~&wire4)))) : (($unsigned((^~wire3)) << $signed(wire3[(1'h1):(1'h0)])) > (wire1[(4'hc):(4'h9)] ?
                         (8'hbd) : $unsigned($unsigned(wire3)))));
  module6 #() modinst3072 (wire3071, clk, wire2, wire0, wire3, wire1);
  assign wire3073 = $signed((-wire5[(1'h1):(1'h0)]));
  module2467 #() modinst3075 (.wire2470(wire1), .wire2469(wire2), .clk(clk), .y(wire3074), .wire2471(wire5), .wire2472(wire3), .wire2468(wire3073));
  module2467 #() modinst3077 (wire3076, clk, wire0, wire3, wire2, wire3071, wire5);
  assign wire3078 = wire2[(4'h9):(3'h7)];
  assign wire3079 = {((wire1 + (-(wire5 ? (8'hb0) : wire1))) ?
                            ((|(wire3073 ?
                                wire3 : wire5)) && (8'hb5)) : $unsigned((+$unsigned(wire3071)))),
                        wire5};
  always
    @(posedge clk) begin
      reg3080 <= (({(wire3079[(5'h16):(3'h4)] > wire3073),
              {((8'hbd) ? wire3 : wire3), $unsigned((7'h55))},
              $unsigned($unsigned(wire3074))} <= (~&($unsigned(wire3078) ?
              (^wire3073) : {wire3071}))) ?
          {$unsigned(((-wire3) > wire3079))} : $signed($unsigned(wire3[(4'hd):(4'h9)])));
      reg3081 <= (-{$signed($signed((reg3080 & wire3076)))});
      reg3082 = (~(~|((^~wire3079) >= (^~reg3081))));
      for (forvar3083 = (1'h0); (forvar3083 < (3'h5)); forvar3083 = (forvar3083 + (1'h1)))
        begin
          reg3084 = ($unsigned((~&$unsigned($unsigned((8'h9c))))) ?
              $unsigned(reg3081[(5'h12):(3'h4)]) : $unsigned(wire0));
          if ({($unsigned(reg3080) * $signed(wire3073)),
              (^wire4),
              $signed($unsigned((~^$unsigned(wire3074))))})
            begin
              reg3085 <= (|$unsigned($unsigned({(wire5 ? wire3 : wire0),
                  (+wire2),
                  $unsigned(reg3082)})));
              reg3086 = ((((wire3076 || $unsigned(forvar3083)) >= $signed($signed(wire3078))) & (reg3082 == reg3081[(4'h9):(3'h7)])) & wire5);
            end
          else
            begin
              reg3085 <= wire3076[(4'hc):(2'h2)];
              reg3086 = $signed((~|$unsigned(wire3074)));
              reg3087 <= {(~&{forvar3083}),
                  {$unsigned(reg3086[(3'h6):(1'h0)]),
                      (~^wire3[(4'hb):(3'h5)]),
                      $signed(wire3076[(4'hd):(4'h8)])},
                  $unsigned((((wire3078 & reg3081) ^~ (wire3071 ?
                      wire4 : reg3084)) || ((7'h44) >= $signed(wire3))))};
            end
          reg3088 = $signed($unsigned({(&$unsigned(wire3074)),
              $unsigned(reg3085),
              {(wire5 & forvar3083)}}));
          for (forvar3089 = (1'h0); (forvar3089 < (2'h3)); forvar3089 = (forvar3089 + (1'h1)))
            begin
              reg3090 <= (~^(wire3078 ?
                  (+forvar3083[(2'h2):(1'h0)]) : {{$signed(reg3081),
                          (reg3088 + reg3084),
                          reg3085},
                      wire3[(5'h16):(5'h11)],
                      wire2}));
              reg3091 <= wire3079[(5'h18):(4'hc)];
              reg3092 = ((wire3078 ?
                  reg3090[(3'h7):(2'h3)] : $unsigned(($unsigned(reg3090) << (wire1 ?
                      wire3078 : wire3073)))) > reg3081[(5'h12):(4'h9)]);
            end
          if ({(reg3092[(3'h5):(2'h3)] ?
                  ({(~(7'h45)),
                          (wire3073 >> wire3074),
                          wire3074[(4'hf):(4'hf)]} ?
                      (wire3076[(3'h6):(2'h3)] ^ $unsigned(wire3073)) : reg3080) : reg3087)})
            begin
              reg3093 = {$signed(wire1),
                  $signed((forvar3083[(2'h3):(2'h3)] != ($signed(wire3) << {wire1,
                      wire3071,
                      wire5}))),
                  wire3071[(5'h12):(3'h6)]};
              reg3094 <= (($signed($unsigned(wire2[(1'h0):(1'h0)])) ?
                      (($unsigned(reg3090) ?
                          $signed(wire0) : (~&(8'hbd))) == forvar3083) : ($unsigned((~^wire3076)) > reg3080)) ?
                  $unsigned(wire4[(4'hb):(4'ha)]) : wire3073[(4'h9):(2'h2)]);
              reg3095 <= $signed($unsigned((({(7'h54)} ?
                      {wire3076, wire0, forvar3083} : $unsigned(wire3073)) ?
                  (reg3091[(3'h5):(3'h4)] && (wire3 - wire3073)) : wire3[(3'h6):(3'h4)])));
              reg3096 = forvar3089[(2'h2):(1'h1)];
              reg3097 = (+$unsigned((reg3085[(4'hb):(4'hb)] ?
                  reg3081[(3'h4):(3'h4)] : (~&reg3085[(4'hb):(1'h1)]))));
              reg3098 = (!{$signed(((|reg3094) | reg3081)),
                  (-$unsigned($signed(forvar3083)))});
              reg3099 <= {$unsigned((^~reg3092)),
                  (wire2 ?
                      $signed({(wire3076 <<< reg3087),
                          $unsigned(reg3080),
                          (forvar3089 + wire1)}) : (!((wire3079 ?
                              wire3073 : reg3088) ?
                          $unsigned((7'h47)) : $signed(reg3090)))),
                  ($signed({reg3085[(3'h4):(3'h4)]}) ?
                      (((&reg3084) <<< wire5) ?
                          {(8'ha5)} : $signed((&(8'haf)))) : forvar3089)};
            end
          else
            begin
              reg3093 = (-(8'ha1));
              reg3094 <= ({(((wire1 >>> wire3074) ?
                              (reg3087 | wire3076) : wire3079) ?
                          (wire3074 > (reg3092 ? reg3092 : wire2)) : (7'h4b)),
                      $signed(wire2[(4'hd):(4'hb)]),
                      $unsigned((^(forvar3083 >>> wire5)))} ?
                  $signed((|(reg3090 ?
                      (~^wire3076) : (wire1 >> reg3087)))) : (&(~$signed({wire3071,
                      (7'h49),
                      reg3082}))));
              reg3096 = $signed(((-({reg3092, wire3079} ?
                  wire3 : (wire3073 ?
                      reg3098 : wire3074))) | (((^~wire3071) > $signed(wire3078)) ?
                  $unsigned(wire3076) : forvar3083[(3'h5):(3'h4)])));
              reg3097 = $unsigned({reg3095,
                  $signed((reg3087 >> (wire2 ? (8'hb7) : wire3073)))});
              reg3099 <= $unsigned(((-(wire3076[(3'h4):(1'h1)] ?
                      wire3073[(4'hb):(4'h9)] : (^~reg3084))) ?
                  (~^(reg3088[(5'h16):(2'h3)] ?
                      (wire3076 ?
                          reg3087 : reg3086) : ((8'hb3) + wire3071))) : reg3088));
              reg3100 <= $unsigned((reg3086[(4'h8):(3'h7)] ?
                  (&{wire3073}) : (&$signed(wire3071[(5'h15):(4'hb)]))));
            end
          reg3101 <= ($unsigned($signed((8'hbb))) ? reg3096 : $signed(reg3098));
        end
      reg3102 = ($unsigned((reg3100 < reg3095)) ?
          reg3097[(3'h5):(3'h4)] : (^wire3074));
      reg3103 <= (wire4 ?
          $unsigned((((~^(8'hb8)) << (wire3 & (8'ha3))) ^~ (-(reg3082 ?
              reg3082 : wire5)))) : (reg3102 ?
              {((forvar3083 ? reg3102 : reg3090) ?
                      wire3074[(5'h17):(4'hf)] : $signed(reg3088)),
                  (!reg3080)} : ((8'ha8) >>> ((7'h47) ?
                  {reg3087, forvar3083} : (wire3 < reg3090)))));
      reg3104 <= reg3096;
    end
  assign wire3105 = (7'h46);
  always
    @(posedge clk) begin
      for (forvar3106 = (1'h0); (forvar3106 < (2'h2)); forvar3106 = (forvar3106 + (1'h1)))
        begin
          for (forvar3107 = (1'h0); (forvar3107 < (3'h6)); forvar3107 = (forvar3107 + (1'h1)))
            begin
              reg3108 <= ((~^(reg3080[(3'h4):(1'h1)] ?
                      $signed((wire3105 ~^ wire3105)) : (~&wire3079[(5'h13):(5'h11)]))) ?
                  ($signed((((8'hbc) * wire3105) ?
                          reg3087[(3'h7):(2'h3)] : (wire3078 ?
                              wire3079 : wire3))) ?
                      reg3081 : ({wire3078[(5'h15):(4'hc)]} == (wire5 ?
                          wire4[(2'h3):(1'h1)] : ((8'ha1) ?
                              wire3076 : wire1)))) : $signed(((&(reg3099 && wire3078)) > (reg3103[(2'h2):(1'h0)] + (reg3091 ?
                      wire4 : wire4)))));
              reg3109 <= ($unsigned((+$unsigned($signed(wire1)))) ~^ $unsigned((^~$signed((wire1 ?
                  wire3 : reg3100)))));
              reg3110 <= forvar3106;
              reg3111 = ($signed(reg3087) < $unsigned($unsigned((~^((7'h48) <= reg3081)))));
              reg3112 = ((~^reg3110) | $signed(((reg3104 || reg3101) >> reg3095)));
            end
          reg3113 = ((-$signed(reg3087[(3'h4):(1'h0)])) <= reg3085[(4'h9):(4'h8)]);
          reg3114 = $unsigned((8'ha4));
          reg3115 <= ($unsigned(reg3111[(5'h13):(4'he)]) ?
              ((|(8'hb4)) ?
                  wire3073 : (^~($unsigned((7'h42)) >>> (reg3100 ?
                      (7'h52) : (8'hbf))))) : (+($unsigned((8'h9f)) ?
                  $unsigned((~^wire4)) : reg3112[(1'h0):(1'h0)])));
        end
      reg3116 = ($unsigned((~reg3085[(3'h5):(3'h4)])) * ((~^($signed(forvar3107) * (8'hb6))) ?
          (|(+(wire3073 ? wire3076 : reg3109))) : (reg3094 > $signed(((7'h54) ?
              wire3071 : reg3085)))));
    end
  always
    @(posedge clk) begin
      for (forvar3117 = (1'h0); (forvar3117 < (1'h1)); forvar3117 = (forvar3117 + (1'h1)))
        begin
          for (forvar3118 = (1'h0); (forvar3118 < (3'h4)); forvar3118 = (forvar3118 + (1'h1)))
            begin
              reg3119 <= (forvar3117[(3'h5):(1'h0)] ?
                  $unsigned(reg3100) : wire3073);
            end
          for (forvar3120 = (1'h0); (forvar3120 < (3'h4)); forvar3120 = (forvar3120 + (1'h1)))
            begin
              reg3121 = wire3073[(2'h3):(1'h1)];
            end
          reg3122 <= wire5;
          if (($unsigned($unsigned(($signed(wire3) ?
              $unsigned((8'hab)) : $unsigned((7'h41))))) - $unsigned((((reg3100 >> wire2) ~^ $unsigned(reg3101)) ?
              ((|reg3110) <<< reg3103) : reg3095[(1'h1):(1'h0)]))))
            begin
              reg3123 = $signed((~$unsigned({(^~(8'ha6)),
                  $unsigned(reg3087),
                  $unsigned(forvar3118)})));
              reg3124 = (((~{(wire2 ^ (7'h41)), ((8'ha6) < wire3073)}) ?
                  $unsigned($signed($signed(wire3105))) : ({(|reg3109),
                      wire3} * wire4[(4'ha):(1'h1)])) + forvar3120[(4'hc):(3'h7)]);
              reg3125 = (reg3085 << (reg3115 ^ $signed((-$unsigned(wire4)))));
              reg3126 <= reg3087[(3'h4):(1'h0)];
              reg3127 = (|{({$signed(wire3105), (!reg3081)} ?
                      ((~reg3125) ^~ {reg3099}) : (^~$signed(wire5))),
                  (~^$unsigned($signed((7'h56))))});
            end
          else
            begin
              reg3123 = ($unsigned((^$unsigned($signed(forvar3120)))) || ($unsigned(reg3094[(3'h6):(3'h6)]) ^~ ($unsigned($signed(reg3122)) ?
                  (!(forvar3120 ?
                      reg3122 : (8'h9e))) : ((^reg3095) != reg3104[(5'h16):(5'h12)]))));
              reg3124 = reg3080;
            end
          reg3128 <= $unsigned($unsigned((wire1[(1'h1):(1'h0)] < ({reg3110,
              reg3127,
              wire4} || wire3073[(2'h2):(1'h1)]))));
        end
      reg3129 <= $unsigned(($signed(wire3078[(2'h3):(1'h1)]) ?
          reg3119[(5'h12):(5'h10)] : (!reg3081)));
      if ((8'hb8))
        begin
          if ((~|$signed($signed(wire3078))))
            begin
              reg3130 = (reg3127 ? reg3125 : $signed($unsigned(reg3095)));
              reg3131 <= reg3110[(1'h1):(1'h0)];
              reg3132 = $signed(reg3103[(4'h9):(3'h6)]);
            end
          else
            begin
              reg3131 <= (~wire1[(1'h0):(1'h0)]);
              reg3133 <= forvar3118;
              reg3134 <= (~|$signed($unsigned($unsigned((reg3130 ?
                  (7'h52) : reg3085)))));
              reg3135 <= (7'h4d);
              reg3136 <= $signed((~(8'hb0)));
              reg3137 = (~&(~|$signed(($unsigned((8'hb5)) ?
                  $unsigned(reg3130) : reg3127[(3'h4):(1'h1)]))));
            end
          reg3138 = wire4;
          if ((+$unsigned({reg3101[(3'h6):(2'h3)]})))
            begin
              reg3139 = wire1;
              reg3140 <= (~&((~^(~^(-wire3074))) ~^ $unsigned(reg3129)));
              reg3141 <= reg3137[(2'h2):(1'h0)];
              reg3142 <= (reg3108 ?
                  ((8'hac) ?
                      (((~&reg3080) ^ (wire2 <= wire0)) & $signed((reg3133 - reg3138))) : reg3119) : reg3119);
              reg3143 = reg3123;
            end
          else
            begin
              reg3139 = $signed(reg3121[(3'h5):(2'h3)]);
              reg3143 = $unsigned(reg3095[(4'h8):(3'h6)]);
            end
          reg3144 <= reg3124[(5'h13):(4'h8)];
          for (forvar3145 = (1'h0); (forvar3145 < (3'h5)); forvar3145 = (forvar3145 + (1'h1)))
            begin
              reg3146 <= wire3078;
              reg3147 = (~reg3099);
              reg3148 <= $unsigned(reg3131[(4'ha):(4'h9)]);
              reg3149 <= reg3122;
              reg3150 <= (($signed($signed($unsigned(wire1))) < (reg3144[(3'h7):(3'h5)] != ($unsigned(wire3105) ?
                      forvar3120[(1'h1):(1'h1)] : (wire3073 != (7'h52))))) ?
                  wire4 : forvar3118[(3'h4):(3'h4)]);
              reg3151 <= $signed($unsigned($signed(reg3101)));
            end
          for (forvar3152 = (1'h0); (forvar3152 < (2'h2)); forvar3152 = (forvar3152 + (1'h1)))
            begin
              reg3153 <= reg3103[(4'ha):(4'h8)];
              reg3154 = wire4;
              reg3155 <= (~reg3126[(1'h1):(1'h1)]);
              reg3156 <= $signed(reg3155[(2'h3):(2'h3)]);
              reg3157 <= reg3149[(1'h1):(1'h1)];
              reg3158 = (!$unsigned({(&(reg3134 ? reg3126 : reg3144)),
                  ($unsigned(reg3143) >> wire2)}));
            end
          for (forvar3159 = (1'h0); (forvar3159 < (3'h5)); forvar3159 = (forvar3159 + (1'h1)))
            begin
              reg3160 = reg3135[(2'h2):(2'h2)];
              reg3161 = {$unsigned(($unsigned((reg3094 || reg3109)) + $signed((&reg3156)))),
                  reg3150[(2'h2):(1'h0)]};
              reg3162 <= (reg3131[(2'h2):(2'h2)] ?
                  $unsigned($unsigned((((8'ha1) ? (8'hba) : (7'h53)) ?
                      reg3155 : ((8'ha2) ?
                          reg3151 : reg3131)))) : reg3149[(1'h1):(1'h0)]);
              reg3163 <= $signed(reg3124);
              reg3164 = $signed(wire5[(5'h11):(2'h2)]);
              reg3165 <= $unsigned(reg3129[(3'h6):(2'h3)]);
            end
        end
      else
        begin
          reg3130 = reg3094;
          for (forvar3131 = (1'h0); (forvar3131 < (3'h5)); forvar3131 = (forvar3131 + (1'h1)))
            begin
              reg3132 = (~&reg3094[(2'h2):(1'h1)]);
              reg3137 = {(8'hb2)};
              reg3138 = {$unsigned(((reg3136 ? reg3087 : $signed(wire2)) ?
                      {$unsigned(reg3123)} : (reg3119[(2'h2):(1'h1)] <= {(8'h9d),
                          (8'hbb),
                          reg3141})))};
            end
          for (forvar3139 = (1'h0); (forvar3139 < (1'h0)); forvar3139 = (forvar3139 + (1'h1)))
            begin
              reg3140 <= (((^(^~(forvar3159 <= reg3094))) <<< reg3158) >= (!reg3147));
              reg3143 = reg3085[(4'hd):(4'hb)];
              reg3144 <= $signed((7'h54));
              reg3145 = wire4[(2'h3):(1'h0)];
              reg3147 = $signed((^$unsigned((^~{reg3136, reg3149, reg3104}))));
              reg3148 <= wire3079;
            end
          for (forvar3149 = (1'h0); (forvar3149 < (3'h4)); forvar3149 = (forvar3149 + (1'h1)))
            begin
              reg3152 = ((8'h9c) ? reg3135[(4'hb):(3'h7)] : $signed(reg3151));
              reg3153 <= reg3163[(4'he):(4'hc)];
              reg3154 = (((((!reg3136) <= $unsigned((7'h42))) ?
                          reg3115 : ((8'ha5) ?
                              $unsigned(reg3152) : reg3146[(5'h16):(3'h4)])) ?
                      wire1[(4'hb):(2'h2)] : $signed(reg3129[(5'h12):(4'h9)])) ?
                  ((({wire1} ? (|reg3161) : $unsigned(reg3161)) ?
                      (~&$signed(reg3121)) : (~^reg3140)) <= reg3140) : (~&(~reg3127[(1'h1):(1'h1)])));
              reg3158 = reg3126;
            end
          reg3159 = reg3134[(5'h11):(4'hd)];
          reg3162 <= (reg3164 ^~ (reg3149[(2'h3):(1'h1)] ~^ ($unsigned($unsigned(reg3145)) ?
              (+$unsigned(wire3079)) : wire5)));
          reg3163 <= (8'hbc);
        end
      reg3166 = {forvar3131[(5'h19):(4'hf)],
          ({wire0[(5'h18):(1'h1)],
              {{reg3125, (8'ha2), reg3138}, $unsigned(reg3081)},
              $signed((wire3078 || reg3132))} & reg3148),
          $unsigned($unsigned((!(!reg3164))))};
      if ((reg3123 == reg3109[(4'hf):(3'h5)]))
        begin
          reg3167 <= $unsigned((reg3143 ?
              $signed((~&$unsigned(reg3159))) : {(~&reg3150),
                  (8'ha2),
                  reg3140[(4'hb):(3'h6)]}));
          reg3168 <= reg3152[(4'ha):(4'h8)];
        end
      else
        begin
          reg3169 = $unsigned((7'h4d));
          reg3170 <= {(-(!(reg3151[(3'h5):(3'h5)] >>> (~|reg3163)))),
              ((((reg3151 && forvar3117) ?
                  {reg3160, forvar3152, (8'hba)} : {(7'h51),
                      reg3119}) >= $signed((wire3076 ?
                  (8'h9f) : reg3132))) * $signed(wire2))};
          reg3171 <= ($signed(reg3151[(1'h1):(1'h1)]) ?
              (($unsigned(reg3104) ? (|(~^reg3148)) : reg3162) ?
                  wire3073 : ((^{reg3155, (7'h57), (8'hba)}) ?
                      $unsigned(reg3133[(3'h7):(3'h6)]) : reg3091[(3'h6):(2'h3)])) : (($unsigned($signed(reg3122)) * {reg3110,
                      reg3101[(4'hb):(2'h3)]}) ?
                  wire1 : reg3170[(3'h4):(1'h1)]));
          reg3172 = (7'h53);
          if (($unsigned($unsigned({(wire3074 ? reg3169 : reg3123), reg3145})) ?
              $signed((~|{(reg3135 ? reg3161 : reg3123),
                  $signed((8'haa))})) : {$signed((^{reg3119,
                      forvar3145,
                      forvar3149})),
                  $unsigned($signed(wire3076)),
                  $unsigned(reg3124)}))
            begin
              reg3173 <= reg3103;
              reg3174 = $signed((!($unsigned(reg3142[(4'hf):(3'h5)]) > reg3090[(2'h2):(2'h2)])));
              reg3175 = forvar3120[(2'h3):(2'h2)];
            end
          else
            begin
              reg3174 = $signed(($signed($signed((reg3104 | reg3126))) <<< (!$unsigned({wire3074}))));
              reg3176 <= reg3122;
              reg3177 <= (((^~$unsigned((8'hbe))) != reg3167) - (~^(~wire3078[(1'h0):(1'h0)])));
              reg3178 = (|(wire3105 ?
                  $unsigned(((~|wire4) >= $unsigned(reg3134))) : {(~&(^~wire3105)),
                      $signed((~^reg3137)),
                      reg3150[(2'h3):(1'h0)]}));
              reg3179 <= $signed(({($signed(reg3126) > (8'hb1)),
                  reg3133[(4'h8):(4'h8)],
                  reg3100} - $signed(((reg3126 ?
                  (8'hb5) : reg3130) & $unsigned(reg3164)))));
              reg3180 = forvar3139[(1'h0):(1'h0)];
              reg3181 <= forvar3152[(4'h8):(2'h2)];
            end
        end
      if ($unsigned((|$unsigned(((7'h42) <= reg3170[(4'h8):(1'h1)])))))
        begin
          reg3182 = (8'ha8);
        end
      else
        begin
          reg3182 = $unsigned(((reg3156 * reg3123) - reg3174[(4'hd):(4'h8)]));
          reg3183 <= {{((reg3169 << (~^reg3163)) ?
                      $unsigned($unsigned((8'ha0))) : reg3162),
                  (&({reg3180, reg3157, reg3153} * reg3174[(5'h16):(1'h0)])),
                  reg3099[(1'h0):(1'h0)]},
              (+$unsigned((~&reg3152[(2'h3):(1'h0)])))};
          reg3184 <= reg3139[(3'h5):(3'h4)];
        end
      for (forvar3185 = (1'h0); (forvar3185 < (1'h1)); forvar3185 = (forvar3185 + (1'h1)))
        begin
          if (forvar3185)
            begin
              reg3186 <= $signed($unsigned(reg3081[(1'h1):(1'h0)]));
              reg3187 = (~|((^wire5[(4'h8):(3'h6)]) << ($unsigned(((8'hbe) ?
                  (8'hba) : reg3081)) >> {$signed(reg3183),
                  $unsigned(reg3175),
                  reg3149})));
              reg3188 <= {$unsigned({$unsigned($unsigned(reg3125))})};
              reg3189 = reg3124[(4'h9):(3'h4)];
              reg3190 = $unsigned(($unsigned({$signed(reg3184),
                  $signed(reg3136)}) >= $signed(({(8'had)} ?
                  (reg3164 <<< reg3179) : {wire1, reg3171, (8'ha9)}))));
              reg3191 <= (7'h4a);
              reg3192 = reg3143[(4'hc):(1'h1)];
            end
          else
            begin
              reg3186 <= (8'ha7);
            end
        end
    end
  assign wire3193 = (($unsigned(((&reg3100) ?
                        {(7'h43)} : (~^(8'hbc)))) << ((~(&reg3176)) ?
                        reg3087 : reg3094)) == (~|$unsigned((|$signed(reg3094)))));
  module2467 #() modinst3195 (wire3194, clk, reg3103, reg3176, reg3153, reg3171, wire1);
  assign wire3196 = (-(^((reg3129[(3'h5):(2'h3)] ^~ ((7'h4e) == wire1)) ?
                        $signed({reg3165,
                            reg3173,
                            reg3094}) : $unsigned(reg3151[(2'h3):(2'h2)]))));
  assign wire3197 = ((reg3094[(1'h1):(1'h1)] ?
                            {wire3073[(4'ha):(4'h8)]} : reg3165) ?
                        (!$signed(reg3119)) : wire3078[(3'h5):(2'h3)]);
  module71 #() modinst3199 (wire3198, clk, reg3122, reg3167, reg3104, wire3074, wire5, reg3165);
  always
    @(posedge clk) begin
      for (forvar3200 = (1'h0); (forvar3200 < (1'h1)); forvar3200 = (forvar3200 + (1'h1)))
        begin
          for (forvar3201 = (1'h0); (forvar3201 < (2'h2)); forvar3201 = (forvar3201 + (1'h1)))
            begin
              reg3202 = $unsigned({{{(-reg3167)},
                      ($signed(wire3193) < reg3183),
                      $unsigned(reg3167[(3'h4):(1'h0)])},
                  ({(reg3179 ? (8'hbb) : (8'had)),
                      (~reg3184)} + $signed((-(7'h4b))))});
              reg3203 <= reg3133;
              reg3204 <= (~&$unsigned(forvar3201[(4'hf):(1'h1)]));
              reg3205 = wire3194;
            end
          reg3206 <= (|$signed({reg3162[(2'h2):(1'h1)],
              $signed({reg3104, reg3108})}));
        end
      reg3207 <= (~reg3100);
      reg3208 <= reg3168;
    end
  assign wire3209 = (^~(($unsigned((|reg3162)) ?
                            $unsigned($signed(reg3208)) : $unsigned((wire3197 <= (7'h49)))) ?
                        (!reg3099) : (($signed(reg3203) ?
                            $signed(reg3179) : $signed(reg3140)) | {$unsigned((7'h4d))})));
  assign wire3210 = (((!(wire3194[(2'h2):(2'h2)] ? reg3148 : reg3184)) ?
                            $signed($signed($signed((8'hb5)))) : (reg3149[(2'h2):(2'h2)] ~^ wire0)) ?
                        ((wire3078[(5'h12):(3'h4)] + ($signed(reg3173) ?
                                (reg3087 ? reg3148 : reg3131) : {wire0,
                                    (8'had),
                                    reg3155})) ?
                            $unsigned({(reg3080 > reg3095)}) : (((7'h53) <<< $signed((7'h54))) ?
                                $signed($unsigned(reg3188)) : {(!(7'h4b)),
                                    $signed(reg3173),
                                    $signed(reg3085)})) : reg3177[(4'hd):(4'ha)]);
  assign wire3211 = $signed((-{({reg3148} || (reg3134 ^ reg3156)),
                        (&$signed(wire3079)),
                        wire3071}));
  always
    @(posedge clk) begin
      reg3212 <= {(wire3209 >>> (7'h43)),
          ((^$unsigned($signed(reg3100))) ?
              {(reg3140 + (~^reg3131))} : (^~$unsigned($unsigned(wire3105))))};
      reg3213 <= {{wire3210[(5'h16):(4'hc)],
              $signed($signed((wire3071 < reg3090)))},
          reg3165};
      reg3214 = wire1[(4'hd):(4'hd)];
      reg3215 = reg3167;
    end
  module326 #() modinst3217 (.wire327(reg3099), .wire328(reg3181), .y(wire3216), .wire330(wire3197), .wire331(reg3080), .wire329(reg3153), .clk(clk));
  assign wire3218 = reg3184[(2'h2):(1'h1)];
  assign wire3219 = (~^((wire3073 <<< reg3186) | wire3197));
  always
    @(posedge clk) begin
      for (forvar3220 = (1'h0); (forvar3220 < (3'h5)); forvar3220 = (forvar3220 + (1'h1)))
        begin
          for (forvar3221 = (1'h0); (forvar3221 < (2'h2)); forvar3221 = (forvar3221 + (1'h1)))
            begin
              reg3222 = reg3153[(1'h1):(1'h1)];
            end
          for (forvar3223 = (1'h0); (forvar3223 < (3'h5)); forvar3223 = (forvar3223 + (1'h1)))
            begin
              reg3224 <= reg3162;
              reg3225 <= {(8'ha2),
                  reg3162[(4'he):(2'h3)],
                  ($signed($unsigned($signed(reg3207))) ?
                      ({(reg3146 != reg3100),
                          (wire3079 ? reg3099 : (7'h4f))} > ((+reg3179) ?
                          reg3090 : reg3186[(4'hd):(3'h4)])) : (~&$signed({wire3198})))};
              reg3226 = $signed(wire3197);
              reg3227 = (($unsigned(wire3219[(4'h8):(1'h1)]) ?
                      $signed(wire5) : {(~|(~&reg3222))}) ?
                  (((~&(reg3212 | reg3144)) | (-(wire3209 == reg3141))) ?
                      $signed($unsigned(reg3225[(2'h3):(1'h1)])) : (wire3193[(4'hb):(2'h2)] ?
                          (~|$unsigned(wire3218)) : ((reg3122 < wire1) - (7'h40)))) : reg3204);
              reg3228 = $signed({({(reg3144 ? reg3146 : wire3219),
                          $unsigned(wire3071)} ?
                      ((wire5 ^~ wire3073) + wire2) : (^$unsigned(reg3146)))});
              reg3229 <= (~&(reg3183[(2'h3):(1'h1)] != (($unsigned(reg3080) << (7'h44)) ?
                  $signed($unsigned(reg3228)) : $signed($unsigned(reg3149)))));
            end
          reg3230 = reg3142[(4'ha):(1'h0)];
          reg3231 <= {{(($unsigned(reg3126) && (8'hb1)) == wire3198),
                  (~&$signed($signed(forvar3220)))}};
          if (reg3176)
            begin
              reg3232 <= (^((&((-wire3198) ^ $signed(wire3210))) && $unsigned($signed($unsigned(wire3105)))));
              reg3233 = (&{(reg3104 ?
                      $unsigned(reg3151[(3'h5):(3'h4)]) : (|(reg3229 ?
                          reg3181 : wire4))),
                  (~$unsigned((7'h44)))});
              reg3234 <= (((reg3081 ?
                      ((!reg3231) >>> (reg3212 ?
                          reg3146 : wire3074)) : (&(reg3136 ?
                          reg3140 : reg3184))) ?
                  reg3153 : wire3078) <<< (&($signed(reg3233[(4'hb):(4'h8)]) ?
                  wire3074[(4'hc):(2'h2)] : reg3115)));
              reg3235 = $unsigned((reg3207 ?
                  (7'h55) : ({$signed(reg3231),
                      $signed(reg3081)} < $signed(reg3141))));
            end
          else
            begin
              reg3233 = {$signed(reg3206),
                  reg3233[(5'h1d):(4'hf)],
                  $unsigned((^$signed(wire5)))};
              reg3235 = (~(^(reg3191[(5'h1f):(4'hd)] ?
                  (~(reg3153 ?
                      reg3129 : wire3209)) : $signed($unsigned(reg3163)))));
              reg3236 = $unsigned({((reg3233[(3'h7):(1'h1)] >= (reg3232 >>> (7'h4f))) ?
                      $unsigned(wire3209) : ({reg3153} ?
                          reg3095[(4'h8):(1'h1)] : reg3227)),
                  $unsigned($signed((reg3177 ^~ reg3188))),
                  $signed((^(^~wire5)))});
              reg3237 <= {{(~^$signed($unsigned(reg3177))),
                      ({$signed(wire3194),
                          (reg3142 ? reg3167 : reg3203)} * reg3235)},
                  ({($unsigned(reg3162) ?
                          reg3188[(3'h6):(1'h1)] : (~&wire3))} ~^ (8'hbf))};
              reg3238 = $signed(reg3204);
              reg3239 = ((!reg3208[(4'hc):(4'ha)]) ^~ ($signed(($unsigned(reg3146) & wire5)) >>> (reg3184[(5'h12):(4'hc)] > $unsigned((8'hb5)))));
            end
          reg3240 = ($signed((8'ha7)) ?
              reg3173[(3'h7):(3'h7)] : reg3134[(4'hb):(2'h2)]);
        end
      reg3241 = (+wire3219[(3'h7):(2'h3)]);
      for (forvar3242 = (1'h0); (forvar3242 < (3'h5)); forvar3242 = (forvar3242 + (1'h1)))
        begin
          reg3243 <= ({$signed($signed($signed(reg3094)))} ?
              (reg3184[(5'h11):(4'hf)] ?
                  $unsigned(($unsigned(wire3073) == (reg3141 >> reg3230))) : ((reg3135 ?
                      reg3168 : ((7'h52) ?
                          reg3225 : wire3079)) > (((8'h9e) ~^ reg3239) ^ (7'h51)))) : ((reg3109 <= ($unsigned((8'ha3)) ?
                      (reg3129 ^~ forvar3242) : (&reg3103))) ?
                  reg3095 : (forvar3242 <= $unsigned($signed(reg3126)))));
          reg3244 <= $signed({$signed((reg3110 ?
                  $unsigned(forvar3223) : $unsigned(wire2))),
              $unsigned($unsigned((reg3142 ? wire3194 : reg3224)))});
        end
      for (forvar3245 = (1'h0); (forvar3245 < (1'h0)); forvar3245 = (forvar3245 + (1'h1)))
        begin
          if ((((reg3103[(4'h9):(3'h4)] ?
                  (~|{wire3076}) : (|wire3197[(5'h19):(5'h19)])) * ($signed({reg3080}) & $unsigned((reg3226 ?
                  (7'h55) : reg3232)))) ?
              reg3208[(1'h0):(1'h0)] : reg3101))
            begin
              reg3246 <= (~(|(~wire1[(4'h9):(2'h2)])));
              reg3247 <= ((~&(|$unsigned((^reg3233)))) ?
                  reg3240[(2'h3):(2'h3)] : ((((~reg3228) > (reg3237 ?
                      wire5 : forvar3223)) ^~ {((7'h48) | (7'h4d))}) < (~^($signed(reg3103) ?
                      reg3135 : $signed((8'hab))))));
              reg3248 = reg3109;
            end
          else
            begin
              reg3248 = forvar3245[(5'h11):(1'h1)];
              reg3249 <= wire3196[(1'h0):(1'h0)];
              reg3250 <= ($unsigned(($signed((^~reg3246)) ?
                      (-$unsigned(wire3196)) : (reg3081[(5'h11):(3'h6)] ?
                          (wire3216 ? (8'hb9) : reg3115) : forvar3221))) ?
                  (^(~|(reg3228[(2'h3):(1'h0)] << (-wire4)))) : (8'ha9));
              reg3251 = $signed(reg3081[(5'h11):(3'h5)]);
            end
          for (forvar3252 = (1'h0); (forvar3252 < (3'h6)); forvar3252 = (forvar3252 + (1'h1)))
            begin
              reg3253 = reg3240;
              reg3254 = (wire3196[(1'h0):(1'h0)] - $unsigned(((8'ha7) && reg3104)));
              reg3255 = $unsigned($unsigned($signed($signed({reg3119,
                  reg3235}))));
            end
          for (forvar3256 = (1'h0); (forvar3256 < (3'h4)); forvar3256 = (forvar3256 + (1'h1)))
            begin
              reg3257 <= {((|$unsigned(wire3211[(5'h11):(1'h1)])) ?
                      ($unsigned({reg3156,
                          reg3227}) >>> reg3091) : reg3254[(4'hc):(1'h1)])};
              reg3258 = (~&reg3087);
              reg3259 <= forvar3242;
              reg3260 = (|((+$unsigned((^(7'h48)))) ?
                  (~^$unsigned($unsigned(wire3219))) : (($unsigned(forvar3223) ^~ reg3237[(5'h12):(3'h5)]) == reg3234)));
            end
          for (forvar3261 = (1'h0); (forvar3261 < (1'h0)); forvar3261 = (forvar3261 + (1'h1)))
            begin
              reg3262 = $unsigned(($unsigned(((8'hb8) || $signed(wire5))) ?
                  (((8'hba) ?
                      (reg3101 > wire3210) : (8'haa)) <<< ((wire3196 & reg3234) ?
                      $unsigned(reg3184) : (8'hb0))) : (^(7'h49))));
              reg3263 = (+(~reg3250));
              reg3264 <= ((^~{(((8'hb7) ? reg3244 : reg3140) == (&reg3129)),
                  $signed((reg3227 ? reg3254 : (8'hbc))),
                  reg3204[(1'h0):(1'h0)]}) == ((((reg3136 ? reg3207 : reg3165) ?
                      reg3155[(3'h5):(2'h3)] : (wire3071 ? reg3232 : reg3155)) ?
                  (!$unsigned(reg3244)) : ({wire3105,
                      (7'h49)} ^~ (^~forvar3221))) == $unsigned($unsigned({reg3207,
                  reg3103,
                  wire3211}))));
              reg3265 <= (reg3095[(4'h9):(2'h2)] || {({reg3155[(3'h4):(2'h3)]} ?
                      reg3179[(4'ha):(3'h6)] : ($signed(reg3253) ?
                          (-wire3079) : reg3188[(4'hb):(2'h3)]))});
            end
          reg3266 <= (&(!(!reg3094[(3'h7):(2'h3)])));
        end
      if (($unsigned(reg3204) ? reg3091[(4'he):(2'h2)] : reg3254))
        begin
          if (({((wire5 ^ $unsigned(reg3148)) ?
                  $unsigned((~^reg3250)) : (~^$signed(wire3193))),
              reg3227[(4'h8):(2'h3)]} << (8'ha9)))
            begin
              reg3267 = (($unsigned(reg3135) - $signed(($unsigned(reg3080) || reg3163))) ?
                  (|$signed(reg3264)) : ((+(reg3207[(5'h14):(3'h5)] ^ (!reg3162))) - wire3079[(1'h0):(1'h0)]));
              reg3268 <= (reg3259 ?
                  reg3090 : (wire3216 ?
                      $signed($unsigned(reg3101)) : $unsigned($signed(reg3126[(3'h4):(2'h2)]))));
              reg3269 <= reg3191[(4'hd):(4'hb)];
              reg3270 = reg3235[(1'h0):(1'h0)];
              reg3271 = (!reg3167);
              reg3272 <= wire3219[(3'h4):(3'h4)];
            end
          else
            begin
              reg3267 = (&reg3173[(4'hc):(2'h3)]);
              reg3268 <= wire4[(4'ha):(3'h4)];
              reg3269 <= wire1;
              reg3272 <= $signed({$signed($signed($unsigned(reg3091))),
                  $signed((&(reg3235 ? reg3162 : (7'h4c)))),
                  reg3269[(4'hc):(2'h3)]});
            end
          for (forvar3273 = (1'h0); (forvar3273 < (3'h6)); forvar3273 = (forvar3273 + (1'h1)))
            begin
              reg3274 = $signed(reg3179);
            end
        end
      else
        begin
          reg3268 <= (-(((7'h45) * $unsigned((reg3222 ~^ reg3177))) ?
              reg3156[(1'h1):(1'h0)] : $signed(wire3073)));
          for (forvar3269 = (1'h0); (forvar3269 < (1'h0)); forvar3269 = (forvar3269 + (1'h1)))
            begin
              reg3270 = (8'ha8);
              reg3272 <= {(+forvar3269[(2'h2):(1'h0)]), reg3234};
              reg3273 = (reg3167[(3'h7):(2'h3)] >> $unsigned($signed(((|reg3104) ?
                  reg3150[(2'h2):(2'h2)] : $signed(reg3100)))));
              reg3275 <= {(+$signed(((reg3272 ? reg3091 : reg3250) ?
                      (reg3267 ? reg3094 : reg3119) : $unsigned(reg3251)))),
                  $unsigned((((wire3 << reg3109) ? (7'h48) : reg3241) ?
                      reg3155 : {reg3191[(5'h17):(3'h4)]}))};
            end
        end
    end
  always
    @(posedge clk) begin
      if ({(reg3246 ?
              (reg3173 ?
                  $unsigned($unsigned((7'h49))) : ((reg3104 ? wire5 : reg3140) ?
                      $unsigned(reg3237) : (wire3219 ?
                          reg3213 : reg3091))) : $unsigned((^(reg3207 >> reg3268)))),
          (~&$signed(reg3148))})
        begin
          for (forvar3276 = (1'h0); (forvar3276 < (3'h4)); forvar3276 = (forvar3276 + (1'h1)))
            begin
              reg3277 <= (^($unsigned(($signed(wire3073) ?
                  $unsigned((7'h42)) : (reg3234 ?
                      reg3212 : (8'hbb)))) != reg3151));
              reg3278 = (^~$unsigned(reg3131[(4'ha):(4'h9)]));
              reg3279 = (reg3148[(4'ha):(2'h3)] ?
                  (!$signed(wire3194)) : reg3133);
            end
          reg3280 <= wire1;
          reg3281 = {reg3247[(4'ha):(4'h9)],
              reg3181[(4'hd):(4'h9)],
              ((-$unsigned(reg3162)) ?
                  {$signed((reg3188 ? wire3078 : (8'hb3)))} : reg3151)};
        end
      else
        begin
          reg3276 = ($unsigned(reg3148) ?
              wire3105[(5'h10):(4'hb)] : reg3109[(4'hf):(3'h4)]);
          if ((&((8'h9d) ? reg3265 : (!$unsigned({(8'hbc)})))))
            begin
              reg3278 = {(reg3191[(4'hf):(4'he)] ?
                      reg3276[(2'h3):(2'h2)] : reg3213[(2'h2):(2'h2)])};
              reg3279 = reg3278[(2'h2):(1'h1)];
              reg3280 <= (((~^((^wire3197) && $signed(reg3153))) >= reg3229) && ((7'h53) ?
                  $signed((8'ha2)) : {reg3173[(1'h1):(1'h0)]}));
              reg3282 <= wire3076;
              reg3283 <= $signed(reg3229);
              reg3284 <= (($signed(reg3149[(1'h0):(1'h0)]) + reg3173) <= reg3176);
            end
          else
            begin
              reg3278 = $signed(reg3085[(5'h11):(3'h4)]);
              reg3280 <= wire3211[(4'hb):(2'h3)];
              reg3282 <= ((^~{{{reg3224}, (~&reg3279), ((8'h9d) >>> reg3265)},
                  reg3237}) && $unsigned(reg3266[(1'h0):(1'h0)]));
              reg3285 = $signed(reg3229);
              reg3286 <= (!(reg3100[(4'ha):(1'h0)] ?
                  reg3279[(3'h4):(2'h2)] : ((((8'hb0) || wire3209) ?
                          $unsigned((8'h9d)) : (reg3184 ? wire3219 : reg3119)) ?
                      wire3071 : reg3191)));
              reg3287 = wire3;
              reg3288 = $signed((~&$signed($signed((reg3259 ?
                  reg3144 : wire3196)))));
            end
          reg3289 <= ({reg3135[(1'h0):(1'h0)],
              reg3206[(5'h15):(3'h6)]} | $signed(($unsigned($unsigned((7'h4d))) ?
              ((7'h53) && (reg3279 ? wire2 : reg3246)) : ({reg3179,
                      reg3257,
                      reg3149} ?
                  (&reg3284) : (reg3153 ? (8'hb9) : reg3110)))));
        end
      reg3290 <= $unsigned($unsigned((reg3150[(3'h5):(2'h3)] ?
          ((wire1 ? reg3213 : reg3151) & {(7'h44),
              wire3105,
              (8'hb5)}) : $unsigned((wire3209 ? reg3126 : wire3219)))));
      reg3291 <= reg3278;
      reg3292 <= (reg3191[(5'h10):(3'h6)] <= reg3144[(1'h1):(1'h1)]);
      if ({{$signed({$unsigned(reg3144)}),
              wire3194[(3'h4):(1'h0)],
              $unsigned($unsigned(wire3210))}})
        begin
          for (forvar3293 = (1'h0); (forvar3293 < (3'h5)); forvar3293 = (forvar3293 + (1'h1)))
            begin
              reg3294 = reg3103;
              reg3295 <= $unsigned((|reg3286[(4'he):(4'he)]));
            end
          reg3296 <= reg3104;
        end
      else
        begin
          reg3293 = (~(~|{(~$unsigned(reg3181)),
              ({reg3104, reg3288, reg3115} ?
                  (^(8'had)) : reg3265[(4'hc):(3'h7)])}));
          reg3294 = ($signed((+$unsigned((wire3071 ? (8'ha2) : reg3157)))) ?
              {$signed(reg3115),
                  (reg3285 ?
                      ((reg3186 || reg3259) ~^ $signed(reg3142)) : reg3128[(5'h15):(3'h7)])} : ((&(~^reg3087[(2'h3):(1'h1)])) ?
                  (~^(reg3153[(2'h2):(1'h0)] * (~&reg3115))) : {$unsigned((&reg3168))}));
          reg3295 <= ($unsigned(reg3144) ?
              ((reg3134[(5'h16):(5'h16)] ~^ {reg3136[(3'h6):(2'h3)],
                  ((8'hbf) ? wire3076 : reg3225)}) || reg3287) : ((|reg3157) ?
                  ($unsigned($signed(reg3285)) | reg3146) : (|(!$signed((8'hbe))))));
          for (forvar3296 = (1'h0); (forvar3296 < (3'h5)); forvar3296 = (forvar3296 + (1'h1)))
            begin
              reg3297 <= (7'h4f);
              reg3298 = ({((^~{reg3156,
                      reg3266}) <<< forvar3296[(1'h1):(1'h1)]),
                  $unsigned(reg3297[(3'h7):(3'h4)]),
                  {($signed(reg3173) - (wire0 ~^ (8'hbd))),
                      (reg3108[(3'h5):(3'h5)] ^~ (wire3218 | (7'h40))),
                      (|wire3211[(5'h1a):(2'h2)])}} > $unsigned($unsigned((wire3074[(4'he):(3'h4)] ?
                  (wire2 ? reg3156 : reg3297) : $unsigned(reg3168)))));
              reg3299 <= {{{reg3163[(3'h7):(1'h1)],
                          ((wire3076 ? reg3272 : reg3272) ^~ {reg3134,
                              reg3144,
                              reg3165}),
                          ($signed((8'had)) - $signed(reg3204))},
                      reg3162[(4'h9):(1'h0)],
                      reg3281[(1'h0):(1'h0)]},
                  (($signed((7'h55)) >= ($signed(reg3104) >> reg3229[(5'h11):(4'ha)])) <= (!$unsigned(reg3285[(4'h9):(1'h1)]))),
                  reg3094[(2'h2):(2'h2)]};
              reg3300 <= $unsigned({$signed($unsigned(wire3074[(4'hb):(1'h1)])),
                  wire3210[(5'h17):(5'h16)],
                  $unsigned($unsigned((wire3 ? wire3 : reg3213)))});
            end
          reg3301 <= (~&($unsigned((!reg3131)) ~^ $unsigned(reg3249[(4'h8):(3'h6)])));
          reg3302 <= ($unsigned({wire3076[(5'h19):(4'hb)],
                  reg3148[(4'ha):(3'h6)]}) ?
              reg3183 : $unsigned(reg3212));
        end
      reg3303 <= (reg3142[(5'h10):(4'ha)] >= forvar3276[(2'h3):(1'h0)]);
      reg3304 = ($unsigned(((8'hba) * $unsigned($signed(reg3232)))) ?
          (^reg3168) : wire3196);
    end
  always
    @(posedge clk) begin
      reg3305 <= reg3212;
      if ($signed($signed(($signed($unsigned((8'ha3))) ?
          $unsigned($unsigned(reg3264)) : reg3149))))
        begin
          reg3306 = ((reg3299[(1'h0):(1'h0)] >>> reg3305[(5'h17):(5'h14)]) ?
              $unsigned($unsigned($unsigned($unsigned(reg3153)))) : (|$signed({(wire3198 ?
                      reg3184 : reg3101),
                  $signed(reg3133),
                  reg3163[(1'h1):(1'h0)]})));
          for (forvar3307 = (1'h0); (forvar3307 < (1'h0)); forvar3307 = (forvar3307 + (1'h1)))
            begin
              reg3308 <= $signed($unsigned($signed(wire3218[(5'h17):(5'h10)])));
              reg3309 = ($unsigned((~&reg3165[(4'hb):(4'ha)])) && (&(~&((reg3177 >> wire3197) || (~|reg3171)))));
              reg3310 = {wire3193[(4'he):(4'ha)]};
              reg3311 = $signed((wire3193 ?
                  ($unsigned($signed(reg3213)) ?
                      (&reg3115) : (!(wire3216 ?
                          reg3126 : reg3133))) : reg3146[(5'h17):(4'he)]));
            end
          if ((($unsigned(reg3249) < (($unsigned(reg3224) + (wire3196 ?
              reg3305 : reg3090)) ~^ $unsigned(reg3141))) - (((reg3291[(3'h7):(3'h4)] ^~ $unsigned((7'h42))) ?
                  (8'hb5) : ((reg3173 == reg3155) ?
                      reg3231[(2'h3):(2'h2)] : (|reg3295))) ?
              reg3115[(3'h4):(3'h4)] : (&(^~{reg3155})))))
            begin
              reg3312 <= ((!reg3265) == $signed(reg3305));
              reg3313 <= {reg3171};
            end
          else
            begin
              reg3314 = reg3269;
              reg3315 <= $signed($unsigned($unsigned(reg3231[(4'hf):(4'hc)])));
              reg3316 <= $unsigned((~^$unsigned(reg3269[(5'h15):(4'hf)])));
              reg3317 = $signed(reg3234);
              reg3318 = reg3170[(1'h0):(1'h0)];
              reg3319 <= $unsigned(reg3171[(3'h6):(3'h6)]);
              reg3320 = ((((&$unsigned(reg3133)) == (~^{reg3186,
                      reg3146,
                      reg3176})) != ($signed($unsigned(reg3170)) ?
                      (wire5[(5'h11):(4'hf)] ?
                          reg3090[(4'hc):(2'h3)] : wire3211) : $unsigned({reg3225,
                          reg3126}))) ?
                  {reg3134} : (reg3299 ?
                      ($signed((reg3257 ^ reg3280)) < reg3309) : (((reg3208 - reg3126) > {reg3299,
                          reg3184}) + reg3312)));
            end
          for (forvar3321 = (1'h0); (forvar3321 < (3'h4)); forvar3321 = (forvar3321 + (1'h1)))
            begin
              reg3322 = (reg3101 | reg3275);
              reg3323 <= reg3081;
              reg3324 = (~|$unsigned((&$signed((^reg3091)))));
              reg3325 <= $signed((reg3140[(4'h8):(3'h7)] ?
                  $signed(reg3085) : reg3264[(4'he):(3'h7)]));
            end
          for (forvar3326 = (1'h0); (forvar3326 < (1'h0)); forvar3326 = (forvar3326 + (1'h1)))
            begin
              reg3327 = reg3203;
              reg3328 <= $unsigned({(&(reg3319[(2'h2):(1'h1)] + (~^wire3076)))});
              reg3329 = $signed(reg3320[(4'hd):(1'h1)]);
              reg3330 = (reg3329 <<< wire3194);
              reg3331 = reg3167[(1'h0):(1'h0)];
            end
          reg3332 <= ((&reg3249[(1'h0):(1'h0)]) ? reg3126 : wire3078);
        end
      else
        begin
          reg3306 = {$unsigned(($unsigned((reg3264 ? reg3275 : wire3076)) ?
                  reg3146[(4'hb):(3'h4)] : (reg3300 ?
                      (wire3078 ? reg3249 : reg3186) : reg3099))),
              $unsigned(reg3328),
              $unsigned($unsigned((^reg3250[(3'h6):(2'h2)])))};
          for (forvar3307 = (1'h0); (forvar3307 < (2'h2)); forvar3307 = (forvar3307 + (1'h1)))
            begin
              reg3309 = ({($unsigned($unsigned(reg3324)) ?
                      $unsigned(reg3104[(2'h2):(2'h2)]) : (~&$unsigned((7'h42))))} <= (reg3224 ?
                  (~(~&(reg3099 == reg3284))) : $unsigned(reg3110)));
              reg3310 = ((8'hb1) ?
                  (forvar3326 ?
                      (((~&reg3319) ?
                          $signed(wire3196) : ((8'hbe) || reg3299)) >>> ((!reg3295) + $signed(reg3291))) : {{(wire3219 >>> forvar3307),
                              (8'hb6)},
                          reg3094[(2'h3):(1'h0)],
                          (~(reg3309 <<< reg3231))}) : $unsigned($unsigned(reg3284[(1'h1):(1'h1)])));
              reg3312 <= reg3087;
              reg3314 = reg3119;
            end
          reg3317 = {$signed(($unsigned(reg3141[(1'h0):(1'h0)]) * wire3211[(1'h1):(1'h0)])),
              reg3249[(4'h9):(1'h1)]};
          for (forvar3318 = (1'h0); (forvar3318 < (3'h5)); forvar3318 = (forvar3318 + (1'h1)))
            begin
              reg3320 = reg3186;
              reg3321 <= {$signed({reg3268})};
              reg3322 = $unsigned(reg3167);
              reg3323 <= reg3310[(4'h9):(2'h2)];
              reg3325 <= reg3090;
              reg3326 = wire5;
              reg3327 = (~|($unsigned((7'h55)) && (-reg3299[(5'h10):(4'h8)])));
            end
          reg3329 = (-(({(reg3225 << reg3229)} & ($signed(reg3155) + (~&reg3140))) != $unsigned($unsigned($signed((7'h40))))));
          for (forvar3330 = (1'h0); (forvar3330 < (2'h3)); forvar3330 = (forvar3330 + (1'h1)))
            begin
              reg3331 = (reg3330[(5'h12):(4'hb)] <= (reg3203[(4'hb):(3'h4)] ?
                  reg3108 : reg3213));
              reg3332 <= (!reg3332);
              reg3333 = reg3110[(1'h1):(1'h0)];
            end
          reg3334 <= (&reg3331);
        end
      reg3335 <= reg3303;
    end
  always
    @(posedge clk) begin
      reg3336 = $signed($unsigned(((-reg3171[(4'ha):(3'h6)]) ?
          reg3290[(4'h9):(3'h6)] : ((8'hbc) + (reg3165 ? (8'ha2) : reg3207)))));
      if ($signed(reg3302))
        begin
          reg3337 = {$unsigned($signed(((reg3232 && reg3135) ?
                  wire1 : reg3119))),
              (((^reg3284) == ($signed(reg3090) ?
                  (reg3332 | (8'hbf)) : reg3087)) ^ ((!(reg3237 ?
                      reg3128 : reg3177)) ?
                  (((8'hb8) - wire3210) << $unsigned((7'h50))) : ($unsigned(reg3207) ?
                      $unsigned(reg3225) : (~&reg3269))))};
          if ((reg3237[(5'h15):(4'hd)] - wire3198))
            begin
              reg3338 <= reg3090[(3'h7):(3'h4)];
              reg3339 = (|reg3203[(2'h2):(2'h2)]);
              reg3340 <= reg3313[(3'h7):(1'h0)];
              reg3341 <= $unsigned(reg3131);
              reg3342 <= (((($unsigned(reg3122) ?
                              $unsigned(reg3179) : (7'h48)) ?
                          (((7'h46) >> (8'hb8)) <<< reg3303) : reg3341) ?
                      (~|reg3275[(3'h6):(2'h2)]) : (^(reg3315 ?
                          wire1[(4'hd):(2'h3)] : (~^reg3191)))) ?
                  (~(reg3099[(2'h2):(1'h0)] ?
                      {{reg3284, wire4},
                          reg3153[(4'h8):(2'h3)]} : ((reg3319 >> reg3103) ?
                          $signed(wire3105) : (~&(8'ha9))))) : reg3340[(3'h6):(3'h5)]);
              reg3343 <= $signed({reg3286, reg3316});
              reg3344 = reg3212;
            end
          else
            begin
              reg3339 = ($unsigned(($unsigned(reg3191) ^ $signed((reg3315 ?
                  reg3188 : reg3122)))) <= $unsigned(reg3191[(4'h9):(2'h3)]));
              reg3344 = wire3211[(3'h7):(2'h3)];
              reg3345 <= reg3321[(1'h1):(1'h1)];
              reg3346 <= ($unsigned((reg3266 ?
                  ($unsigned(reg3156) <<< ((7'h55) ?
                      wire3198 : (8'ha4))) : reg3259[(1'h1):(1'h0)])) >>> $unsigned($signed($signed(wire3078[(5'h10):(4'hf)]))));
              reg3347 = ({reg3296[(1'h0):(1'h0)],
                  $signed(($unsigned(reg3135) ? (~reg3108) : $signed(reg3094))),
                  wire3219[(1'h1):(1'h1)]} << $signed($unsigned($signed(wire3194))));
              reg3348 = (wire3193[(5'h1a):(5'h10)] ?
                  reg3126 : ((~&reg3149) ?
                      ((reg3128 ?
                          (reg3332 & wire3073) : reg3280) == (^~wire3196)) : (+(8'hb2))));
              reg3349 <= $signed(wire3074);
            end
          if (($unsigned(((~^wire3105[(4'h9):(2'h3)]) < $unsigned((reg3290 ?
                  reg3149 : wire3)))) ?
              reg3295[(3'h5):(1'h1)] : wire3194))
            begin
              reg3350 = (!$signed(wire3210));
              reg3351 = (((~|(8'ha0)) ^~ reg3244[(4'hf):(1'h1)]) ?
                  $signed($unsigned(((reg3303 | reg3247) ?
                      reg3087 : $unsigned(reg3313)))) : (&reg3319));
              reg3352 <= reg3080[(5'h18):(5'h10)];
            end
          else
            begin
              reg3350 = ((((8'ha5) <= reg3340[(5'h11):(3'h4)]) && (~(reg3171[(4'h9):(3'h4)] ^~ (reg3249 ?
                  reg3101 : wire3211)))) == reg3100);
              reg3351 = $unsigned($unsigned(reg3128));
            end
        end
      else
        begin
          reg3337 = $signed(({reg3081[(4'ha):(2'h3)],
                  $signed($unsigned(reg3171))} ?
              ($unsigned((reg3177 ^ reg3325)) ~^ reg3085[(2'h2):(2'h2)]) : reg3292));
          reg3339 = wire3210[(5'h13):(5'h10)];
        end
    end
  module1773 #() modinst3354 (.clk(clk), .wire1774(reg3104), .wire1775(reg3308), .wire1777(reg3234), .y(wire3353), .wire1776(reg3349), .wire1778(reg3247));
  always
    @(posedge clk) begin
      reg3355 = $signed(reg3085[(4'hf):(4'h8)]);
    end
  module326 #() modinst3357 (.wire329(reg3108), .wire330(reg3302), .wire331(wire3074), .clk(clk), .y(wire3356), .wire328(reg3280), .wire327(reg3283));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module6  (y, clk, wire7, wire8, wire9, wire10);
  output wire [(32'h936):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire7;
  input wire signed [(5'h1a):(1'h0)] wire8;
  input wire [(5'h17):(1'h0)] wire9;
  input wire signed [(3'h7):(1'h0)] wire10;
  wire [(3'h4):(1'h0)] wire69;
  wire [(5'h1a):(1'h0)] wire70;
  wire [(5'h1b):(1'h0)] wire844;
  wire [(5'h1f):(1'h0)] wire3069;
  reg [(4'hf):(1'h0)] reg919 = (1'h0);
  reg [(3'h6):(1'h0)] reg915 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg914 = (1'h0);
  reg [(4'hd):(1'h0)] reg913 = (1'h0);
  reg [(5'h15):(1'h0)] reg912 = (1'h0);
  reg [(4'hb):(1'h0)] reg911 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg909 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg906 = (1'h0);
  reg [(5'h1d):(1'h0)] reg905 = (1'h0);
  reg [(5'h16):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg903 = (1'h0);
  reg [(4'hc):(1'h0)] reg897 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg894 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg890 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg889 = (1'h0);
  reg [(4'hb):(1'h0)] reg888 = (1'h0);
  reg [(5'h14):(1'h0)] reg887 = (1'h0);
  reg [(5'h1c):(1'h0)] reg886 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg885 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg883 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg882 = (1'h0);
  reg [(4'h8):(1'h0)] reg880 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg879 = (1'h0);
  reg [(4'hc):(1'h0)] reg875 = (1'h0);
  reg [(2'h2):(1'h0)] reg874 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg872 = (1'h0);
  reg [(5'h16):(1'h0)] reg869 = (1'h0);
  reg [(5'h13):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg866 = (1'h0);
  reg [(3'h6):(1'h0)] reg864 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg861 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg860 = (1'h0);
  reg [(2'h2):(1'h0)] reg858 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg854 = (1'h0);
  reg [(5'h18):(1'h0)] reg853 = (1'h0);
  reg [(5'h17):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg62 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg61 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg55 = (1'h0);
  reg [(5'h1b):(1'h0)] reg54 = (1'h0);
  reg [(5'h13):(1'h0)] reg53 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg52 = (1'h0);
  reg [(5'h16):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg49 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg48 = (1'h0);
  reg [(5'h17):(1'h0)] reg46 = (1'h0);
  reg [(4'h9):(1'h0)] reg45 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg41 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg39 = (1'h0);
  reg [(3'h5):(1'h0)] reg34 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg30 = (1'h0);
  reg [(4'hc):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg21 = (1'h0);
  reg [(3'h7):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg18 = (1'h0);
  reg [(5'h14):(1'h0)] reg13 = (1'h0);
  reg [(4'hf):(1'h0)] reg12 = (1'h0);
  reg [(5'h11):(1'h0)] reg11 = (1'h0);
  reg [(5'h12):(1'h0)] reg922 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg921 = (1'h0);
  reg [(3'h4):(1'h0)] reg920 = (1'h0);
  reg [(5'h14):(1'h0)] reg918 = (1'h0);
  reg [(5'h14):(1'h0)] reg917 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar916 = (1'h0);
  reg [(4'hc):(1'h0)] reg910 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar908 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg907 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg902 = (1'h0);
  reg [(4'h9):(1'h0)] reg901 = (1'h0);
  reg [(4'hd):(1'h0)] reg900 = (1'h0);
  reg [(5'h17):(1'h0)] forvar899 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg898 = (1'h0);
  reg [(2'h3):(1'h0)] reg896 = (1'h0);
  reg [(5'h13):(1'h0)] reg893 = (1'h0);
  reg [(5'h19):(1'h0)] reg892 = (1'h0);
  reg [(5'h1c):(1'h0)] reg891 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar884 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg881 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg870 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar868 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg878 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg877 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg876 = (1'h0);
  reg [(4'hb):(1'h0)] reg873 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg871 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar870 = (1'h0);
  reg [(5'h19):(1'h0)] reg867 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar865 = (1'h0);
  reg [(5'h14):(1'h0)] reg863 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg862 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg859 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg857 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg856 = (1'h0);
  reg [(5'h1e):(1'h0)] reg855 = (1'h0);
  reg [(3'h5):(1'h0)] forvar852 = (1'h0);
  reg [(5'h16):(1'h0)] reg850 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg849 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar848 = (1'h0);
  reg [(5'h13):(1'h0)] reg847 = (1'h0);
  reg [(5'h1c):(1'h0)] reg846 = (1'h0);
  reg [(5'h1b):(1'h0)] reg68 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg66 = (1'h0);
  reg [(5'h14):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg63 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg59 = (1'h0);
  reg [(5'h17):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg47 = (1'h0);
  reg [(3'h6):(1'h0)] forvar44 = (1'h0);
  reg [(3'h5):(1'h0)] reg43 = (1'h0);
  reg [(4'hb):(1'h0)] reg42 = (1'h0);
  reg [(4'ha):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg38 = (1'h0);
  reg [(5'h10):(1'h0)] reg37 = (1'h0);
  reg [(5'h17):(1'h0)] reg36 = (1'h0);
  reg [(2'h3):(1'h0)] reg35 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar33 = (1'h0);
  reg [(4'hb):(1'h0)] forvar31 = (1'h0);
  reg [(5'h10):(1'h0)] reg28 = (1'h0);
  reg [(3'h6):(1'h0)] reg27 = (1'h0);
  reg [(5'h1e):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg24 = (1'h0);
  reg [(4'hd):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg19 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar15 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg14 = (1'h0);
  assign y = {wire69,
                 wire70,
                 wire844,
                 wire3069,
                 reg919,
                 reg915,
                 reg914,
                 reg913,
                 reg912,
                 reg911,
                 reg909,
                 reg906,
                 reg905,
                 reg904,
                 reg903,
                 reg897,
                 reg895,
                 reg894,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 reg886,
                 reg885,
                 reg883,
                 reg882,
                 reg880,
                 reg879,
                 reg875,
                 reg874,
                 reg872,
                 reg869,
                 reg868,
                 reg866,
                 reg864,
                 reg861,
                 reg860,
                 reg858,
                 reg854,
                 reg853,
                 reg851,
                 reg67,
                 reg62,
                 reg61,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg49,
                 reg48,
                 reg46,
                 reg45,
                 reg41,
                 reg39,
                 reg34,
                 reg32,
                 reg30,
                 reg29,
                 reg26,
                 reg23,
                 reg21,
                 reg20,
                 reg18,
                 reg13,
                 reg12,
                 reg11,
                 reg922,
                 reg921,
                 reg920,
                 reg918,
                 reg917,
                 forvar916,
                 reg910,
                 forvar908,
                 reg907,
                 reg902,
                 reg901,
                 reg900,
                 forvar899,
                 reg898,
                 reg896,
                 reg893,
                 reg892,
                 reg891,
                 forvar884,
                 reg881,
                 reg870,
                 forvar868,
                 reg878,
                 reg877,
                 reg876,
                 reg873,
                 reg871,
                 forvar870,
                 reg867,
                 forvar865,
                 reg863,
                 reg862,
                 reg859,
                 reg857,
                 reg856,
                 reg855,
                 forvar852,
                 reg850,
                 reg849,
                 forvar848,
                 reg847,
                 reg846,
                 reg68,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg50,
                 reg47,
                 forvar44,
                 reg43,
                 reg42,
                 reg40,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 forvar33,
                 forvar31,
                 reg28,
                 reg27,
                 reg25,
                 reg24,
                 reg22,
                 reg19,
                 reg17,
                 reg16,
                 forvar15,
                 reg14,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg11 <= ((~&$unsigned(($unsigned(wire7) == wire10))) ^~ ($signed((~|$signed(wire10))) && (~|($unsigned(wire8) ?
          $unsigned(wire10) : $signed(wire10)))));
      reg12 <= (({$unsigned((wire9 ? (7'h55) : wire7)),
                  (wire10 | (wire8 ? wire9 : wire8))} ?
              ($signed((wire8 ? wire8 : wire9)) >> (^{reg11})) : reg11) ?
          (wire10[(1'h1):(1'h1)] * (~&$unsigned({(8'hac),
              wire10}))) : $unsigned((wire9[(4'hc):(1'h1)] ?
              $unsigned(wire10[(3'h5):(3'h4)]) : (wire8 ?
                  wire8 : (reg11 ^~ wire9)))));
      reg13 <= {(~|wire8)};
      reg14 = (^$signed($signed($unsigned((reg12 ? wire7 : wire7)))));
      if ((^(-(&(wire10[(3'h4):(2'h3)] || $signed(wire7))))))
        begin
          for (forvar15 = (1'h0); (forvar15 < (1'h0)); forvar15 = (forvar15 + (1'h1)))
            begin
              reg16 = wire7[(4'hd):(3'h7)];
              reg17 = $signed(reg11[(5'h10):(5'h10)]);
              reg18 <= $signed($signed({($unsigned(reg16) ?
                      (reg16 != reg14) : (wire9 || reg16)),
                  (wire8[(5'h18):(3'h5)] ?
                      (reg16 ? reg12 : reg12) : reg14[(3'h7):(3'h6)])}));
              reg19 = $unsigned(((wire8 ?
                  reg14 : reg13[(4'hb):(4'h9)]) == $unsigned($signed(wire9))));
              reg20 <= ($unsigned(((reg16[(3'h4):(2'h3)] < reg18[(2'h3):(1'h0)]) ?
                      $signed($unsigned(wire10)) : ((wire10 ?
                          wire7 : reg13) >>> (~^reg12)))) ?
                  wire10 : reg17);
              reg21 <= reg20[(3'h4):(2'h2)];
            end
          if (($unsigned(wire9[(3'h5):(1'h0)]) ?
              ((-$signed($unsigned(reg16))) ^ (reg20 ?
                  reg12 : $signed((reg16 != reg12)))) : wire7))
            begin
              reg22 = reg17[(4'ha):(3'h5)];
              reg23 <= reg13[(3'h6):(2'h3)];
              reg24 = $unsigned($signed(reg17[(4'h8):(2'h3)]));
              reg25 = (7'h55);
              reg26 <= ((&({$unsigned(reg23),
                      {reg12},
                      (wire7 ? reg16 : (7'h54))} ?
                  reg22[(3'h4):(1'h1)] : ((reg13 ?
                      reg19 : reg19) ^~ (|reg24)))) || (!$signed($signed(((7'h53) + reg16)))));
              reg27 = (((reg16[(2'h2):(1'h1)] ^ reg16[(1'h1):(1'h0)]) ?
                  (-({reg18, (8'hb8), reg20} ?
                      (!reg12) : {reg21,
                          (8'ha0)})) : $signed(reg13)) >>> ((7'h43) ?
                  ((+reg21[(1'h0):(1'h0)]) ?
                      forvar15[(4'hc):(1'h1)] : $signed(reg25[(5'h1b):(5'h18)])) : forvar15[(4'hd):(4'hc)]));
              reg28 = (reg11 ?
                  reg12 : $signed((&($unsigned(wire9) ?
                      reg12[(1'h0):(1'h0)] : (wire9 ? (8'hbe) : reg16)))));
            end
          else
            begin
              reg22 = $signed(reg23);
              reg24 = ((wire7[(4'h9):(3'h4)] >> ($unsigned((reg13 ?
                  reg21 : reg11)) > (^(~&(8'haa))))) >= $unsigned((^{reg11[(3'h7):(3'h7)],
                  reg17})));
              reg26 <= $unsigned($unsigned($unsigned((wire7[(3'h4):(3'h4)] == forvar15[(4'hc):(4'ha)]))));
              reg29 <= reg26[(1'h0):(1'h0)];
              reg30 <= (+$unsigned(wire8));
            end
          for (forvar31 = (1'h0); (forvar31 < (3'h6)); forvar31 = (forvar31 + (1'h1)))
            begin
              reg32 <= {((^$signed((reg28 - (7'h40)))) ?
                      wire7[(4'h8):(1'h1)] : (~(~^{reg27}))),
                  ($signed(((-forvar15) << $unsigned(reg18))) ?
                      reg21[(4'hf):(2'h3)] : reg29[(4'ha):(4'h8)]),
                  reg30[(4'he):(2'h2)]};
            end
          for (forvar33 = (1'h0); (forvar33 < (1'h1)); forvar33 = (forvar33 + (1'h1)))
            begin
              reg34 <= (~&forvar33[(4'he):(3'h7)]);
              reg35 = forvar31;
            end
          if ((({(&reg11[(4'h8):(3'h5)])} <= (|(+reg27[(3'h4):(2'h2)]))) ?
              $unsigned($signed((+wire9))) : $unsigned($signed(({reg11,
                  reg19,
                  (8'ha7)} <<< {reg25})))))
            begin
              reg36 = forvar15;
              reg37 = (!(~wire10));
              reg38 = {reg12, (~reg36), reg17[(4'hc):(3'h7)]};
              reg39 <= $signed((reg27[(2'h3):(2'h3)] <<< reg25[(5'h10):(4'hd)]));
              reg40 = (7'h4e);
            end
          else
            begin
              reg36 = {forvar33};
              reg39 <= reg22;
              reg40 = ({($unsigned((reg23 < wire9)) ?
                          (~&$signed(wire10)) : {$unsigned(reg28)}),
                      reg18[(2'h2):(1'h0)],
                      (-($unsigned(reg22) <<< (7'h45)))} ?
                  $unsigned({(^$signed(reg40))}) : reg11);
              reg41 <= {wire10[(2'h2):(1'h0)],
                  ($signed(reg18[(2'h2):(1'h1)]) && ((~^$signed(reg12)) ?
                      reg19 : $unsigned((wire9 ~^ reg17)))),
                  $signed(reg18[(2'h2):(1'h1)])};
              reg42 = (($signed((+{reg35, wire7, (7'h48)})) ?
                  {reg35} : (forvar15[(4'hf):(1'h1)] ~^ $unsigned(reg14[(3'h6):(3'h5)]))) <= $unsigned(wire9));
              reg43 = forvar33;
            end
        end
      else
        begin
          for (forvar15 = (1'h0); (forvar15 < (3'h6)); forvar15 = (forvar15 + (1'h1)))
            begin
              reg18 <= reg43;
              reg20 <= $unsigned(reg26);
              reg21 <= $signed($signed(reg28[(3'h5):(3'h4)]));
            end
          reg23 <= $unsigned($unsigned($unsigned((^(^forvar15)))));
          reg26 <= reg32[(4'h9):(3'h4)];
        end
      for (forvar44 = (1'h0); (forvar44 < (3'h4)); forvar44 = (forvar44 + (1'h1)))
        begin
          if ($unsigned(reg32[(4'h8):(2'h2)]))
            begin
              reg45 <= (((^~$signed($signed(forvar15))) >>> $unsigned(((reg19 < reg37) >> wire8[(5'h12):(1'h0)]))) ?
                  (!$signed((~|(~|(7'h42))))) : (&$signed(((reg25 || reg28) ?
                      (reg19 ? reg29 : reg37) : (reg37 >> (8'hb5))))));
              reg46 <= ({(7'h51),
                      reg12[(1'h0):(1'h0)],
                      $unsigned(reg37[(4'he):(4'hd)])} ?
                  $unsigned($unsigned({(reg19 ? reg36 : reg14),
                      reg30[(5'h1c):(5'h19)]})) : {($signed((reg11 ?
                          reg16 : wire10)) | wire9),
                      (+($unsigned(reg12) ~^ reg43[(1'h1):(1'h0)]))});
              reg47 = (^~{((reg20[(3'h6):(1'h0)] <<< (reg39 ? reg22 : reg38)) ?
                      $unsigned(forvar33[(1'h0):(1'h0)]) : (&(|forvar15)))});
              reg48 <= $signed($signed((!forvar44[(1'h1):(1'h0)])));
              reg49 <= reg24;
            end
          else
            begin
              reg47 = ($unsigned({{$signed((8'hbf)),
                          {reg28, reg48, reg16},
                          ((8'haf) ^~ reg28)}}) ?
                  ((|reg20) ?
                      $unsigned(({reg43,
                          reg29,
                          (7'h46)} <= $unsigned(reg48))) : reg39[(2'h3):(1'h0)]) : (reg35[(2'h3):(2'h3)] ?
                      wire10[(3'h5):(3'h4)] : {reg22,
                          ((reg29 ? reg16 : (8'haf)) ?
                              (forvar33 ? reg48 : reg28) : (reg12 < reg19)),
                          (reg12 ? $unsigned(wire7) : $signed(reg25))}));
              reg48 <= ((reg34 >= reg34[(2'h3):(1'h1)]) ?
                  $signed(reg17[(4'h8):(3'h7)]) : reg48[(4'h8):(2'h3)]);
              reg49 <= (reg40[(4'h8):(3'h4)] ?
                  (({(reg20 ? (7'h43) : reg36), reg23} << ((reg22 && reg28) ?
                      reg30[(3'h6):(2'h2)] : forvar44[(3'h4):(2'h2)])) >> reg42[(3'h6):(3'h5)]) : ($unsigned({wire8}) << reg37));
              reg50 = {$signed(reg18), wire9[(5'h16):(4'h8)]};
              reg51 <= ($unsigned(($signed(reg40) ?
                  {$signed(wire9),
                      forvar15} : $unsigned($unsigned((7'h50))))) >>> $unsigned($signed((8'hab))));
              reg52 <= $signed(($unsigned(reg45) ?
                  $signed(($signed(reg27) ?
                      $unsigned(reg26) : (reg38 ?
                          (7'h51) : (7'h47)))) : (~|(reg34 < $unsigned(reg30)))));
              reg53 <= $unsigned($unsigned(reg34[(2'h2):(2'h2)]));
            end
          if ($signed(((&((reg30 >= (7'h45)) + (8'haf))) ?
              reg43[(2'h3):(1'h1)] : ((^reg22[(4'h8):(4'h8)]) >= {{reg35},
                  (reg21 ? reg32 : (8'h9c))}))))
            begin
              reg54 <= ($signed((reg23 >= $signed($unsigned((7'h49))))) ?
                  {$unsigned(reg45), reg32[(4'h9):(2'h2)]} : reg34);
              reg55 <= $unsigned(((((7'h53) ? {reg37, reg41, reg27} : reg25) ?
                  (~|$signed(reg42)) : (!$signed(reg30))) == $signed((8'h9d))));
              reg56 <= {($unsigned(reg30[(4'hd):(2'h2)]) == (reg28 - ($unsigned(reg23) ?
                      (reg40 ? reg29 : reg35) : (^forvar15))))};
              reg57 = reg47;
              reg58 = (|(reg30 >> (~^$signed((reg42 ? wire8 : reg35)))));
            end
          else
            begin
              reg54 <= ($signed(reg29[(4'h9):(4'h8)]) - reg14);
            end
          if (($signed((&((!wire7) ?
              $signed(reg53) : $signed((7'h53))))) >> (reg18 ?
              (^~$unsigned((-reg41))) : $signed($signed(reg30[(1'h0):(1'h0)])))))
            begin
              reg59 = (&(~^reg18));
            end
          else
            begin
              reg59 = ($signed($unsigned(($unsigned(reg29) ?
                      (~&reg14) : (reg19 ? reg45 : reg53)))) ?
                  $unsigned((~^(wire9 | reg43))) : ({$unsigned({(8'hab),
                          reg28}),
                      {$signed((8'ha9)),
                          $signed(reg13)}} ^~ (($unsigned((8'hba)) ?
                          reg38 : (wire10 ? forvar31 : reg55)) ?
                      $unsigned(wire9[(4'hf):(4'he)]) : reg21)));
            end
          reg60 = (~&({reg47[(4'ha):(1'h0)],
              (wire7 ? reg47 : (-forvar33))} <<< (~&(-reg29[(4'hc):(4'hc)]))));
          if (((^({$unsigned(reg41)} ?
              {$signed((7'h45)), (~|reg46)} : ({reg16} ?
                  (+reg42) : (-reg35)))) ~^ $unsigned(reg58)))
            begin
              reg61 <= reg12[(1'h1):(1'h1)];
              reg62 <= $signed({($unsigned(forvar15[(3'h6):(1'h1)]) || forvar15)});
              reg63 = reg18;
              reg64 = forvar33;
              reg65 = $unsigned($unsigned((^$unsigned(reg38))));
              reg66 = $signed(reg19);
            end
          else
            begin
              reg63 = reg37[(2'h2):(1'h0)];
              reg64 = {{{((~|wire7) * (~reg46))},
                      (reg30 ? reg21 : (^reg37[(3'h7):(2'h3)])),
                      $signed({forvar44})},
                  (~|($signed(reg25) ?
                      {{reg23},
                          forvar33,
                          {reg37, forvar15}} : $unsigned((~&reg19))))};
              reg67 <= (~|((($signed(reg41) ? (~^reg52) : (&reg14)) ?
                  ((reg25 + reg20) << $unsigned(reg20)) : ((reg24 ?
                          reg26 : reg62) ?
                      ((8'hbe) ?
                          (7'h56) : reg35) : ((8'hbe) != reg37))) + reg21));
            end
          reg68 = reg48;
        end
    end
  assign wire69 = (({{$signed(reg52), $unsigned(reg13), reg54[(4'hd):(3'h6)]},
                              ((reg32 <= wire10) ? $signed(reg20) : (7'h46))} ?
                          reg55 : ($unsigned((reg23 ? reg12 : reg53)) ?
                              {(^~reg67),
                                  $signed(reg26)} : $signed($signed(reg54)))) ?
                      (((-reg23[(3'h7):(1'h0)]) ?
                          ((reg12 <= reg12) ?
                              {reg61} : (reg49 ?
                                  reg51 : reg13)) : $signed((~(8'hb2)))) & $signed($unsigned(wire7))) : (7'h53));
  assign wire70 = $unsigned((({((7'h49) | (7'h4c)), (reg52 && (7'h52))} ?
                      ((8'hac) == (reg30 ?
                          (7'h4f) : (8'h9c))) : (|reg11[(4'he):(3'h4)])) ~^ reg29[(4'hc):(1'h0)]));
  module71 #() modinst845 (wire844, clk, reg18, reg48, reg12, reg26, reg29, reg11);
  always
    @(posedge clk) begin
      if ((reg41[(4'h9):(1'h0)] ?
          reg11[(4'hd):(3'h4)] : $unsigned($signed(({(7'h51)} << (reg39 && reg48))))))
        begin
          reg846 = {$signed($unsigned($signed(reg29))),
              ({(reg52 ? $unsigned(reg18) : $signed(wire8)),
                      (reg52[(3'h5):(3'h4)] && $unsigned(reg48)),
                      ((reg48 ? reg18 : reg41) * (reg53 ~^ (7'h52)))} ?
                  $unsigned($signed(wire9[(4'hf):(4'hf)])) : {$signed($signed(reg56)),
                      $signed($unsigned(reg23)),
                      (!(^~reg45))}),
              ($signed(reg30) ?
                  $unsigned((reg11 ? reg26 : $signed(reg46))) : reg11)};
        end
      else
        begin
          reg846 = {$unsigned($unsigned((~$unsigned((7'h4d))))),
              (|reg62),
              $unsigned(reg13[(5'h12):(2'h3)])};
          reg847 = (reg13 ?
              $signed(((reg48 - reg29) >= {$unsigned(reg51)})) : ((($unsigned((8'ha7)) ^~ (^reg48)) && $unsigned((wire10 & reg26))) >> ((reg45 ?
                  $unsigned((7'h4c)) : $signed((8'ha0))) ^~ (^~reg32))));
          for (forvar848 = (1'h0); (forvar848 < (1'h0)); forvar848 = (forvar848 + (1'h1)))
            begin
              reg849 = (((|(^$unsigned(reg29))) ?
                  (!reg39) : ($signed($signed(reg29)) <<< (~|{forvar848,
                      (8'ha6)}))) ^~ wire69[(3'h4):(2'h3)]);
              reg850 = reg26[(1'h0):(1'h0)];
              reg851 <= (+$signed(reg49[(3'h4):(2'h2)]));
            end
          for (forvar852 = (1'h0); (forvar852 < (2'h2)); forvar852 = (forvar852 + (1'h1)))
            begin
              reg853 <= $signed(wire69[(3'h4):(3'h4)]);
              reg854 <= $unsigned((-$signed($signed($signed((8'hbc))))));
              reg855 = reg853[(2'h3):(2'h3)];
              reg856 = (!($signed(reg54[(2'h2):(2'h2)]) ?
                  (~reg847) : (^reg851)));
              reg857 = ((~&$unsigned(reg39[(1'h1):(1'h1)])) && wire69);
              reg858 <= {(8'hb6),
                  $signed(($unsigned($signed(reg853)) ?
                      ($unsigned(reg29) ^~ $unsigned(reg26)) : (wire9 ^ {wire9}))),
                  reg55};
            end
          if ((!($unsigned(reg46[(5'h12):(5'h12)]) >> {(|reg851[(4'ha):(3'h6)]),
              $unsigned($signed(reg855))})))
            begin
              reg859 = ((^~$unsigned($signed($signed((7'h55))))) ?
                  $unsigned($signed((-$signed(reg851)))) : $signed({(!(reg45 ?
                          reg847 : reg847)),
                      {reg39[(1'h0):(1'h0)], (reg67 ? (7'h46) : reg41)}}));
              reg860 <= $unsigned(reg34);
              reg861 <= reg46;
              reg862 = $unsigned(wire8);
              reg863 = {(8'ha4)};
              reg864 <= reg34[(2'h2):(2'h2)];
            end
          else
            begin
              reg860 <= (reg20[(3'h5):(1'h1)] ?
                  (((reg30[(3'h6):(1'h0)] != $signed(reg23)) ?
                          $unsigned((~&reg861)) : (|((7'h48) ?
                              reg29 : forvar852))) ?
                      $unsigned($unsigned(reg21[(3'h5):(3'h5)])) : (7'h4f)) : reg851);
              reg862 = $unsigned((reg54 ?
                  ((reg39 ? (reg855 ? reg856 : reg51) : $signed(reg861)) ?
                      $unsigned($signed(reg859)) : reg854) : {($signed(wire69) | (8'ha9))}));
              reg864 <= $signed(reg863);
            end
          for (forvar865 = (1'h0); (forvar865 < (2'h2)); forvar865 = (forvar865 + (1'h1)))
            begin
              reg866 <= (!wire70[(3'h7):(1'h0)]);
            end
          reg867 = $unsigned(reg862[(4'h9):(4'h8)]);
        end
      if (reg855)
        begin
          reg868 <= $unsigned(($signed(reg867) && (8'ha7)));
          reg869 <= reg56;
          for (forvar870 = (1'h0); (forvar870 < (1'h1)); forvar870 = (forvar870 + (1'h1)))
            begin
              reg871 = $signed(reg26[(4'hd):(2'h2)]);
            end
          reg872 <= (wire9 < (~|reg850));
          if ($unsigned($unsigned((8'hab))))
            begin
              reg873 = $signed(reg54[(5'h19):(5'h16)]);
              reg874 <= ($signed({(forvar852[(1'h1):(1'h1)] > reg869),
                      {reg847, wire10},
                      (^$unsigned((8'hb1)))}) ?
                  (~$unsigned((^~{reg11}))) : ($unsigned($signed(reg846[(3'h7):(1'h0)])) ~^ (^{(wire70 ?
                          reg868 : reg853)})));
              reg875 <= reg858[(1'h1):(1'h0)];
              reg876 = {(reg856[(1'h1):(1'h0)] == ((|reg846[(4'h8):(3'h7)]) ?
                      reg863 : wire9[(2'h3):(2'h2)])),
                  reg866,
                  ((~^$unsigned(reg11)) ?
                      $unsigned((-$signed((8'hb6)))) : reg858[(2'h2):(1'h1)])};
              reg877 = reg39[(1'h0):(1'h0)];
              reg878 = ((reg861 ?
                  (reg846[(5'h12):(5'h12)] >>> {reg863,
                      (reg853 <<< reg48),
                      reg53[(3'h4):(2'h3)]}) : reg859) > {(wire8 ?
                      (^wire10) : (reg12[(4'he):(2'h2)] <<< ((8'haa) ?
                          wire9 : reg13))),
                  wire8[(1'h0):(1'h0)]});
            end
          else
            begin
              reg874 <= ((reg855[(5'h12):(5'h11)] ?
                      {reg62} : $unsigned(($signed(reg51) != $signed(reg61)))) ?
                  wire10[(1'h0):(1'h0)] : reg846);
              reg876 = reg23;
              reg879 <= reg862;
            end
        end
      else
        begin
          for (forvar868 = (1'h0); (forvar868 < (1'h1)); forvar868 = (forvar868 + (1'h1)))
            begin
              reg870 = (7'h4c);
              reg872 <= forvar865[(1'h0):(1'h0)];
            end
          if (reg860)
            begin
              reg874 <= reg12[(2'h3):(2'h2)];
              reg875 <= $unsigned($unsigned(reg18[(4'hc):(1'h1)]));
              reg879 <= (-(($signed(wire10) != $unsigned(((8'h9d) || reg846))) | (~&$signed($signed((7'h41))))));
              reg880 <= ((((-wire9[(4'hf):(4'ha)]) <= wire10[(3'h6):(3'h6)]) ?
                      ($signed(wire70[(5'h16):(4'he)]) || wire7) : reg30[(4'h8):(1'h1)]) ?
                  ($signed((^$unsigned(reg847))) + reg56[(4'ha):(2'h2)]) : reg868[(1'h1):(1'h1)]);
              reg881 = wire9[(5'h11):(3'h5)];
              reg882 <= $unsigned({(reg860 ?
                      (^(reg13 ? (8'hb9) : reg39)) : {reg864,
                          (reg32 || reg18)}),
                  {((reg867 ? reg876 : wire844) ?
                          $unsigned(reg875) : {(8'hab)})},
                  (7'h4e)});
              reg883 <= (|$signed(((reg48 + reg872[(5'h11):(4'ha)]) ?
                  $unsigned(reg20[(1'h0):(1'h0)]) : ((7'h4c) >>> (reg61 + reg46)))));
            end
          else
            begin
              reg873 = forvar848[(1'h1):(1'h0)];
              reg876 = $unsigned({{reg26[(5'h10):(2'h2)],
                      $unsigned($signed(reg52))},
                  (reg51[(3'h4):(2'h3)] ?
                      ($unsigned(wire9) ?
                          $unsigned(reg849) : reg18[(4'hf):(4'ha)]) : $signed((reg23 ?
                          reg51 : reg56))),
                  $unsigned((reg39[(2'h2):(1'h0)] ^ (reg860 ?
                      reg878 : forvar870)))});
              reg879 <= {(+$unsigned($unsigned((reg866 - reg876)))),
                  (+$signed(forvar868[(3'h7):(3'h5)]))};
            end
          for (forvar884 = (1'h0); (forvar884 < (3'h4)); forvar884 = (forvar884 + (1'h1)))
            begin
              reg885 <= reg48[(4'h9):(4'h9)];
              reg886 <= $unsigned((^~{(^~$unsigned((7'h4d)))}));
              reg887 <= $signed(reg32);
              reg888 <= $signed(((+reg859[(2'h3):(1'h1)]) >>> (~&(8'h9f))));
              reg889 <= $unsigned(reg52);
              reg890 <= $unsigned($signed($signed(reg867[(2'h3):(1'h0)])));
              reg891 = {(8'hbc)};
            end
          if ({reg61})
            begin
              reg892 = (|$signed((reg49[(3'h4):(2'h3)] <<< $signed({wire10}))));
              reg893 = (reg890 ?
                  reg868 : $unsigned($signed($unsigned((+forvar868)))));
              reg894 <= ((^$unsigned($signed($signed((8'h9d))))) ?
                  ({$signed((reg861 << reg62)),
                      (~$signed(reg850)),
                      $unsigned(reg49[(3'h4):(1'h0)])} ~^ $unsigned(reg862[(3'h5):(3'h4)])) : (-{$signed($signed((8'hbf))),
                      reg875[(3'h5):(2'h3)]}));
              reg895 <= (~reg11);
              reg896 = (((^(&(~forvar884))) ?
                  (&(~reg850[(5'h16):(2'h2)])) : $signed(forvar884[(3'h5):(3'h4)])) + (((^~(reg23 ?
                      (8'ha5) : forvar848)) || ($unsigned((8'hb3)) < {reg887,
                      reg30})) ?
                  ((~&$unsigned(reg56)) ?
                      (^$unsigned(reg39)) : $unsigned((reg892 != reg859))) : (~^reg870[(3'h4):(1'h0)])));
              reg897 <= {(8'h9f), $signed(reg889[(5'h17):(4'hf)])};
            end
          else
            begin
              reg892 = reg880;
              reg893 = $unsigned({(^reg850[(5'h15):(5'h14)]),
                  reg23[(5'h16):(4'h8)],
                  ($signed((reg896 ? reg867 : reg895)) <= $unsigned(reg23))});
            end
          reg898 = $unsigned({{$unsigned($unsigned(reg886))}});
        end
      for (forvar899 = (1'h0); (forvar899 < (2'h3)); forvar899 = (forvar899 + (1'h1)))
        begin
          reg900 = (~^reg32);
          if (reg879[(3'h6):(3'h6)])
            begin
              reg901 = (($unsigned(((wire9 ? reg29 : reg853) && (~^reg846))) ?
                  $signed(reg51[(4'ha):(4'h9)]) : $signed($unsigned(((8'ha8) ?
                      reg860 : reg45)))) && reg874);
              reg902 = $unsigned($signed({$signed($signed((7'h4e))),
                  ((reg866 >= reg67) ? reg856 : $unsigned((7'h4b))),
                  ($unsigned(reg874) ~^ reg885)}));
              reg903 <= $unsigned((!(reg890[(1'h0):(1'h0)] ?
                  reg39[(1'h1):(1'h1)] : ($unsigned(reg878) ?
                      $signed(wire9) : $signed(reg29)))));
              reg904 <= reg29;
            end
          else
            begin
              reg901 = (~&(~{$unsigned({reg866, reg13}),
                  $unsigned($signed(reg871)),
                  forvar848[(2'h3):(2'h3)]}));
              reg902 = {(reg886 >= $unsigned(reg881[(5'h13):(5'h12)])),
                  ((((~^reg877) ? $signed(reg892) : reg56[(3'h4):(1'h0)]) ?
                          reg885 : ((reg903 ? reg863 : (7'h43)) ?
                              (&(8'ha7)) : (reg21 ? forvar868 : reg895))) ?
                      reg876 : reg850[(1'h1):(1'h1)])};
            end
          reg905 <= {(~&(|forvar868)),
              $signed({((reg850 || (8'ha5)) != {(8'ha2), reg904}),
                  ({forvar865, reg55, reg873} && (reg55 ? reg863 : reg857))}),
              ((forvar848 - {{reg904, reg860}, (reg52 ? reg903 : wire844)}) ?
                  $unsigned((((7'h44) ? wire7 : reg61) ?
                      $signed(reg882) : ((8'ha6) ?
                          reg871 : forvar868))) : reg857[(3'h5):(2'h2)])};
          if ($unsigned(((7'h40) ?
              (~&(+(!reg874))) : ((!forvar899) <= reg851[(4'hb):(1'h1)]))))
            begin
              reg906 <= reg864;
              reg907 = (!((8'ha0) != reg856));
            end
          else
            begin
              reg907 = $signed(($unsigned(reg867[(4'hd):(1'h0)]) << {$signed(reg54[(5'h1a):(3'h5)]),
                  $signed($signed((8'ha7))),
                  (((7'h57) ? reg18 : reg13) ?
                      reg846[(5'h15):(1'h0)] : (~|(8'ha9)))}));
            end
          for (forvar908 = (1'h0); (forvar908 < (3'h6)); forvar908 = (forvar908 + (1'h1)))
            begin
              reg909 <= $unsigned((reg904[(1'h1):(1'h0)] ~^ reg876));
              reg910 = {reg885[(5'h17):(4'hc)],
                  ((^$signed($signed(reg883))) ?
                      $unsigned(reg885[(1'h1):(1'h1)]) : $signed(forvar868[(5'h13):(5'h12)])),
                  reg849[(2'h3):(2'h2)]};
              reg911 <= (forvar884[(1'h1):(1'h0)] ?
                  $signed(reg864[(3'h5):(3'h4)]) : (&$signed(((^~reg51) ?
                      forvar848[(2'h2):(1'h0)] : reg894))));
              reg912 <= reg900;
              reg913 <= $unsigned((7'h4f));
              reg914 <= {(forvar884[(3'h6):(3'h6)] >>> ({reg869, reg21} ?
                      (((8'h9c) ~^ reg869) << reg11) : reg860)),
                  $signed({(wire70[(4'hd):(1'h1)] >= $unsigned(reg868)),
                      $unsigned($signed(reg872)),
                      {$signed(reg864), reg898}}),
                  $signed($signed(reg863[(4'h9):(1'h1)]))};
              reg915 <= $signed($unsigned($signed(reg879)));
            end
          for (forvar916 = (1'h0); (forvar916 < (1'h0)); forvar916 = (forvar916 + (1'h1)))
            begin
              reg917 = (7'h4a);
              reg918 = $signed(((^~$unsigned((wire9 ?
                  reg909 : reg883))) ^~ ($unsigned($unsigned(reg873)) ?
                  (~|(reg875 > (7'h56))) : $unsigned(reg903[(5'h13):(4'h8)]))));
              reg919 <= $signed({($unsigned($unsigned(reg915)) ?
                      ({reg62} ? $unsigned(reg895) : (&reg915)) : reg39)});
              reg920 = ((^~reg41) >= (($unsigned($signed(reg882)) ?
                      $unsigned(reg905[(4'h8):(3'h4)]) : reg877) ?
                  reg896 : ($unsigned(reg851) + reg855)));
              reg921 = $unsigned($unsigned((+reg20)));
            end
          reg922 = (forvar870 || (~^reg864[(3'h5):(1'h1)]));
        end
    end
  module923 #() modinst3070 (.y(wire3069), .wire925(wire7), .wire924(reg919), .clk(clk), .wire928(reg21), .wire926(reg880), .wire927(reg879));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module923
#(parameter param3066 = (((^~(((7'h4b) - (8'ha6)) ? (-(8'ha6)) : (8'hbe))) ? (((+(8'hae)) ? (|(8'h9c)) : (~(8'ha0))) >>> (((7'h4f) != (8'hb8)) ? {(7'h44), (8'hba)} : ((7'h4a) ? (7'h57) : (7'h49)))) : ({(^(8'hab))} ? (^(~&(7'h4e))) : {{(8'hba)}})) >> (({((7'h43) >= (8'ha4)), (~(8'hbf)), ((8'hb0) > (8'hab))} >>> ((^~(8'h9c)) & ((8'hbb) ? (7'h40) : (8'ha7)))) ^~ ((((7'h4b) >= (8'hbb)) >> {(8'ha1)}) ? ({(8'haa), (8'hb7)} ~^ (~&(7'h44))) : ({(8'hb1)} ? (~&(8'hb4)) : (+(7'h4e)))))), 
parameter param3067 = ({(&{(param3066 != (8'ha5)), param3066}), (|(^(&param3066))), (^~(param3066 ? ((8'hb3) ^ param3066) : (^param3066)))} >= (^((!((7'h57) ^ param3066)) ? (^((8'hb0) <= param3066)) : param3066))), 
parameter param3068 = (^~(param3066 ? param3067 : {((param3066 && param3067) ? ((8'hb3) + param3066) : ((7'h4d) == param3067))})))
(y, clk, wire924, wire925, wire926, wire927, wire928);
  output wire [(32'h3166):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire924;
  input wire [(4'h8):(1'h0)] wire925;
  input wire signed [(4'h8):(1'h0)] wire926;
  input wire [(5'h19):(1'h0)] wire927;
  input wire [(5'h19):(1'h0)] wire928;
  wire [(5'h19):(1'h0)] wire2804;
  wire [(2'h2):(1'h0)] wire2339;
  wire [(3'h5):(1'h0)] wire2338;
  wire signed [(5'h1a):(1'h0)] wire2337;
  wire signed [(4'h8):(1'h0)] wire2260;
  wire signed [(4'hb):(1'h0)] wire2195;
  wire [(5'h1b):(1'h0)] wire1772;
  wire signed [(5'h17):(1'h0)] wire1013;
  wire signed [(5'h18):(1'h0)] wire1327;
  wire [(5'h1f):(1'h0)] wire1770;
  wire [(5'h1d):(1'h0)] wire3064;
  reg signed [(4'ha):(1'h0)] reg3062 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3059 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3058 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3055 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3054 = (1'h0);
  reg [(5'h15):(1'h0)] reg3051 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3049 = (1'h0);
  reg [(4'ha):(1'h0)] reg3048 = (1'h0);
  reg [(5'h12):(1'h0)] reg3045 = (1'h0);
  reg [(2'h3):(1'h0)] reg3044 = (1'h0);
  reg [(2'h2):(1'h0)] reg3043 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3042 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3040 = (1'h0);
  reg [(4'h8):(1'h0)] reg3036 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3035 = (1'h0);
  reg [(3'h5):(1'h0)] reg3034 = (1'h0);
  reg [(4'hf):(1'h0)] reg3033 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3032 = (1'h0);
  reg [(4'ha):(1'h0)] reg3030 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3027 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3026 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3024 = (1'h0);
  reg [(4'hb):(1'h0)] reg3020 = (1'h0);
  reg [(5'h14):(1'h0)] reg3017 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3016 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3014 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3011 = (1'h0);
  reg [(5'h16):(1'h0)] reg3010 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3008 = (1'h0);
  reg [(5'h13):(1'h0)] reg3004 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3002 = (1'h0);
  reg [(5'h14):(1'h0)] reg2996 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2995 = (1'h0);
  reg [(5'h17):(1'h0)] reg2992 = (1'h0);
  reg [(3'h5):(1'h0)] reg2991 = (1'h0);
  reg [(5'h17):(1'h0)] reg2990 = (1'h0);
  reg [(5'h12):(1'h0)] reg2987 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2984 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2983 = (1'h0);
  reg [(4'ha):(1'h0)] reg2982 = (1'h0);
  reg [(4'hb):(1'h0)] reg2979 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2977 = (1'h0);
  reg [(4'hf):(1'h0)] reg2974 = (1'h0);
  reg [(4'hd):(1'h0)] reg2973 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2972 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2971 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2968 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2966 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2964 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2962 = (1'h0);
  reg [(5'h13):(1'h0)] reg2961 = (1'h0);
  reg [(4'hf):(1'h0)] reg2960 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2958 = (1'h0);
  reg [(3'h5):(1'h0)] reg2955 = (1'h0);
  reg [(5'h15):(1'h0)] reg2954 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2953 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2951 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2947 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2946 = (1'h0);
  reg [(5'h10):(1'h0)] reg2942 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2936 = (1'h0);
  reg [(5'h11):(1'h0)] reg2935 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2932 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2928 = (1'h0);
  reg [(4'ha):(1'h0)] reg2926 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2924 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2919 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2918 = (1'h0);
  reg [(5'h12):(1'h0)] reg2916 = (1'h0);
  reg [(4'hd):(1'h0)] reg2915 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2913 = (1'h0);
  reg [(5'h13):(1'h0)] reg2911 = (1'h0);
  reg [(4'hf):(1'h0)] reg2909 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2907 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2905 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2902 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2899 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2897 = (1'h0);
  reg [(4'ha):(1'h0)] reg2895 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2894 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2893 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2891 = (1'h0);
  reg [(4'hb):(1'h0)] reg2888 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2887 = (1'h0);
  reg [(2'h3):(1'h0)] reg2881 = (1'h0);
  reg [(5'h10):(1'h0)] reg2879 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2878 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2877 = (1'h0);
  reg [(4'h9):(1'h0)] reg2874 = (1'h0);
  reg [(5'h12):(1'h0)] reg2873 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2872 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2870 = (1'h0);
  reg [(4'hf):(1'h0)] reg2867 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2866 = (1'h0);
  reg [(4'he):(1'h0)] reg2865 = (1'h0);
  reg [(2'h2):(1'h0)] reg2864 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2863 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2862 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2861 = (1'h0);
  reg [(4'hb):(1'h0)] reg2854 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2853 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2851 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2848 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2846 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2845 = (1'h0);
  reg [(5'h11):(1'h0)] reg2842 = (1'h0);
  reg [(4'h8):(1'h0)] reg2835 = (1'h0);
  reg [(4'he):(1'h0)] reg2829 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2828 = (1'h0);
  reg [(4'ha):(1'h0)] reg2826 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2823 = (1'h0);
  reg [(4'hb):(1'h0)] reg2822 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2816 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2814 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2812 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2811 = (1'h0);
  reg [(5'h19):(1'h0)] reg2810 = (1'h0);
  reg [(5'h16):(1'h0)] reg2809 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2806 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2461 = (1'h0);
  reg [(5'h19):(1'h0)] reg2460 = (1'h0);
  reg [(5'h13):(1'h0)] reg2457 = (1'h0);
  reg [(3'h4):(1'h0)] reg2456 = (1'h0);
  reg [(4'ha):(1'h0)] reg2455 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2453 = (1'h0);
  reg [(4'h8):(1'h0)] reg2452 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2451 = (1'h0);
  reg [(3'h7):(1'h0)] reg2449 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2448 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2447 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2440 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2439 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2438 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2436 = (1'h0);
  reg [(4'he):(1'h0)] reg2435 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2433 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2432 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2430 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2429 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2428 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2427 = (1'h0);
  reg [(3'h5):(1'h0)] reg2425 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2423 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2421 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2419 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2418 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2415 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2413 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2411 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2405 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2404 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2401 = (1'h0);
  reg [(5'h11):(1'h0)] reg2398 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2397 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2396 = (1'h0);
  reg [(5'h19):(1'h0)] reg2394 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2391 = (1'h0);
  reg [(4'hc):(1'h0)] reg2390 = (1'h0);
  reg [(3'h6):(1'h0)] reg2389 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2388 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2387 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2385 = (1'h0);
  reg [(5'h19):(1'h0)] reg2383 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2382 = (1'h0);
  reg [(3'h7):(1'h0)] reg2381 = (1'h0);
  reg [(2'h3):(1'h0)] reg2380 = (1'h0);
  reg [(5'h16):(1'h0)] reg2378 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2368 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2367 = (1'h0);
  reg [(3'h6):(1'h0)] reg2363 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2362 = (1'h0);
  reg [(5'h16):(1'h0)] reg2360 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2359 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2358 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2357 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2356 = (1'h0);
  reg [(3'h4):(1'h0)] reg2341 = (1'h0);
  reg [(5'h12):(1'h0)] reg2353 = (1'h0);
  reg [(5'h11):(1'h0)] reg2351 = (1'h0);
  reg [(4'h8):(1'h0)] reg2349 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2347 = (1'h0);
  reg [(4'hb):(1'h0)] reg2345 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2344 = (1'h0);
  reg [(3'h4):(1'h0)] reg2342 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2340 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2336 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2331 = (1'h0);
  reg [(3'h5):(1'h0)] reg2329 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2328 = (1'h0);
  reg [(5'h11):(1'h0)] reg2327 = (1'h0);
  reg [(3'h4):(1'h0)] reg2323 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2321 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2320 = (1'h0);
  reg [(3'h6):(1'h0)] reg2319 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2316 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2315 = (1'h0);
  reg [(5'h12):(1'h0)] reg2313 = (1'h0);
  reg [(5'h14):(1'h0)] reg2312 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2309 = (1'h0);
  reg [(2'h2):(1'h0)] reg2307 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2306 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2265 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2304 = (1'h0);
  reg [(4'hf):(1'h0)] reg2302 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2301 = (1'h0);
  reg [(5'h13):(1'h0)] reg2298 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2297 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2296 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2293 = (1'h0);
  reg [(4'hb):(1'h0)] reg2292 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2291 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2290 = (1'h0);
  reg [(5'h10):(1'h0)] reg2287 = (1'h0);
  reg [(5'h14):(1'h0)] reg2286 = (1'h0);
  reg [(5'h19):(1'h0)] reg2285 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2283 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2282 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2281 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2279 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2276 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2274 = (1'h0);
  reg [(5'h10):(1'h0)] reg2273 = (1'h0);
  reg [(5'h11):(1'h0)] reg2271 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2270 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2269 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2268 = (1'h0);
  reg [(5'h12):(1'h0)] reg2267 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2266 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2264 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2263 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2255 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2248 = (1'h0);
  reg [(4'h8):(1'h0)] reg2247 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2246 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2242 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2235 = (1'h0);
  reg [(4'hc):(1'h0)] reg2234 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2232 = (1'h0);
  reg [(5'h12):(1'h0)] reg2230 = (1'h0);
  reg [(5'h15):(1'h0)] reg2228 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2225 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2224 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2223 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2222 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2221 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2217 = (1'h0);
  reg [(5'h18):(1'h0)] reg2216 = (1'h0);
  reg [(4'hb):(1'h0)] reg2215 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2213 = (1'h0);
  reg [(5'h16):(1'h0)] reg2209 = (1'h0);
  reg [(2'h3):(1'h0)] reg2203 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2202 = (1'h0);
  reg [(5'h19):(1'h0)] reg2199 = (1'h0);
  reg [(4'hc):(1'h0)] reg1057 = (1'h0);
  reg [(4'hc):(1'h0)] reg1054 = (1'h0);
  reg [(5'h18):(1'h0)] reg1052 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1050 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1047 = (1'h0);
  reg [(5'h13):(1'h0)] reg1046 = (1'h0);
  reg [(5'h15):(1'h0)] reg1044 = (1'h0);
  reg [(3'h4):(1'h0)] reg1043 = (1'h0);
  reg [(5'h17):(1'h0)] reg1036 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1025 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1023 = (1'h0);
  reg [(5'h13):(1'h0)] reg1020 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1002 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1010 = (1'h0);
  reg [(5'h12):(1'h0)] reg1009 = (1'h0);
  reg [(5'h17):(1'h0)] reg1005 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1001 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg997 = (1'h0);
  reg [(5'h11):(1'h0)] reg996 = (1'h0);
  reg [(3'h5):(1'h0)] reg995 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg994 = (1'h0);
  reg [(2'h2):(1'h0)] reg991 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg990 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg989 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg988 = (1'h0);
  reg [(4'hb):(1'h0)] reg986 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg985 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg982 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg981 = (1'h0);
  reg [(3'h5):(1'h0)] reg979 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg978 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg961 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg976 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg972 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg970 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg966 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg964 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg963 = (1'h0);
  reg [(5'h1b):(1'h0)] reg962 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg959 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg957 = (1'h0);
  reg [(5'h16):(1'h0)] reg956 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg955 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg952 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg945 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg944 = (1'h0);
  reg [(5'h1d):(1'h0)] reg943 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg941 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg940 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg936 = (1'h0);
  reg [(2'h3):(1'h0)] reg933 = (1'h0);
  reg signed [(4'he):(1'h0)] reg932 = (1'h0);
  reg [(5'h1d):(1'h0)] reg931 = (1'h0);
  reg [(4'he):(1'h0)] reg1333 = (1'h0);
  reg [(5'h11):(1'h0)] reg1335 = (1'h0);
  reg [(4'hc):(1'h0)] reg1338 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1339 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1343 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1344 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1345 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1346 = (1'h0);
  reg [(5'h11):(1'h0)] reg1347 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1349 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1351 = (1'h0);
  reg [(4'hd):(1'h0)] reg1352 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1353 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1355 = (1'h0);
  reg [(5'h14):(1'h0)] reg1357 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1359 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1362 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1365 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1369 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1370 = (1'h0);
  reg [(4'hd):(1'h0)] reg1371 = (1'h0);
  reg [(5'h17):(1'h0)] reg1372 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1373 = (1'h0);
  reg [(5'h14):(1'h0)] reg1374 = (1'h0);
  reg [(4'hf):(1'h0)] reg1375 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3063 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3061 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3060 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3057 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3056 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3053 = (1'h0);
  reg [(5'h11):(1'h0)] reg3052 = (1'h0);
  reg [(5'h12):(1'h0)] forvar3050 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3047 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3044 = (1'h0);
  reg [(5'h11):(1'h0)] reg3046 = (1'h0);
  reg [(3'h4):(1'h0)] reg3041 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3039 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar3038 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3037 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3031 = (1'h0);
  reg [(5'h14):(1'h0)] reg3029 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3028 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3025 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar3023 = (1'h0);
  reg [(3'h7):(1'h0)] reg3022 = (1'h0);
  reg [(4'hf):(1'h0)] reg3021 = (1'h0);
  reg [(4'ha):(1'h0)] reg3019 = (1'h0);
  reg [(4'he):(1'h0)] reg3018 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar3015 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3013 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3012 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3009 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3006 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3005 = (1'h0);
  reg [(5'h15):(1'h0)] reg3007 = (1'h0);
  reg [(3'h4):(1'h0)] reg3006 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3005 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3003 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3001 = (1'h0);
  reg [(5'h12):(1'h0)] reg3000 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2999 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2998 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2997 = (1'h0);
  reg [(5'h16):(1'h0)] reg2994 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2993 = (1'h0);
  reg [(5'h19):(1'h0)] reg2989 = (1'h0);
  reg [(5'h13):(1'h0)] reg2988 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2986 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2985 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2981 = (1'h0);
  reg [(4'hd):(1'h0)] reg2980 = (1'h0);
  reg [(4'hd):(1'h0)] reg2978 = (1'h0);
  reg [(4'ha):(1'h0)] reg2976 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2975 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2970 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2969 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2967 = (1'h0);
  reg [(5'h16):(1'h0)] reg2965 = (1'h0);
  reg [(2'h2):(1'h0)] reg2963 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2959 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2957 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar2956 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2952 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2950 = (1'h0);
  reg [(4'h8):(1'h0)] reg2949 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2948 = (1'h0);
  reg [(4'ha):(1'h0)] reg2945 = (1'h0);
  reg [(3'h5):(1'h0)] reg2944 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2943 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2941 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2940 = (1'h0);
  reg [(3'h5):(1'h0)] reg2939 = (1'h0);
  reg [(5'h11):(1'h0)] reg2938 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2937 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2934 = (1'h0);
  reg [(5'h15):(1'h0)] reg2933 = (1'h0);
  reg [(5'h18):(1'h0)] reg2931 = (1'h0);
  reg [(2'h3):(1'h0)] reg2930 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2929 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2927 = (1'h0);
  reg [(5'h18):(1'h0)] reg2925 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2923 = (1'h0);
  reg [(4'hc):(1'h0)] reg2922 = (1'h0);
  reg [(3'h5):(1'h0)] reg2921 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2920 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2917 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2914 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar2912 = (1'h0);
  reg [(5'h17):(1'h0)] reg2910 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2908 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2906 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2904 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2903 = (1'h0);
  reg [(4'ha):(1'h0)] reg2901 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2900 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2898 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2894 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2886 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2885 = (1'h0);
  reg [(3'h4):(1'h0)] reg2896 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2892 = (1'h0);
  reg [(3'h5):(1'h0)] reg2890 = (1'h0);
  reg [(5'h10):(1'h0)] reg2889 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar2886 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2885 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2884 = (1'h0);
  reg [(3'h7):(1'h0)] reg2883 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2882 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2880 = (1'h0);
  reg [(5'h14):(1'h0)] reg2876 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2875 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2871 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2860 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2869 = (1'h0);
  reg [(5'h13):(1'h0)] reg2868 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2860 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2859 = (1'h0);
  reg [(5'h17):(1'h0)] reg2858 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2857 = (1'h0);
  reg [(5'h14):(1'h0)] reg2856 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2855 = (1'h0);
  reg [(4'hd):(1'h0)] reg2852 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2850 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2849 = (1'h0);
  reg [(5'h16):(1'h0)] reg2847 = (1'h0);
  reg [(5'h18):(1'h0)] reg2844 = (1'h0);
  reg [(5'h15):(1'h0)] reg2843 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2841 = (1'h0);
  reg [(4'hc):(1'h0)] reg2840 = (1'h0);
  reg [(4'hc):(1'h0)] reg2839 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2838 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2837 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2836 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2834 = (1'h0);
  reg [(5'h10):(1'h0)] reg2833 = (1'h0);
  reg [(4'he):(1'h0)] reg2832 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2831 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2830 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2827 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2825 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2824 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2821 = (1'h0);
  reg [(5'h12):(1'h0)] reg2820 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2819 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2818 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2817 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar2815 = (1'h0);
  reg [(5'h15):(1'h0)] reg2813 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2808 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2807 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2466 = (1'h0);
  reg [(3'h4):(1'h0)] reg2465 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2464 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2463 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2462 = (1'h0);
  reg [(4'hc):(1'h0)] reg2459 = (1'h0);
  reg [(3'h6):(1'h0)] reg2458 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2454 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2450 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2446 = (1'h0);
  reg [(5'h11):(1'h0)] reg2445 = (1'h0);
  reg [(5'h15):(1'h0)] reg2444 = (1'h0);
  reg [(4'hf):(1'h0)] reg2443 = (1'h0);
  reg [(2'h3):(1'h0)] reg2442 = (1'h0);
  reg [(5'h14):(1'h0)] reg2441 = (1'h0);
  reg [(4'hf):(1'h0)] reg2437 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2434 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2431 = (1'h0);
  reg [(5'h17):(1'h0)] reg2426 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2424 = (1'h0);
  reg [(5'h17):(1'h0)] reg2422 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2420 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2417 = (1'h0);
  reg [(4'hf):(1'h0)] reg2416 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2408 = (1'h0);
  reg [(5'h18):(1'h0)] reg2402 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2400 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2399 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2414 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2412 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2410 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2409 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2408 = (1'h0);
  reg [(5'h12):(1'h0)] reg2407 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2406 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2403 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2402 = (1'h0);
  reg [(3'h4):(1'h0)] reg2400 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2399 = (1'h0);
  reg [(4'h8):(1'h0)] reg2395 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2393 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2392 = (1'h0);
  reg [(4'h8):(1'h0)] reg2386 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2384 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2379 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2377 = (1'h0);
  reg [(4'hc):(1'h0)] reg2376 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2375 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2374 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2373 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2372 = (1'h0);
  reg [(5'h10):(1'h0)] reg2371 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2370 = (1'h0);
  reg [(3'h5):(1'h0)] reg2369 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2366 = (1'h0);
  reg [(4'hc):(1'h0)] reg2365 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2364 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2361 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2355 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2354 = (1'h0);
  reg [(3'h6):(1'h0)] reg2352 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2350 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2348 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2346 = (1'h0);
  reg [(5'h12):(1'h0)] reg2343 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar2341 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2335 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2334 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2333 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2332 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2330 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2326 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2325 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2324 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2322 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2318 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2317 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2314 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2311 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2310 = (1'h0);
  reg [(4'hb):(1'h0)] reg2308 = (1'h0);
  reg [(4'ha):(1'h0)] reg2305 = (1'h0);
  reg [(3'h5):(1'h0)] reg2299 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2275 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2266 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2303 = (1'h0);
  reg [(4'he):(1'h0)] reg2300 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2299 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2295 = (1'h0);
  reg [(5'h17):(1'h0)] reg2294 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2289 = (1'h0);
  reg [(4'h9):(1'h0)] reg2288 = (1'h0);
  reg [(4'hb):(1'h0)] reg2284 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2280 = (1'h0);
  reg [(5'h11):(1'h0)] reg2278 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2277 = (1'h0);
  reg [(4'h9):(1'h0)] reg2275 = (1'h0);
  reg [(2'h3):(1'h0)] reg2272 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2265 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2262 = (1'h0);
  reg [(2'h3):(1'h0)] reg2261 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2259 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2258 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2257 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2256 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2236 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2254 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2253 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2252 = (1'h0);
  reg [(4'ha):(1'h0)] reg2251 = (1'h0);
  reg [(5'h18):(1'h0)] reg2250 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2249 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2245 = (1'h0);
  reg [(3'h4):(1'h0)] reg2244 = (1'h0);
  reg [(5'h14):(1'h0)] reg2243 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2241 = (1'h0);
  reg [(4'hc):(1'h0)] reg2240 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2239 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2238 = (1'h0);
  reg [(5'h16):(1'h0)] reg2237 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2236 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2233 = (1'h0);
  reg [(5'h14):(1'h0)] reg2231 = (1'h0);
  reg [(2'h2):(1'h0)] reg2229 = (1'h0);
  reg [(2'h3):(1'h0)] reg2227 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2226 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar2214 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2212 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar2220 = (1'h0);
  reg [(2'h3):(1'h0)] reg2219 = (1'h0);
  reg [(2'h2):(1'h0)] reg2218 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2214 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar2212 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2211 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2210 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2208 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2207 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2206 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2205 = (1'h0);
  reg [(3'h6):(1'h0)] reg2204 = (1'h0);
  reg [(5'h17):(1'h0)] reg2201 = (1'h0);
  reg [(5'h18):(1'h0)] reg2200 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2198 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2197 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1368 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1367 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1366 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1364 = (1'h0);
  reg [(4'hb):(1'h0)] reg1363 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1361 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1360 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1358 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1356 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1354 = (1'h0);
  reg [(2'h2):(1'h0)] reg1331 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1330 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1350 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1348 = (1'h0);
  reg [(5'h10):(1'h0)] reg1342 = (1'h0);
  reg [(5'h12):(1'h0)] reg1341 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1340 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1337 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1336 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1334 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1332 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1331 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1330 = (1'h0);
  reg [(4'hd):(1'h0)] reg1329 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1058 = (1'h0);
  reg [(2'h3):(1'h0)] reg1056 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1055 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1053 = (1'h0);
  reg [(5'h14):(1'h0)] reg1051 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1049 = (1'h0);
  reg [(4'hb):(1'h0)] reg1048 = (1'h0);
  reg [(4'hb):(1'h0)] reg1045 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1042 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1041 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1040 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1039 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1038 = (1'h0);
  reg [(4'hd):(1'h0)] reg1037 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1035 = (1'h0);
  reg [(5'h17):(1'h0)] reg1034 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1033 = (1'h0);
  reg [(3'h4):(1'h0)] reg1032 = (1'h0);
  reg [(4'h9):(1'h0)] reg1031 = (1'h0);
  reg [(5'h15):(1'h0)] reg1030 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1029 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1028 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1027 = (1'h0);
  reg [(4'hd):(1'h0)] reg1026 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1024 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1022 = (1'h0);
  reg [(2'h3):(1'h0)] reg1021 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1019 = (1'h0);
  reg [(4'h8):(1'h0)] reg1018 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1017 = (1'h0);
  reg [(2'h3):(1'h0)] reg1016 = (1'h0);
  reg [(5'h17):(1'h0)] reg1015 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1014 = (1'h0);
  reg [(5'h15):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1011 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1003 = (1'h0);
  reg [(2'h3):(1'h0)] forvar999 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1008 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1007 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1006 = (1'h0);
  reg [(4'h9):(1'h0)] reg1004 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1003 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1002 = (1'h0);
  reg [(5'h12):(1'h0)] reg1000 = (1'h0);
  reg [(5'h15):(1'h0)] reg999 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg998 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg993 = (1'h0);
  reg [(5'h19):(1'h0)] reg992 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg987 = (1'h0);
  reg [(5'h19):(1'h0)] reg984 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg983 = (1'h0);
  reg [(2'h2):(1'h0)] forvar980 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar977 = (1'h0);
  reg [(4'ha):(1'h0)] reg975 = (1'h0);
  reg [(4'hd):(1'h0)] reg974 = (1'h0);
  reg [(5'h1c):(1'h0)] reg973 = (1'h0);
  reg [(5'h18):(1'h0)] reg971 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg969 = (1'h0);
  reg [(5'h18):(1'h0)] reg968 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg967 = (1'h0);
  reg [(4'hb):(1'h0)] reg965 = (1'h0);
  reg [(3'h7):(1'h0)] forvar961 = (1'h0);
  reg [(3'h7):(1'h0)] reg960 = (1'h0);
  reg [(4'hf):(1'h0)] reg958 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg954 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg953 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg951 = (1'h0);
  reg [(5'h17):(1'h0)] reg950 = (1'h0);
  reg [(4'hd):(1'h0)] reg949 = (1'h0);
  reg [(4'hd):(1'h0)] reg948 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg947 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar946 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar942 = (1'h0);
  reg [(5'h10):(1'h0)] forvar929 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg939 = (1'h0);
  reg [(5'h18):(1'h0)] reg938 = (1'h0);
  reg [(3'h6):(1'h0)] reg937 = (1'h0);
  reg [(5'h18):(1'h0)] forvar936 = (1'h0);
  reg [(4'he):(1'h0)] reg935 = (1'h0);
  reg [(5'h17):(1'h0)] reg934 = (1'h0);
  reg [(5'h16):(1'h0)] reg930 = (1'h0);
  reg [(4'ha):(1'h0)] reg929 = (1'h0);
  assign y = {wire2804,
                 wire2339,
                 wire2338,
                 wire2337,
                 wire2260,
                 wire2195,
                 wire1772,
                 wire1013,
                 wire1327,
                 wire1770,
                 wire3064,
                 reg3062,
                 reg3059,
                 reg3058,
                 reg3055,
                 reg3054,
                 reg3051,
                 reg3049,
                 reg3048,
                 reg3045,
                 reg3044,
                 reg3043,
                 reg3042,
                 reg3040,
                 reg3036,
                 reg3035,
                 reg3034,
                 reg3033,
                 reg3032,
                 reg3030,
                 reg3027,
                 reg3026,
                 reg3024,
                 reg3020,
                 reg3017,
                 reg3016,
                 reg3014,
                 reg3011,
                 reg3010,
                 reg3008,
                 reg3004,
                 reg3002,
                 reg2996,
                 reg2995,
                 reg2992,
                 reg2991,
                 reg2990,
                 reg2987,
                 reg2984,
                 reg2983,
                 reg2982,
                 reg2979,
                 reg2977,
                 reg2974,
                 reg2973,
                 reg2972,
                 reg2971,
                 reg2968,
                 reg2966,
                 reg2964,
                 reg2962,
                 reg2961,
                 reg2960,
                 reg2958,
                 reg2955,
                 reg2954,
                 reg2953,
                 reg2951,
                 reg2947,
                 reg2946,
                 reg2942,
                 reg2936,
                 reg2935,
                 reg2932,
                 reg2928,
                 reg2926,
                 reg2924,
                 reg2919,
                 reg2918,
                 reg2916,
                 reg2915,
                 reg2913,
                 reg2911,
                 reg2909,
                 reg2907,
                 reg2905,
                 reg2902,
                 reg2899,
                 reg2897,
                 reg2895,
                 reg2894,
                 reg2893,
                 reg2891,
                 reg2888,
                 reg2887,
                 reg2881,
                 reg2879,
                 reg2878,
                 reg2877,
                 reg2874,
                 reg2873,
                 reg2872,
                 reg2870,
                 reg2867,
                 reg2866,
                 reg2865,
                 reg2864,
                 reg2863,
                 reg2862,
                 reg2861,
                 reg2854,
                 reg2853,
                 reg2851,
                 reg2848,
                 reg2846,
                 reg2845,
                 reg2842,
                 reg2835,
                 reg2829,
                 reg2828,
                 reg2826,
                 reg2823,
                 reg2822,
                 reg2816,
                 reg2814,
                 reg2812,
                 reg2811,
                 reg2810,
                 reg2809,
                 reg2806,
                 reg2461,
                 reg2460,
                 reg2457,
                 reg2456,
                 reg2455,
                 reg2453,
                 reg2452,
                 reg2451,
                 reg2449,
                 reg2448,
                 reg2447,
                 reg2440,
                 reg2439,
                 reg2438,
                 reg2436,
                 reg2435,
                 reg2433,
                 reg2432,
                 reg2430,
                 reg2429,
                 reg2428,
                 reg2427,
                 reg2425,
                 reg2423,
                 reg2421,
                 reg2419,
                 reg2418,
                 reg2415,
                 reg2413,
                 reg2411,
                 reg2405,
                 reg2404,
                 reg2401,
                 reg2398,
                 reg2397,
                 reg2396,
                 reg2394,
                 reg2391,
                 reg2390,
                 reg2389,
                 reg2388,
                 reg2387,
                 reg2385,
                 reg2383,
                 reg2382,
                 reg2381,
                 reg2380,
                 reg2378,
                 reg2368,
                 reg2367,
                 reg2363,
                 reg2362,
                 reg2360,
                 reg2359,
                 reg2358,
                 reg2357,
                 reg2356,
                 reg2341,
                 reg2353,
                 reg2351,
                 reg2349,
                 reg2347,
                 reg2345,
                 reg2344,
                 reg2342,
                 reg2340,
                 reg2336,
                 reg2331,
                 reg2329,
                 reg2328,
                 reg2327,
                 reg2323,
                 reg2321,
                 reg2320,
                 reg2319,
                 reg2316,
                 reg2315,
                 reg2313,
                 reg2312,
                 reg2309,
                 reg2307,
                 reg2306,
                 reg2265,
                 reg2304,
                 reg2302,
                 reg2301,
                 reg2298,
                 reg2297,
                 reg2296,
                 reg2293,
                 reg2292,
                 reg2291,
                 reg2290,
                 reg2287,
                 reg2286,
                 reg2285,
                 reg2283,
                 reg2282,
                 reg2281,
                 reg2279,
                 reg2276,
                 reg2274,
                 reg2273,
                 reg2271,
                 reg2270,
                 reg2269,
                 reg2268,
                 reg2267,
                 reg2266,
                 reg2264,
                 reg2263,
                 reg2255,
                 reg2248,
                 reg2247,
                 reg2246,
                 reg2242,
                 reg2235,
                 reg2234,
                 reg2232,
                 reg2230,
                 reg2228,
                 reg2225,
                 reg2224,
                 reg2223,
                 reg2222,
                 reg2221,
                 reg2217,
                 reg2216,
                 reg2215,
                 reg2213,
                 reg2209,
                 reg2203,
                 reg2202,
                 reg2199,
                 reg1057,
                 reg1054,
                 reg1052,
                 reg1050,
                 reg1047,
                 reg1046,
                 reg1044,
                 reg1043,
                 reg1036,
                 reg1025,
                 reg1023,
                 reg1020,
                 reg1002,
                 reg1010,
                 reg1009,
                 reg1005,
                 reg1001,
                 reg997,
                 reg996,
                 reg995,
                 reg994,
                 reg991,
                 reg990,
                 reg989,
                 reg988,
                 reg986,
                 reg985,
                 reg982,
                 reg981,
                 reg979,
                 reg978,
                 reg961,
                 reg976,
                 reg972,
                 reg970,
                 reg966,
                 reg964,
                 reg963,
                 reg962,
                 reg959,
                 reg957,
                 reg956,
                 reg955,
                 reg952,
                 reg945,
                 reg944,
                 reg943,
                 reg941,
                 reg940,
                 reg936,
                 reg933,
                 reg932,
                 reg931,
                 reg1333,
                 reg1335,
                 reg1338,
                 reg1339,
                 reg1343,
                 reg1344,
                 reg1345,
                 reg1346,
                 reg1347,
                 reg1349,
                 reg1351,
                 reg1352,
                 reg1353,
                 reg1355,
                 reg1357,
                 reg1359,
                 reg1362,
                 reg1365,
                 reg1369,
                 reg1370,
                 reg1371,
                 reg1372,
                 reg1373,
                 reg1374,
                 reg1375,
                 reg3063,
                 reg3061,
                 reg3060,
                 forvar3057,
                 reg3056,
                 reg3053,
                 reg3052,
                 forvar3050,
                 reg3047,
                 forvar3044,
                 reg3046,
                 reg3041,
                 reg3039,
                 forvar3038,
                 reg3037,
                 forvar3031,
                 reg3029,
                 reg3028,
                 reg3025,
                 forvar3023,
                 reg3022,
                 reg3021,
                 reg3019,
                 reg3018,
                 forvar3015,
                 reg3013,
                 reg3012,
                 reg3009,
                 forvar3006,
                 reg3005,
                 reg3007,
                 reg3006,
                 forvar3005,
                 reg3003,
                 reg3001,
                 reg3000,
                 forvar2999,
                 reg2998,
                 forvar2997,
                 reg2994,
                 forvar2993,
                 reg2989,
                 reg2988,
                 reg2986,
                 reg2985,
                 forvar2981,
                 reg2980,
                 reg2978,
                 reg2976,
                 reg2975,
                 reg2970,
                 reg2969,
                 forvar2967,
                 reg2965,
                 reg2963,
                 reg2959,
                 reg2957,
                 forvar2956,
                 reg2952,
                 reg2950,
                 reg2949,
                 forvar2948,
                 reg2945,
                 reg2944,
                 reg2943,
                 reg2941,
                 reg2940,
                 reg2939,
                 reg2938,
                 reg2937,
                 reg2934,
                 reg2933,
                 reg2931,
                 reg2930,
                 forvar2929,
                 reg2927,
                 reg2925,
                 reg2923,
                 reg2922,
                 reg2921,
                 reg2920,
                 reg2917,
                 reg2914,
                 forvar2912,
                 reg2910,
                 reg2908,
                 reg2906,
                 reg2904,
                 reg2903,
                 reg2901,
                 reg2900,
                 reg2898,
                 forvar2894,
                 reg2886,
                 forvar2885,
                 reg2896,
                 reg2892,
                 reg2890,
                 reg2889,
                 forvar2886,
                 reg2885,
                 reg2884,
                 reg2883,
                 forvar2882,
                 reg2880,
                 reg2876,
                 reg2875,
                 reg2871,
                 forvar2860,
                 reg2869,
                 reg2868,
                 reg2860,
                 reg2859,
                 reg2858,
                 reg2857,
                 reg2856,
                 reg2855,
                 reg2852,
                 forvar2850,
                 reg2849,
                 reg2847,
                 reg2844,
                 reg2843,
                 reg2841,
                 reg2840,
                 reg2839,
                 reg2838,
                 reg2837,
                 reg2836,
                 reg2834,
                 reg2833,
                 reg2832,
                 reg2831,
                 reg2830,
                 forvar2827,
                 reg2825,
                 reg2824,
                 reg2821,
                 reg2820,
                 forvar2819,
                 reg2818,
                 reg2817,
                 forvar2815,
                 reg2813,
                 forvar2808,
                 forvar2807,
                 reg2466,
                 reg2465,
                 reg2464,
                 reg2463,
                 reg2462,
                 reg2459,
                 reg2458,
                 reg2454,
                 reg2450,
                 reg2446,
                 reg2445,
                 reg2444,
                 reg2443,
                 reg2442,
                 reg2441,
                 reg2437,
                 reg2434,
                 reg2431,
                 reg2426,
                 reg2424,
                 reg2422,
                 forvar2420,
                 reg2417,
                 reg2416,
                 reg2408,
                 reg2402,
                 forvar2400,
                 reg2399,
                 reg2414,
                 reg2412,
                 reg2410,
                 reg2409,
                 forvar2408,
                 reg2407,
                 reg2406,
                 reg2403,
                 forvar2402,
                 reg2400,
                 forvar2399,
                 reg2395,
                 reg2393,
                 forvar2392,
                 reg2386,
                 reg2384,
                 reg2379,
                 forvar2377,
                 reg2376,
                 reg2375,
                 reg2374,
                 forvar2373,
                 reg2372,
                 reg2371,
                 reg2370,
                 reg2369,
                 forvar2366,
                 reg2365,
                 forvar2364,
                 reg2361,
                 reg2355,
                 reg2354,
                 reg2352,
                 reg2350,
                 reg2348,
                 reg2346,
                 reg2343,
                 forvar2341,
                 reg2335,
                 reg2334,
                 reg2333,
                 reg2332,
                 reg2330,
                 reg2326,
                 reg2325,
                 reg2324,
                 reg2322,
                 reg2318,
                 reg2317,
                 reg2314,
                 reg2311,
                 reg2310,
                 reg2308,
                 reg2305,
                 reg2299,
                 forvar2275,
                 forvar2266,
                 reg2303,
                 reg2300,
                 forvar2299,
                 reg2295,
                 reg2294,
                 reg2289,
                 reg2288,
                 reg2284,
                 reg2280,
                 reg2278,
                 reg2277,
                 reg2275,
                 reg2272,
                 forvar2265,
                 forvar2262,
                 reg2261,
                 reg2259,
                 reg2258,
                 reg2257,
                 reg2256,
                 reg2236,
                 reg2254,
                 reg2253,
                 reg2252,
                 reg2251,
                 reg2250,
                 reg2249,
                 reg2245,
                 reg2244,
                 reg2243,
                 reg2241,
                 reg2240,
                 reg2239,
                 reg2238,
                 reg2237,
                 forvar2236,
                 reg2233,
                 reg2231,
                 reg2229,
                 reg2227,
                 reg2226,
                 forvar2214,
                 reg2212,
                 forvar2220,
                 reg2219,
                 reg2218,
                 reg2214,
                 forvar2212,
                 reg2211,
                 reg2210,
                 reg2208,
                 reg2207,
                 forvar2206,
                 reg2205,
                 reg2204,
                 reg2201,
                 reg2200,
                 forvar2198,
                 forvar2197,
                 reg1368,
                 reg1367,
                 forvar1366,
                 reg1364,
                 reg1363,
                 reg1361,
                 forvar1360,
                 reg1358,
                 reg1356,
                 forvar1354,
                 reg1331,
                 forvar1330,
                 reg1350,
                 forvar1348,
                 reg1342,
                 reg1341,
                 reg1340,
                 reg1337,
                 reg1336,
                 reg1334,
                 reg1332,
                 forvar1331,
                 reg1330,
                 reg1329,
                 reg1058,
                 reg1056,
                 reg1055,
                 reg1053,
                 reg1051,
                 reg1049,
                 reg1048,
                 reg1045,
                 reg1042,
                 reg1041,
                 forvar1040,
                 reg1039,
                 reg1038,
                 reg1037,
                 forvar1035,
                 reg1034,
                 forvar1033,
                 reg1032,
                 reg1031,
                 reg1030,
                 reg1029,
                 reg1028,
                 forvar1027,
                 reg1026,
                 forvar1024,
                 reg1022,
                 reg1021,
                 reg1019,
                 reg1018,
                 forvar1017,
                 reg1016,
                 reg1015,
                 forvar1014,
                 reg1012,
                 reg1011,
                 forvar1003,
                 forvar999,
                 reg1008,
                 reg1007,
                 reg1006,
                 reg1004,
                 reg1003,
                 forvar1002,
                 reg1000,
                 reg999,
                 reg998,
                 reg993,
                 reg992,
                 reg987,
                 reg984,
                 reg983,
                 forvar980,
                 forvar977,
                 reg975,
                 reg974,
                 reg973,
                 reg971,
                 reg969,
                 reg968,
                 reg967,
                 reg965,
                 forvar961,
                 reg960,
                 reg958,
                 reg954,
                 reg953,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 forvar946,
                 forvar942,
                 forvar929,
                 reg939,
                 reg938,
                 reg937,
                 forvar936,
                 reg935,
                 reg934,
                 reg930,
                 reg929,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((({((wire924 ? wire926 : wire926) ? (-wire925) : (^wire928))} ?
              $signed(wire927[(3'h6):(3'h4)]) : (-(&wire924[(4'h8):(2'h3)]))) ?
          (|wire925) : {$signed({wire927[(2'h2):(2'h2)]}),
              wire926[(4'h8):(3'h4)]}))
        begin
          if ({wire926[(2'h3):(2'h2)],
              {{$unsigned((-wire924)), (^~wire925)},
                  $unsigned(({wire927, wire928} == wire924[(1'h1):(1'h0)])),
                  wire927},
              $unsigned((~^wire927))})
            begin
              reg929 = $signed((|$unsigned({wire924[(4'hb):(4'h8)],
                  wire925,
                  (wire928 ? wire926 : (7'h4c))})));
              reg930 = $signed($unsigned(wire928[(5'h11):(2'h3)]));
              reg931 <= $signed(wire926[(1'h1):(1'h1)]);
              reg932 <= reg930;
              reg933 <= (reg930 ?
                  reg929[(4'h9):(4'h8)] : (reg931[(5'h1a):(5'h19)] | wire924));
              reg934 = $signed((|($signed(reg932[(3'h6):(3'h4)]) != $unsigned((+(8'ha3))))));
            end
          else
            begin
              reg929 = (~|(7'h47));
            end
          reg935 = wire924;
          for (forvar936 = (1'h0); (forvar936 < (1'h0)); forvar936 = (forvar936 + (1'h1)))
            begin
              reg937 = (((7'h4c) >= (|$signed($unsigned(wire928)))) && ($signed((&(reg935 || reg933))) != (8'hbc)));
              reg938 = $unsigned(((wire925 && ((&reg934) ?
                      reg937[(1'h1):(1'h0)] : (wire926 ? reg935 : reg931))) ?
                  ($signed((wire924 >>> wire927)) ?
                      {reg935,
                          $signed(wire925)} : (reg931 >> (wire927 > reg930))) : ($signed($signed(wire928)) | (~&(reg929 ~^ wire926)))));
              reg939 = wire926[(1'h0):(1'h0)];
            end
        end
      else
        begin
          for (forvar929 = (1'h0); (forvar929 < (3'h6)); forvar929 = (forvar929 + (1'h1)))
            begin
              reg930 = wire924[(4'hc):(4'ha)];
              reg931 <= reg931[(3'h5):(2'h3)];
              reg932 <= (^~(&$unsigned($signed((reg929 ? reg931 : reg939)))));
              reg933 <= (~^(($signed((reg929 ?
                      forvar936 : reg937)) <= $unsigned(wire926[(4'h8):(3'h6)])) ?
                  $unsigned(wire925) : ((~reg937) ?
                      {(8'hb7),
                          (reg935 ?
                              forvar929 : wire924)} : $unsigned($unsigned(reg937)))));
              reg936 <= reg939;
              reg940 <= {$unsigned(($signed(wire926) != ((&reg934) >= (wire928 != (7'h4e))))),
                  (reg930[(5'h15):(1'h1)] - $unsigned({((8'ha3) - reg936),
                      $unsigned(reg930)})),
                  (wire926 ?
                      $signed((~|(8'hba))) : $signed(($unsigned(wire925) >>> (+wire926))))};
              reg941 <= reg937;
            end
          for (forvar942 = (1'h0); (forvar942 < (3'h5)); forvar942 = (forvar942 + (1'h1)))
            begin
              reg943 <= forvar936;
            end
          reg944 <= forvar942;
          reg945 <= reg930[(3'h4):(3'h4)];
        end
      for (forvar946 = (1'h0); (forvar946 < (2'h2)); forvar946 = (forvar946 + (1'h1)))
        begin
          reg947 = $unsigned($unsigned(reg941));
          if (($signed(((|$signed(reg945)) <<< (reg929[(2'h2):(2'h2)] ?
              $signed(reg943) : $signed((8'hb6))))) > reg938))
            begin
              reg948 = (^$signed((+{$signed(reg939), (forvar946 & reg934)})));
              reg949 = $signed({forvar929});
              reg950 = {$unsigned($unsigned($signed((~&reg929)))), reg948};
              reg951 = {wire926[(1'h0):(1'h0)],
                  ($unsigned($signed({forvar929,
                      forvar936,
                      (7'h4a)})) <= ($unsigned(reg936) ?
                      reg947[(5'h19):(3'h4)] : {(reg938 != reg936)})),
                  (+$unsigned($signed((wire926 ? reg932 : (7'h46)))))};
              reg952 <= ($unsigned(($signed(((8'h9e) && reg948)) ?
                      $signed((8'ha5)) : (reg935 ?
                          (+reg933) : (reg937 ? forvar936 : wire927)))) ?
                  reg938 : reg947[(2'h3):(1'h1)]);
            end
          else
            begin
              reg952 <= $signed(forvar936);
              reg953 = forvar936;
              reg954 = forvar942[(3'h5):(3'h4)];
              reg955 <= $unsigned((~(^$unsigned(reg934))));
              reg956 <= {($unsigned((~|$unsigned(reg939))) ?
                      $signed($unsigned(reg954[(3'h6):(3'h6)])) : (^~$signed({reg932,
                          reg941,
                          wire926}))),
                  ($unsigned((reg947 || forvar936[(5'h14):(4'h9)])) ^ $unsigned(reg951)),
                  reg930};
              reg957 <= (wire926[(2'h3):(2'h2)] << (|{reg944}));
            end
        end
      if ($signed(reg941[(5'h12):(4'hb)]))
        begin
          reg958 = ($unsigned($unsigned($signed($signed(reg934)))) ^~ reg945[(4'ha):(3'h4)]);
          reg959 <= forvar946;
          reg960 = reg947;
          for (forvar961 = (1'h0); (forvar961 < (2'h3)); forvar961 = (forvar961 + (1'h1)))
            begin
              reg962 <= (8'h9f);
              reg963 <= ($signed(($signed($signed(reg934)) & reg954)) > {reg954,
                  $signed($signed({reg931, reg951, reg958}))});
              reg964 <= (~|reg931[(4'h9):(4'h9)]);
              reg965 = (($signed(($unsigned(reg953) >= (&reg930))) ~^ {((reg935 ?
                              (7'h52) : (8'ha1)) ?
                          ((7'h4f) ? reg940 : reg963) : $signed(reg933))}) ?
                  reg936[(4'he):(3'h4)] : $unsigned(reg951[(5'h13):(5'h13)]));
              reg966 <= (+reg929);
              reg967 = $signed((8'hb7));
            end
          if ($signed(({reg950, reg956} ?
              ($signed((~|(7'h44))) ?
                  $unsigned((reg966 | reg949)) : $unsigned((reg965 >> reg952))) : $signed(reg932))))
            begin
              reg968 = reg930;
              reg969 = $signed(reg967[(2'h2):(1'h1)]);
              reg970 <= (((&reg951[(5'h19):(4'he)]) + $unsigned($unsigned($signed(reg951)))) | reg940[(4'he):(3'h6)]);
              reg971 = reg932;
            end
          else
            begin
              reg970 <= reg932;
              reg972 <= reg952;
              reg973 = $signed({($unsigned($signed(reg929)) ?
                      (reg954 == (reg953 ?
                          (8'hbb) : forvar961)) : $unsigned(reg955)),
                  $signed((reg950 < $signed(reg970)))});
              reg974 = (reg955 | $unsigned(((&(reg949 >>> reg940)) ^ ({(7'h52),
                      reg931} ?
                  (reg929 >> reg945) : $signed(reg940)))));
              reg975 = forvar961;
              reg976 <= $unsigned((8'hb9));
            end
        end
      else
        begin
          reg959 <= {(^~(($signed(reg934) < $signed((7'h56))) ?
                  reg952 : {{reg931}}))};
          reg961 <= reg970;
          if (forvar936[(4'hc):(4'h9)])
            begin
              reg965 = ($unsigned(reg975) | (|(7'h4d)));
              reg967 = $unsigned({($unsigned((~&(8'had))) ?
                      ((reg948 ?
                          reg932 : (8'haa)) * reg974[(3'h7):(3'h7)]) : (!(forvar942 - reg970))),
                  (7'h42)});
            end
          else
            begin
              reg965 = (~|(^$unsigned((reg970 >> $unsigned(wire925)))));
              reg966 <= reg971[(5'h16):(4'hf)];
              reg967 = $unsigned($unsigned((7'h51)));
              reg970 <= (reg941[(4'ha):(3'h6)] ?
                  {reg935, (^~forvar946)} : reg956[(1'h1):(1'h1)]);
              reg972 <= {(~$unsigned((+(wire924 ? (8'ha0) : reg934))))};
              reg973 = (((-$unsigned(reg966[(4'hf):(3'h6)])) >= (~&$unsigned(reg939[(4'hf):(4'h8)]))) > reg938);
            end
          reg976 <= $unsigned((((^~wire927) || $unsigned((&(8'hb5)))) ?
              ((~&reg955) | reg933) : reg944));
        end
      for (forvar977 = (1'h0); (forvar977 < (3'h5)); forvar977 = (forvar977 + (1'h1)))
        begin
          reg978 <= ($unsigned($unsigned((~&(^(8'haa))))) ~^ $unsigned($signed((8'haa))));
          reg979 <= $unsigned(reg949[(4'ha):(2'h3)]);
          for (forvar980 = (1'h0); (forvar980 < (3'h4)); forvar980 = (forvar980 + (1'h1)))
            begin
              reg981 <= ({($signed((reg963 ?
                          (8'hbe) : reg938)) << (~^$signed((8'hb0)))),
                      (|$signed(reg936[(3'h7):(2'h3)])),
                      $signed($signed($unsigned(reg974)))} ?
                  (|(((reg930 ? forvar946 : reg978) ?
                          ((8'hb2) * reg950) : (reg940 ? reg959 : forvar929)) ?
                      (8'hb8) : $unsigned((reg973 <= reg972)))) : $signed(((^reg952) ^ {(|forvar942)})));
              reg982 <= (((((reg966 <= forvar936) >= (forvar980 ?
                      reg948 : reg956)) ^~ $unsigned((^~wire928))) ?
                  (((reg973 << forvar946) & reg940[(4'h8):(1'h0)]) ?
                      ($signed(reg962) < (reg949 ^~ reg948)) : ((|reg955) ^ reg964)) : $signed({reg941})) <<< (|{reg969,
                  wire924,
                  (reg976 ? $signed(reg965) : (reg981 != reg931))}));
              reg983 = forvar977[(3'h7):(3'h6)];
              reg984 = reg978;
            end
          reg985 <= reg974;
          reg986 <= $signed((&(8'hb1)));
          if (($unsigned((((reg941 + (8'hae)) ^ (8'ha4)) ?
              ({reg970} + $unsigned(reg953)) : reg945)) >= $unsigned({$unsigned((reg972 ?
                  reg986 : reg979)),
              $signed((reg975 ? reg948 : reg950)),
              $unsigned(reg953[(2'h3):(2'h3)])})))
            begin
              reg987 = $signed(reg941[(4'h8):(3'h5)]);
              reg988 <= ((($signed(reg957[(5'h13):(5'h13)]) > $unsigned(reg961)) ?
                      (~&reg933[(2'h3):(2'h3)]) : $unsigned((((7'h41) ?
                          wire924 : reg972) || reg950))) ?
                  reg937 : ((^~reg964[(2'h2):(2'h2)]) > (~|reg966)));
              reg989 <= ((($unsigned($signed(reg975)) + (~^{reg955})) >>> ((~^(~reg932)) ?
                      (forvar936 ?
                          (reg934 ?
                              reg983 : reg957) : $signed(wire926)) : forvar980)) ?
                  reg933 : ({reg973[(4'hf):(3'h6)]} ?
                      (+(reg948 ?
                          reg938 : $unsigned(reg964))) : ($unsigned(reg982) << ((~|forvar980) ?
                          $signed(reg962) : $unsigned(wire924)))));
              reg990 <= {(~^reg973), reg968[(1'h0):(1'h0)]};
              reg991 <= (~^reg964);
            end
          else
            begin
              reg987 = reg959;
              reg992 = ((8'haa) ^~ (&(!$unsigned((reg989 ?
                  (7'h4e) : reg959)))));
              reg993 = (reg969 ?
                  (|$unsigned($signed((reg975 ?
                      reg934 : reg970)))) : {$signed(reg931)});
              reg994 <= ((reg985[(5'h10):(4'h8)] < (&((~&reg945) ?
                  reg962[(3'h5):(3'h4)] : (reg992 ?
                      reg954 : (7'h40))))) != $signed({($signed(wire924) ?
                      reg949[(4'ha):(4'h9)] : (reg958 <= reg938)),
                  $signed($unsigned(reg929)),
                  reg970}));
            end
        end
      if (reg983[(1'h1):(1'h0)])
        begin
          if ((((!forvar946[(4'he):(2'h3)]) ?
                  (reg956 ?
                      wire924 : {{reg956, reg950},
                          reg933[(1'h0):(1'h0)],
                          (!reg941)}) : $unsigned({(reg936 >> reg974),
                      {reg940}})) ?
              (({(reg985 ? reg964 : (7'h41))} ?
                  $signed($unsigned(reg929)) : ($unsigned(reg988) ?
                      reg951 : $unsigned((8'hb1)))) < wire928) : (($signed((reg972 ?
                      reg958 : reg994)) - ((~&(8'hbb)) ?
                      reg931[(4'ha):(3'h7)] : reg949)) ?
                  (($signed(forvar929) ? $signed(reg948) : $unsigned(reg981)) ?
                      forvar942[(4'hf):(4'hc)] : $signed((reg993 + reg990))) : (8'ha6))))
            begin
              reg995 <= reg958;
              reg996 <= forvar980[(1'h1):(1'h1)];
              reg997 <= (!($signed(reg970) & reg990));
            end
          else
            begin
              reg998 = reg995[(1'h1):(1'h0)];
              reg999 = (7'h56);
              reg1000 = {$unsigned((+(!reg957)))};
              reg1001 <= (~^{(-reg991), (~^reg968), forvar961});
            end
          for (forvar1002 = (1'h0); (forvar1002 < (2'h2)); forvar1002 = (forvar1002 + (1'h1)))
            begin
              reg1003 = (~((+(~|$signed(reg968))) ?
                  $signed(reg955[(4'hb):(3'h4)]) : (wire928 && ((8'ha4) != (reg994 ?
                      (7'h58) : reg1000)))));
              reg1004 = ($unsigned(reg932) ^ reg952);
              reg1005 <= $unsigned($unsigned(reg974));
              reg1006 = $unsigned($unsigned($signed(reg963[(1'h0):(1'h0)])));
              reg1007 = (~|reg1000[(4'hc):(3'h5)]);
              reg1008 = (~(($unsigned((~^reg941)) ?
                  $unsigned(reg990[(5'h13):(3'h6)]) : reg983) != {$unsigned(reg962)}));
              reg1009 <= (+(({reg992, $signed(reg951)} ?
                      ($unsigned((8'hb6)) - (^~wire925)) : ($signed(reg1007) < forvar942)) ?
                  reg959 : $unsigned(reg985[(4'hd):(4'hb)])));
            end
          reg1010 <= (+$unsigned($unsigned({reg973[(5'h10):(4'hb)]})));
        end
      else
        begin
          reg998 = (^~(reg935 ?
              $signed(reg986[(4'hb):(4'ha)]) : $signed($signed((^forvar942)))));
          for (forvar999 = (1'h0); (forvar999 < (2'h3)); forvar999 = (forvar999 + (1'h1)))
            begin
              reg1000 = $unsigned(reg967[(2'h3):(2'h3)]);
              reg1001 <= $unsigned(reg935[(1'h1):(1'h1)]);
              reg1002 <= reg930[(4'hf):(4'hc)];
            end
          for (forvar1003 = (1'h0); (forvar1003 < (3'h4)); forvar1003 = (forvar1003 + (1'h1)))
            begin
              reg1005 <= (reg954 <<< $unsigned($unsigned($signed($unsigned((8'h9e))))));
              reg1006 = reg1003;
              reg1007 = (reg953 ?
                  $signed(forvar936[(3'h5):(2'h2)]) : ({$signed(forvar961),
                      reg950[(1'h0):(1'h0)]} - forvar1003));
              reg1009 <= (~reg1000[(1'h0):(1'h0)]);
              reg1011 = $signed($signed($signed(reg985)));
            end
        end
      reg1012 = $unsigned(($signed(((+reg936) ?
          $unsigned(reg948) : $signed(reg947))) <= {((reg982 ?
                  reg944 : forvar980) ?
              (~&reg997) : $signed(reg952)),
          ((+forvar942) ? ((8'ha2) ? (8'hab) : (8'hac)) : {reg960})}));
    end
  assign wire1013 = (8'haf);
  always
    @(posedge clk) begin
      for (forvar1014 = (1'h0); (forvar1014 < (3'h4)); forvar1014 = (forvar1014 + (1'h1)))
        begin
          reg1015 = (({(-{reg964, reg979, reg931}),
                      {reg996[(4'hd):(1'h0)],
                          $signed((8'hb8)),
                          (reg931 ? reg936 : reg990)}} ?
                  reg940[(3'h6):(2'h2)] : (reg1005[(4'h8):(3'h6)] ?
                      ((|reg1009) <<< {(7'h55), forvar1014, (8'ha1)}) : {reg997,
                          (^~reg1010)})) ?
              (-reg1001[(5'h18):(2'h2)]) : (~reg988[(1'h0):(1'h0)]));
          reg1016 = (&(~((^~reg996) ~^ reg1002)));
        end
      for (forvar1017 = (1'h0); (forvar1017 < (3'h5)); forvar1017 = (forvar1017 + (1'h1)))
        begin
          reg1018 = (!(reg944[(1'h0):(1'h0)] ?
              ($unsigned(reg1001) >> (-(reg1010 ?
                  reg1002 : (8'hac)))) : {wire927, reg1015[(2'h2):(1'h1)]}));
          if ((~^reg997))
            begin
              reg1019 = reg1018;
            end
          else
            begin
              reg1020 <= $signed(({reg976[(5'h11):(1'h0)]} > {$unsigned(reg962[(1'h0):(1'h0)])}));
              reg1021 = (-(~^(((reg961 * reg1005) ?
                  (-reg957) : $signed(reg936)) >> reg982)));
              reg1022 = ({reg963[(3'h6):(3'h6)]} <<< reg932);
            end
          reg1023 <= (~&$signed(forvar1014[(3'h6):(3'h4)]));
          for (forvar1024 = (1'h0); (forvar1024 < (1'h0)); forvar1024 = (forvar1024 + (1'h1)))
            begin
              reg1025 <= $unsigned((|((reg1005[(3'h7):(3'h4)] == ((8'hbe) ?
                      reg994 : reg945)) ?
                  $signed(reg943[(5'h15):(5'h12)]) : forvar1024[(2'h2):(1'h0)])));
              reg1026 = ($signed({(!(8'ha7)), $signed($unsigned((7'h53)))}) ?
                  (-$signed(reg933)) : $signed({($unsigned(reg1001) ?
                          $unsigned(reg976) : {reg1009, reg997, reg986}),
                      $signed((reg976 ^ reg945))}));
            end
          for (forvar1027 = (1'h0); (forvar1027 < (3'h4)); forvar1027 = (forvar1027 + (1'h1)))
            begin
              reg1028 = ((+$unsigned(reg943)) ?
                  reg955 : (reg997 ?
                      {$signed((reg955 > reg997)),
                          reg1005[(2'h3):(2'h2)],
                          $unsigned((+(7'h43)))} : $signed(reg1005[(3'h4):(3'h4)])));
              reg1029 = ($unsigned($unsigned(reg1019)) ?
                  $signed($unsigned((+$unsigned(wire928)))) : {({(reg944 ?
                                  reg1010 : reg1018),
                              {reg956, reg1010},
                              wire925[(3'h5):(2'h2)]} ?
                          (~^$unsigned(reg1016)) : $unsigned((reg933 ?
                              reg932 : (7'h54))))});
              reg1030 = ($unsigned(($signed((reg941 < reg1016)) ?
                  (^~$signed(reg961)) : {(reg1023 ? (8'hb7) : reg985),
                      $signed(reg991),
                      reg964[(1'h0):(1'h0)]})) != ((~^$signed($signed(reg978))) && $unsigned($unsigned((reg941 < reg976)))));
            end
          reg1031 = reg976[(5'h12):(4'he)];
        end
    end
  always
    @(posedge clk) begin
      reg1032 = $unsigned(reg996[(2'h3):(2'h2)]);
      for (forvar1033 = (1'h0); (forvar1033 < (1'h0)); forvar1033 = (forvar1033 + (1'h1)))
        begin
          reg1034 = reg1002[(4'hc):(4'hc)];
          for (forvar1035 = (1'h0); (forvar1035 < (1'h0)); forvar1035 = (forvar1035 + (1'h1)))
            begin
              reg1036 <= reg963[(3'h7):(3'h5)];
              reg1037 = (^(({$signed(reg952), $signed(reg991)} ?
                      $signed({reg1010, reg933}) : $signed({reg994,
                          (7'h50),
                          reg989})) ?
                  (($unsigned(reg976) ?
                      $signed(reg985) : $signed(reg976)) & (wire1013 ?
                      reg981[(3'h4):(2'h2)] : (~reg966))) : (^{reg940[(4'ha):(2'h3)]})));
              reg1038 = (^~reg1025);
              reg1039 = (~^reg1002[(5'h1d):(4'hc)]);
            end
          for (forvar1040 = (1'h0); (forvar1040 < (3'h6)); forvar1040 = (forvar1040 + (1'h1)))
            begin
              reg1041 = reg1010;
              reg1042 = $unsigned($signed(reg966));
              reg1043 <= reg933[(2'h2):(1'h0)];
              reg1044 <= ({$signed({(reg957 ? reg1041 : reg932),
                      (reg1010 ? reg989 : reg981),
                      reg963}),
                  $unsigned($signed($signed(reg979))),
                  ($signed(reg936[(3'h4):(3'h4)]) < (~|$signed(reg1038)))} - (reg961 + reg940[(3'h6):(1'h1)]));
            end
          if (({$unsigned(((reg1043 ? (8'haf) : reg978) ?
                      $signed((7'h42)) : (|wire927)))} ?
              ((reg933 ?
                  forvar1035[(1'h1):(1'h1)] : ((reg978 << forvar1040) <<< (-reg1020))) < (reg931 && reg945)) : (8'ha3)))
            begin
              reg1045 = $signed($signed(reg982));
              reg1046 <= (7'h44);
            end
          else
            begin
              reg1046 <= (8'ha3);
              reg1047 <= reg982[(4'hd):(3'h7)];
              reg1048 = $signed($unsigned($unsigned({{reg1032, reg943},
                  (!forvar1040),
                  $signed(reg964)})));
              reg1049 = $unsigned(($unsigned((!reg989)) ?
                  {reg940,
                      $signed((reg994 | reg1045)),
                      reg943[(4'h9):(3'h5)]} : ((!reg1002) ?
                      (&(^~reg932)) : reg976[(5'h11):(1'h0)])));
              reg1050 <= ($signed($unsigned({(8'ha8)})) ?
                  reg963 : (~|$unsigned($signed((~&reg1002)))));
              reg1051 = (&(^~(reg1041[(4'hb):(3'h5)] ?
                  reg1050 : ($unsigned(reg996) ? reg995 : reg982))));
            end
          if ($unsigned(reg1020[(4'hd):(1'h1)]))
            begin
              reg1052 <= $signed($unsigned($signed({$unsigned((8'hba)),
                  (reg1010 > reg943),
                  $signed(reg955)})));
              reg1053 = forvar1033[(2'h2):(1'h0)];
              reg1054 <= ((!reg941) & ((($signed(reg1009) ?
                  (+reg988) : (!reg940)) > ((reg1051 != (8'hbd)) ?
                  (reg943 ? reg982 : reg990) : $unsigned(reg982))) * (7'h57)));
              reg1055 = $signed(reg940);
              reg1056 = reg964[(2'h2):(2'h2)];
            end
          else
            begin
              reg1053 = $unsigned($unsigned((!((-reg961) ?
                  {reg997, reg961, reg1047} : reg1055[(4'h8):(2'h3)]))));
              reg1055 = reg933[(2'h3):(1'h1)];
              reg1056 = $signed((!({$unsigned(reg1052), {forvar1035}} ?
                  (reg1010 << (reg959 <<< reg1042)) : ((~|(7'h4d)) != $signed(reg972)))));
              reg1057 <= (^~(&reg940[(2'h3):(2'h3)]));
            end
          reg1058 = $unsigned({{$signed($unsigned(reg962))}});
        end
    end
  module1059 #() modinst1328 (wire1327, clk, reg982, reg1002, reg931, reg956, reg932);
  always
    @(posedge clk) begin
      reg1329 = $signed({(~&reg1052[(5'h10):(1'h1)]),
          reg931,
          (reg963 ? reg1057 : ($unsigned((7'h40)) & $signed(reg1054)))});
      if (((^~(reg931 ?
              ((|reg997) - (&reg1054)) : ($unsigned(reg1001) ?
                  $signed(reg976) : (|reg976)))) ?
          $signed(((~&(!wire925)) < $unsigned($signed(wire925)))) : $signed($signed((8'h9c)))))
        begin
          reg1330 = {reg1025[(4'hc):(1'h1)],
              (&reg979),
              ((~^reg957) ?
                  reg996[(3'h6):(3'h6)] : {wire1327[(5'h15):(4'h8)],
                      ((^~reg932) ? reg1054 : reg991[(1'h0):(1'h0)]),
                      ((8'hb1) ? $unsigned(reg962) : (reg962 | reg933))})};
          for (forvar1331 = (1'h0); (forvar1331 < (3'h6)); forvar1331 = (forvar1331 + (1'h1)))
            begin
              reg1332 = (~&wire926[(2'h3):(1'h0)]);
              reg1333 <= ($unsigned($unsigned($unsigned({reg1047}))) - $signed(($unsigned((~^(8'hae))) ?
                  reg966 : ({reg944} ?
                      reg931[(4'ha):(4'ha)] : ((7'h50) ? wire1327 : reg944)))));
              reg1334 = (^~($unsigned(reg988[(1'h1):(1'h0)]) ~^ (~&(!{reg1333,
                  reg959}))));
            end
          reg1335 <= $unsigned(reg1052);
          if ({reg997[(4'hb):(4'h8)]})
            begin
              reg1336 = $unsigned($unsigned(reg997[(5'h15):(5'h13)]));
              reg1337 = $unsigned((~^{((reg1005 ?
                      reg1057 : reg994) ~^ $signed(reg957)),
                  $unsigned(reg991[(1'h0):(1'h0)]),
                  $signed($unsigned(reg932))}));
              reg1338 <= reg1001[(3'h6):(1'h0)];
              reg1339 <= (((8'hb7) <<< reg988) ?
                  reg963 : ((~^reg1050[(1'h1):(1'h1)]) ?
                      reg979 : $signed($signed($signed(reg966)))));
            end
          else
            begin
              reg1338 <= $signed((|(^~(reg1036[(2'h2):(1'h1)] && (reg944 ?
                  reg1050 : (7'h4e))))));
              reg1340 = (~$unsigned(reg972[(4'h9):(3'h6)]));
              reg1341 = $unsigned((~&(~^reg982)));
              reg1342 = (((|reg931) ?
                  $signed($signed({(8'ha5),
                      reg990,
                      reg1036})) : ({reg952[(4'h9):(2'h2)],
                          $unsigned(reg1339),
                          wire926} ?
                      reg985[(5'h13):(1'h0)] : (~(^reg1338)))) * $unsigned((reg964[(1'h0):(1'h0)] & $unsigned(reg1001))));
              reg1343 <= reg961;
              reg1344 <= (~|{{$signed(reg972)}});
              reg1345 <= $signed(($signed($unsigned(((8'h9f) && reg961))) ?
                  reg991 : (8'hbb)));
            end
          reg1346 <= {reg957};
          reg1347 <= reg1335[(4'hd):(4'h8)];
          for (forvar1348 = (1'h0); (forvar1348 < (1'h1)); forvar1348 = (forvar1348 + (1'h1)))
            begin
              reg1349 <= reg1332[(5'h15):(4'h8)];
              reg1350 = wire924[(1'h1):(1'h1)];
              reg1351 <= ((({(reg945 ? (8'hb1) : reg1046)} ?
                  reg1330[(5'h14):(2'h3)] : $unsigned(reg1342)) == ($signed((reg1002 < reg944)) ?
                  $unsigned((reg1333 == reg988)) : (reg943[(1'h0):(1'h0)] ?
                      (reg963 * reg1047) : reg1009))) - reg955);
              reg1352 <= $unsigned((~^({(reg991 > reg996), $unsigned(reg1330)} ?
                  $unsigned((^~reg1330)) : reg1343)));
            end
        end
      else
        begin
          for (forvar1330 = (1'h0); (forvar1330 < (3'h4)); forvar1330 = (forvar1330 + (1'h1)))
            begin
              reg1331 = ((((&$unsigned(reg981)) ?
                  $unsigned((reg1347 ? reg944 : (8'had))) : {(7'h55),
                      (+reg1338),
                      ((7'h50) ? forvar1348 : reg932)}) + $unsigned(((reg1334 ?
                      reg932 : wire927) ?
                  forvar1330 : (reg1052 || reg985)))) >> (8'ha5));
              reg1333 <= reg991[(1'h0):(1'h0)];
              reg1334 = $signed(reg1044[(4'h8):(3'h4)]);
              reg1335 <= (^$unsigned(forvar1331));
              reg1336 = reg990;
              reg1338 <= (^((8'h9c) ?
                  ($signed((reg995 ^~ reg1025)) ?
                      reg963 : (((8'ha3) ?
                          reg1342 : reg986) >> reg1329)) : ({reg933[(1'h1):(1'h1)]} >> reg1329[(4'hd):(4'hb)])));
            end
          if (forvar1330[(4'h9):(3'h4)])
            begin
              reg1339 <= $signed(reg932[(3'h7):(1'h1)]);
              reg1340 = $signed(((($signed((8'hb1)) ?
                          reg995[(2'h3):(1'h1)] : $unsigned((7'h4a))) ?
                      (((8'ha6) ? (7'h4c) : (8'hab)) ?
                          (reg1352 || (8'hb1)) : reg970[(4'h9):(2'h3)]) : (^~(&reg989))) ?
                  (~^({(8'hb6)} >>> reg1340[(4'he):(3'h6)])) : (&reg1054[(4'hc):(4'h9)])));
            end
          else
            begin
              reg1340 = reg990;
              reg1343 <= reg986;
              reg1344 <= (^~($signed(($signed(reg985) != forvar1330)) ?
                  reg941 : reg1010[(4'ha):(3'h5)]));
              reg1345 <= ((~reg1352) == forvar1331);
            end
        end
      reg1353 <= (reg1052 > (^$signed({$unsigned(reg991),
          (reg991 ? (7'h4f) : (8'hb9)),
          reg1330[(4'h9):(3'h5)]})));
    end
  always
    @(posedge clk) begin
      for (forvar1354 = (1'h0); (forvar1354 < (2'h3)); forvar1354 = (forvar1354 + (1'h1)))
        begin
          reg1355 <= reg997[(5'h12):(5'h11)];
          if ($unsigned(reg932[(3'h7):(2'h3)]))
            begin
              reg1356 = $unsigned(($signed(reg963) + (~{reg1355[(5'h1b):(2'h2)],
                  {forvar1354, reg989, reg1343},
                  $signed((7'h53))})));
            end
          else
            begin
              reg1357 <= $signed($unsigned(reg952));
              reg1358 = $unsigned(((reg990[(4'hc):(3'h5)] ?
                  reg1020 : $signed($signed(reg940))) + $unsigned(reg985)));
              reg1359 <= ((^reg1357[(3'h4):(2'h2)]) != $unsigned(reg1353[(3'h6):(3'h6)]));
            end
          for (forvar1360 = (1'h0); (forvar1360 < (1'h0)); forvar1360 = (forvar1360 + (1'h1)))
            begin
              reg1361 = ($signed($signed(reg981)) ?
                  (&reg1339) : ({$unsigned($unsigned(wire927))} >> (|reg1005[(4'he):(4'h8)])));
              reg1362 <= ((~|reg1343) + ((($signed(wire924) & (!reg1358)) ?
                      ((reg1353 ?
                          reg1335 : reg952) ^ {reg1358}) : {(reg989 <= wire927),
                          {reg963, reg944},
                          (~reg1352)}) ?
                  reg961[(3'h7):(3'h7)] : reg962));
              reg1363 = reg962;
              reg1364 = $signed({reg1009});
              reg1365 <= ((({reg981} ?
                      ((~&(8'hba)) ?
                          (~^reg1057) : wire924) : {$unsigned(reg1346),
                          reg963[(2'h3):(2'h2)]}) ?
                  ((((8'ha5) ?
                      (7'h4f) : reg957) ^ reg1363) ^ (((8'hb8) | reg1346) ?
                      $unsigned(reg994) : (reg1355 < wire927))) : $unsigned({$signed((8'h9f)),
                      reg933[(2'h2):(2'h2)]})) ^~ $unsigned((((8'hae) ?
                  $signed(reg997) : reg1363[(4'h8):(1'h1)]) == ((|reg976) ?
                  reg982 : $signed(reg1335)))));
            end
          for (forvar1366 = (1'h0); (forvar1366 < (1'h0)); forvar1366 = (forvar1366 + (1'h1)))
            begin
              reg1367 = (((~|($unsigned(reg1357) ? reg1046 : (-reg1050))) ?
                      reg1025 : $unsigned(wire924[(4'hf):(3'h7)])) ?
                  ($unsigned(reg991) ?
                      reg1057[(3'h7):(3'h5)] : {reg1364}) : $signed($signed(reg1364[(3'h5):(1'h1)])));
              reg1368 = (~&(~|reg1046));
              reg1369 <= reg1047;
              reg1370 <= reg1054[(3'h5):(1'h0)];
              reg1371 <= {(reg991 || wire926[(3'h6):(3'h6)])};
              reg1372 <= reg1352;
            end
          reg1373 <= {($signed({$unsigned(reg996)}) << $signed($unsigned((reg1364 ?
                  reg1043 : reg1372))))};
          reg1374 <= ((~&wire928[(5'h10):(4'he)]) <<< (8'hbd));
        end
    end
  always
    @(posedge clk) begin
      reg1375 <= $signed((|(|$signed(reg961))));
    end
  module1376 #() modinst1771 (.y(wire1770), .clk(clk), .wire1380(reg1374), .wire1381(wire924), .wire1378(reg994), .wire1379(reg1362), .wire1377(reg1050));
  assign wire1772 = reg1005[(1'h1):(1'h0)];
  module1773 #() modinst2196 (.y(wire2195), .clk(clk), .wire1775(reg936), .wire1778(reg1357), .wire1776(reg994), .wire1774(reg1010), .wire1777(reg1005));
  always
    @(posedge clk) begin
      for (forvar2197 = (1'h0); (forvar2197 < (3'h5)); forvar2197 = (forvar2197 + (1'h1)))
        begin
          for (forvar2198 = (1'h0); (forvar2198 < (2'h2)); forvar2198 = (forvar2198 + (1'h1)))
            begin
              reg2199 <= $signed(reg997);
              reg2200 = $unsigned($unsigned((^$unsigned((reg956 ?
                  reg1371 : reg1353)))));
              reg2201 = reg1345;
              reg2202 <= $unsigned((wire1013 ?
                  $unsigned($unsigned($signed(reg1374))) : (-wire1327)));
              reg2203 <= reg1355[(5'h11):(1'h0)];
              reg2204 = {(reg991 ?
                      (8'hb7) : (~|(forvar2198 ?
                          $signed(reg931) : $unsigned(reg996))))};
              reg2205 = $signed(reg1036[(3'h7):(2'h3)]);
            end
          for (forvar2206 = (1'h0); (forvar2206 < (3'h5)); forvar2206 = (forvar2206 + (1'h1)))
            begin
              reg2207 = wire1013[(3'h4):(2'h3)];
              reg2208 = {forvar2198};
              reg2209 <= forvar2206;
              reg2210 = reg1046;
            end
          reg2211 = $signed(reg1050[(4'hf):(4'hc)]);
        end
      if (($unsigned((+reg1338[(4'ha):(3'h7)])) ?
          reg961[(4'hb):(2'h3)] : reg991[(1'h1):(1'h1)]))
        begin
          for (forvar2212 = (1'h0); (forvar2212 < (2'h2)); forvar2212 = (forvar2212 + (1'h1)))
            begin
              reg2213 <= $signed({(({reg991, (8'h9f)} << ((7'h52) >> reg982)) ?
                      reg2200[(5'h14):(5'h10)] : ((reg1353 >>> (7'h55)) <= (+(8'hbc))))});
              reg2214 = reg940;
              reg2215 <= {reg1349[(3'h4):(1'h0)]};
              reg2216 <= (^(+(&(~$unsigned((7'h48))))));
            end
          reg2217 <= ((~|((-forvar2212) ?
                  $unsigned(reg1052[(4'he):(4'h8)]) : ($signed(reg2207) > (reg1346 ?
                      reg963 : (8'h9e))))) ?
              ({$unsigned((reg1005 >> reg1353)), $unsigned(reg988), reg1362} ?
                  reg2205[(1'h0):(1'h0)] : ($signed({reg991}) && reg2210[(5'h13):(4'he)])) : (-(^reg986)));
          reg2218 = (reg1002 ?
              $unsigned(($unsigned(reg972) & $unsigned(reg944))) : $signed(((8'hb3) == ((&wire1772) ?
                  {wire927, (7'h56)} : (reg2211 != reg962)))));
          reg2219 = (|(~($unsigned((reg970 - reg1375)) ?
              reg1338 : $unsigned((^~reg2208)))));
          for (forvar2220 = (1'h0); (forvar2220 < (2'h3)); forvar2220 = (forvar2220 + (1'h1)))
            begin
              reg2221 <= reg970[(4'h9):(1'h0)];
              reg2222 <= reg997;
              reg2223 <= {(&(($signed(reg2216) >> $unsigned(forvar2197)) ?
                      (~^(reg1339 << (8'ha1))) : ($unsigned(reg1373) > $unsigned(reg1362)))),
                  ($signed($signed((reg2203 && wire924))) << (($signed(forvar2212) ^ $unsigned(reg996)) || ($signed(reg976) ?
                      {reg970, reg1025, reg933} : reg1372)))};
              reg2224 <= {{(~&(reg1369[(4'hb):(4'h9)] ?
                          $unsigned(wire928) : (forvar2206 & reg932))),
                      (($unsigned((8'had)) >> (~&reg2203)) >>> (reg1052 < $unsigned((8'h9f))))},
                  (^~((~|(reg1344 >= (8'hb9))) ?
                      $signed((|reg1052)) : ((~|reg1036) - $unsigned(wire1327))))};
            end
          reg2225 <= $signed((-$signed(reg957[(4'hd):(4'ha)])));
        end
      else
        begin
          if ((($signed(reg2222[(1'h0):(1'h0)]) <= ($signed(reg2209) ?
                  (7'h4c) : reg936)) ?
              reg982[(4'he):(3'h5)] : (~reg996[(4'h9):(2'h2)])))
            begin
              reg2212 = $unsigned((reg952 ?
                  reg1355[(3'h5):(3'h5)] : (~^reg990[(5'h12):(4'h8)])));
              reg2213 <= reg2208[(4'he):(3'h6)];
            end
          else
            begin
              reg2212 = (((~wire924) >> (((reg1355 >> wire1770) ?
                      $signed((8'h9e)) : reg2200[(3'h6):(2'h2)]) > {(reg941 ?
                          reg961 : reg1009),
                      (reg1345 ? (8'hb9) : (8'hb8))})) ?
                  wire927 : $unsigned(((~&(reg1357 > reg1374)) >= ((reg2210 ?
                      reg1355 : reg2215) * {reg1044}))));
            end
          for (forvar2214 = (1'h0); (forvar2214 < (2'h3)); forvar2214 = (forvar2214 + (1'h1)))
            begin
              reg2215 <= reg1043;
              reg2216 <= ((^((~^(|reg963)) <= (|$signed((7'h47))))) <<< $unsigned((($signed(reg2205) != $signed((7'h4e))) ?
                  (8'ha8) : $unsigned(reg1020[(5'h11):(4'hc)]))));
              reg2217 <= reg1343[(3'h5):(3'h4)];
            end
          reg2218 = ($signed(($unsigned((reg1370 ?
                  reg1374 : reg2204)) > (reg1020[(4'ha):(4'h9)] <= (reg1359 & reg1352)))) ?
              $unsigned({reg1375[(4'hd):(2'h3)],
                  $signed((wire1772 ? reg1001 : reg1036)),
                  ((wire928 ? reg1373 : reg944) ?
                      (reg933 * reg994) : (reg957 ?
                          reg966 : reg1057))}) : (^wire928));
        end
    end
  always
    @(posedge clk) begin
      reg2226 = (((reg932[(1'h1):(1'h1)] ? (~|(7'h47)) : $signed(reg2223)) ?
          ((8'hb3) ~^ ((reg976 >= reg1371) ?
              (~&reg996) : reg1335)) : {(~&$signed(reg1002)),
              (~&((8'hbf) >> reg962))}) >= (reg991 < reg932));
      reg2227 = ((~$unsigned(reg932)) & reg979[(3'h4):(2'h2)]);
      if (wire925)
        begin
          if (reg990)
            begin
              reg2228 <= (reg981 ?
                  (reg1362 ?
                      (|$unsigned(reg1001)) : reg1372) : reg1346[(4'he):(3'h5)]);
              reg2229 = reg1359[(4'h8):(4'h8)];
              reg2230 <= reg2216;
              reg2231 = {(((reg2227[(2'h3):(1'h0)] & (reg1353 ?
                              reg943 : (7'h53))) ?
                          ((reg979 || wire1770) ?
                              {reg2222,
                                  reg2223,
                                  reg1346} : $unsigned(reg1338)) : ({reg986} ?
                              reg1036[(4'h8):(3'h5)] : reg978[(4'he):(4'h9)])) ?
                      reg1010[(3'h6):(3'h6)] : $unsigned(reg955[(3'h5):(1'h1)]))};
            end
          else
            begin
              reg2228 <= {$signed((!reg1370[(5'h17):(3'h5)])),
                  (~|$signed((reg1353 ?
                      {wire926, reg982, reg1344} : {reg2222}))),
                  reg982[(4'hc):(4'h9)]};
              reg2230 <= $signed((7'h4d));
              reg2232 <= $unsigned({reg1347[(3'h7):(3'h6)],
                  {{(reg1352 ? (8'hae) : (8'hba))},
                      (&(!reg1338)),
                      $signed((reg1002 <<< reg1353))}});
            end
          reg2233 = (~|{reg979[(1'h1):(1'h0)],
              (-((+reg2215) >= (&reg1352))),
              (8'haf)});
          reg2234 <= (reg995[(2'h2):(2'h2)] ?
              $unsigned((reg1054 - reg1047)) : $unsigned({(reg936[(2'h3):(1'h1)] ?
                      ((7'h47) > reg1352) : {reg1345, reg2217, (8'hb3)})}));
          reg2235 <= reg2227;
          for (forvar2236 = (1'h0); (forvar2236 < (3'h6)); forvar2236 = (forvar2236 + (1'h1)))
            begin
              reg2237 = {$unsigned((~&{(~reg964)})),
                  $unsigned((reg1001[(5'h12):(5'h12)] == reg2235))};
              reg2238 = reg1020;
              reg2239 = (+(wire926 >> wire2195[(4'h8):(3'h5)]));
              reg2240 = ({$signed(reg1005),
                  reg956[(5'h13):(3'h5)]} << ((~|(|(~&reg944))) ~^ $signed(wire1770[(2'h3):(1'h1)])));
              reg2241 = (reg1339[(3'h7):(3'h4)] ?
                  $unsigned($signed($signed($signed(reg1044)))) : $signed(((~^(~&reg2228)) <<< $signed($signed(reg2222)))));
            end
          if ($unsigned(wire926[(1'h0):(1'h0)]))
            begin
              reg2242 <= (($signed($signed((reg940 & reg956))) ?
                  $signed(((~^(8'hbb)) ?
                      {reg1374,
                          reg941,
                          reg2239} : (8'hab))) : ($unsigned((^reg972)) ?
                      (^~reg1369) : reg1333)) - $unsigned(({reg933[(2'h3):(1'h0)],
                      $signed(reg2240),
                      (reg933 ? reg2222 : reg952)} ?
                  reg1050[(3'h6):(1'h0)] : reg1345[(2'h2):(1'h0)])));
              reg2243 = $signed({{(~|$signed((7'h49))),
                      reg2239,
                      $unsigned(((8'ha5) != reg1020))},
                  (8'hb6)});
              reg2244 = (({(((7'h54) || reg1345) - $signed(reg2228)),
                  {$unsigned(reg978),
                      (reg988 ? reg2203 : reg2203),
                      (reg1050 * reg1001)},
                  (reg1338 ?
                      (^~reg1009) : (reg1046 ?
                          reg1345 : (8'ha1)))} != (({reg1344, (8'hb5)} ?
                  $unsigned(reg952) : reg995[(1'h1):(1'h0)]) ^ $unsigned($unsigned(reg1373)))) ^~ $signed((reg1005[(1'h0):(1'h0)] ?
                  $signed({reg1352, reg2230}) : ((reg1345 ? (8'ha4) : reg966) ?
                      {reg2228, reg1373} : reg996))));
              reg2245 = (-$unsigned($signed(({reg1369,
                  (7'h55),
                  reg2202} != reg995[(1'h1):(1'h1)]))));
            end
          else
            begin
              reg2243 = (+$signed({(reg2229[(2'h2):(1'h0)] ?
                      (wire1772 == (7'h42)) : (|reg982)),
                  ($signed(reg2242) ? $unsigned((7'h4f)) : (reg972 > reg962)),
                  ((wire1013 ~^ reg2199) ?
                      $signed(reg1373) : reg2229[(2'h2):(1'h0)])}));
              reg2246 <= reg981;
              reg2247 <= (~|(((~$signed(reg1357)) > (!$signed((8'hbd)))) ?
                  (reg1025 ?
                      ((8'hb2) ?
                          (reg1333 + reg2238) : reg1023[(3'h5):(3'h5)]) : reg1349[(2'h3):(2'h2)]) : $unsigned(($unsigned((7'h53)) ?
                      $signed((8'ha0)) : $signed(reg1046)))));
              reg2248 <= (({reg1343[(1'h0):(1'h0)], (-(^~reg2242))} ?
                  $signed((7'h46)) : $signed((reg972 - (reg932 && reg981)))) | wire1772);
              reg2249 = (~&$unsigned((-{wire1013,
                  (!reg989),
                  ((8'hb1) ? (7'h4d) : reg1010)})));
            end
          if ($signed($signed(reg1036)))
            begin
              reg2250 = {(($unsigned((+reg2199)) ? (8'hb4) : $signed((8'ha0))) ?
                      ($signed((^~(7'h4b))) ^~ $signed((reg2246 <= reg2237))) : (+$unsigned((^~reg2243)))),
                  $unsigned($unsigned((reg2235 ^ (^~(8'hbe))))),
                  $unsigned((((reg2246 * reg1046) ?
                      ((7'h4e) ?
                          reg2240 : reg1054) : $signed(reg945)) == {reg1359[(1'h1):(1'h0)],
                      $signed(reg1020)}))};
              reg2251 = reg1036[(4'h9):(2'h2)];
              reg2252 = (~|((^~$unsigned(reg1345[(2'h2):(1'h1)])) && (((|reg2199) ?
                  $unsigned(reg2213) : (reg1353 ?
                      (8'hb3) : reg963)) || $signed($signed((8'h9f))))));
              reg2253 = $signed($signed($unsigned(reg1044)));
              reg2254 = reg2251[(4'ha):(3'h7)];
              reg2255 <= (reg2202 ?
                  reg961[(4'ha):(4'h9)] : $signed({$unsigned((8'ha0))}));
            end
          else
            begin
              reg2255 <= ((~{reg1043, reg2237}) ?
                  $signed({(reg2250 < reg943),
                      {(reg990 ? reg957 : reg2230),
                          {reg933, reg957},
                          {reg1010}},
                      reg2216}) : (^($unsigned((wire928 ? reg944 : (7'h56))) ?
                      {$unsigned(reg1333),
                          (reg1050 ?
                              reg994 : (8'hb9))} : ($unsigned(reg2234) ^ (+reg2227)))));
            end
        end
      else
        begin
          if ($signed(reg2233[(5'h17):(4'hc)]))
            begin
              reg2229 = wire2195[(3'h5):(1'h1)];
              reg2230 <= reg1339;
              reg2231 = $unsigned($signed((~^(reg1365 | (~reg2248)))));
              reg2232 <= ({reg988[(1'h1):(1'h0)],
                      $unsigned($signed($signed((7'h58)))),
                      wire1772[(5'h14):(3'h7)]} ?
                  reg1362 : ((+reg1345[(5'h11):(3'h6)]) ?
                      (+{{reg1020, reg2255, reg2202},
                          reg931,
                          reg985}) : reg2250[(5'h12):(3'h6)]));
              reg2234 <= ({(7'h42),
                  {{$signed(wire928), (reg961 ? reg1373 : reg943)}},
                  ((7'h4a) ?
                      ($signed(reg1369) & (~wire924)) : (reg988 & reg1343[(3'h4):(3'h4)]))} ^~ {($signed((reg966 ?
                          reg2253 : (8'hbe))) ?
                      {(!reg1372)} : $signed($unsigned(reg2216))),
                  reg990});
              reg2236 = (({(reg2237[(5'h10):(4'hf)] ?
                              $unsigned(reg986) : (^~reg1339)),
                          reg1369[(3'h7):(2'h2)]} ?
                      $unsigned(((reg1333 > reg932) ?
                          (reg2243 - reg1373) : $unsigned((7'h55)))) : {reg997}) ?
                  reg2216 : reg2213);
            end
          else
            begin
              reg2229 = ((^~{reg976,
                  reg957,
                  ($unsigned(reg1362) ?
                      (reg2242 ? reg1044 : reg955) : {reg1346,
                          reg2249,
                          reg2254})}) ^ ({(reg2216[(3'h5):(2'h2)] ?
                          ((8'hb2) ^ (8'hb3)) : (&reg1044))} ?
                  {(reg2250[(4'he):(4'h8)] ?
                          $signed(reg1362) : ((8'had) ?
                              reg2233 : reg2239))} : $unsigned({$unsigned(reg2253)})));
              reg2231 = ($signed($signed($unsigned((~^(7'h4a))))) >> reg1370);
              reg2233 = $unsigned(((((!(7'h4a)) != (wire925 ?
                      reg2225 : reg970)) ~^ $signed((reg2246 ?
                      reg1343 : (8'ha2)))) ?
                  reg2248 : ($signed($unsigned(reg1351)) ?
                      $signed((8'haf)) : (!reg936[(5'h1c):(4'h9)]))));
              reg2236 = (($unsigned((7'h4a)) ?
                  {reg2235[(4'hb):(4'h8)]} : {$signed((~|reg1372)),
                      ($unsigned(reg1344) ?
                          $signed(reg1023) : (reg1020 <<< reg957))}) == ($signed(reg2255) & reg1050[(4'hf):(4'h8)]));
              reg2237 = (~reg2235);
              reg2242 <= reg2250[(5'h14):(5'h11)];
            end
          reg2246 <= $unsigned($signed($signed({wire928})));
          reg2249 = (+($signed({reg2221[(3'h5):(2'h3)]}) < reg970));
          if ((~^$signed({(^$unsigned(reg2203))})))
            begin
              reg2250 = $signed({$unsigned(((^reg995) || (wire926 ?
                      reg932 : reg1353)))});
            end
          else
            begin
              reg2250 = reg1009;
              reg2255 <= (-reg962);
              reg2256 = (reg1043 - $unsigned(($unsigned(reg1020) != ($signed(reg2247) ?
                  {reg2237} : reg1373[(4'hd):(3'h7)]))));
              reg2257 = reg1338;
              reg2258 = $unsigned((~|reg976[(5'h11):(4'ha)]));
            end
        end
      reg2259 = (~(+{$unsigned((reg931 ? reg972 : reg1002)),
          ($unsigned(reg933) ? $signed(reg933) : (reg2199 && (8'h9e)))}));
    end
  assign wire2260 = reg976;
  always
    @(posedge clk) begin
      reg2261 = $signed($signed($signed((~|reg1353[(2'h2):(1'h1)]))));
      for (forvar2262 = (1'h0); (forvar2262 < (2'h3)); forvar2262 = (forvar2262 + (1'h1)))
        begin
          reg2263 <= (+(&wire926));
          reg2264 <= {(reg2230 ?
                  $unsigned({((8'hbf) ? wire926 : reg2232),
                      (reg2223 ? reg2213 : reg2235)}) : $unsigned(reg972)),
              (+(((8'ha5) ?
                  $signed(reg976) : ((7'h52) ?
                      reg2246 : reg2225)) ^ $unsigned({reg988})))};
        end
      if ($unsigned({($unsigned(((8'had) ?
              reg961 : (8'hbb))) <<< $unsigned((wire926 + reg1345))),
          reg1339}))
        begin
          for (forvar2265 = (1'h0); (forvar2265 < (3'h4)); forvar2265 = (forvar2265 + (1'h1)))
            begin
              reg2266 <= (&reg2230[(2'h2):(1'h0)]);
              reg2267 <= $unsigned(($signed(reg2248) >> (reg1002 ?
                  $unsigned(reg2247) : $signed({reg1044, reg957, reg966}))));
              reg2268 <= $signed(((reg1047[(5'h16):(3'h4)] ?
                  reg1352[(3'h5):(3'h4)] : reg1373[(4'he):(4'hb)]) * ((+(reg1036 ?
                  (7'h58) : reg2202)) - $unsigned((reg988 & reg990)))));
              reg2269 <= (+reg933);
              reg2270 <= (^reg931);
              reg2271 <= $signed(((((reg982 ?
                          reg2215 : (8'hbf)) <<< $unsigned(reg997)) ?
                      $unsigned((reg2266 ?
                          reg997 : reg2217)) : ({reg945} ^ $signed(reg964))) ?
                  reg1375[(3'h5):(3'h5)] : $signed($signed((forvar2262 ?
                      reg943 : reg2261)))));
            end
          reg2272 = reg2235[(2'h3):(2'h2)];
          if (wire2195[(3'h6):(1'h1)])
            begin
              reg2273 <= ((reg2266[(5'h14):(4'ha)] ?
                      wire2260[(3'h4):(2'h2)] : reg1362) ?
                  ($unsigned(((&reg1054) ?
                      reg978 : (reg2247 ?
                          reg2272 : reg2202))) >>> (reg2232 >>> reg1374)) : ($unsigned((reg1010[(4'h8):(3'h7)] ?
                      (forvar2262 <= wire1327) : $unsigned(reg1352))) >= $unsigned(reg1365)));
              reg2274 <= reg2266;
              reg2275 = (((({reg1044} ? (reg957 ? (7'h45) : reg944) : reg1374) ?
                      (~&$unsigned(reg1010)) : (8'hae)) ?
                  {wire926[(1'h0):(1'h0)],
                      $signed(forvar2265),
                      $signed(forvar2265[(1'h0):(1'h0)])} : $unsigned(reg1044)) << $signed($unsigned((-$unsigned((7'h47))))));
              reg2276 <= ({(reg1371 ?
                      $unsigned(reg2232) : reg2270[(5'h17):(4'hd)]),
                  reg1343[(3'h4):(1'h0)],
                  {reg2267}} ^~ $signed($unsigned(reg1345[(2'h2):(2'h2)])));
              reg2277 = $signed(((((reg2247 << reg936) ?
                          (^reg940) : $unsigned(wire927)) ?
                      reg940 : ($unsigned(reg1001) >= {reg1047, reg1335})) ?
                  reg2235[(4'hf):(4'hb)] : (!((~&wire924) >= reg941[(5'h16):(1'h0)]))));
            end
          else
            begin
              reg2275 = $signed((^reg2269[(1'h1):(1'h1)]));
              reg2277 = (({$unsigned($signed(reg1047))} ?
                      reg2202 : reg2225[(1'h0):(1'h0)]) ?
                  (($signed({reg979, reg994}) >>> ((|reg931) ?
                      reg2202 : (reg982 < reg1050))) ^ $signed($unsigned(reg2224))) : (reg976 ?
                      $unsigned($unsigned((reg962 ?
                          reg1054 : reg985))) : (^~reg1339)));
              reg2278 = $signed({{reg933[(1'h0):(1'h0)], (7'h4f)},
                  $unsigned($signed(wire924))});
              reg2279 <= (&(+{reg2268,
                  {(reg2266 ? (8'ha3) : reg1374),
                      (forvar2265 <= wire928),
                      reg1371[(4'ha):(4'ha)]},
                  reg2247}));
            end
          reg2280 = reg1335;
          if (($unsigned(((!$signed((7'h44))) ?
                  ($signed(wire2195) ^ {reg961}) : ((reg2235 << reg1343) ?
                      (&reg989) : (7'h49)))) ?
              reg985[(5'h1b):(4'hc)] : ($signed((~^reg2223[(5'h17):(2'h3)])) ?
                  (~^$unsigned((~|reg1044))) : $signed($signed(reg1338[(4'ha):(3'h6)])))))
            begin
              reg2281 <= {reg997[(5'h17):(2'h2)],
                  reg1054[(3'h4):(2'h3)],
                  (~{({reg1005} == $unsigned((8'ha1)))})};
              reg2282 <= $signed($signed(((((8'hb9) ? reg959 : reg1020) ?
                  wire928[(5'h18):(5'h18)] : (reg1343 && (7'h4d))) >>> $unsigned(reg2202))));
              reg2283 <= wire1327[(5'h13):(1'h1)];
              reg2284 = ($unsigned(((&(~|reg1047)) ? reg932 : reg1359)) ?
                  ($unsigned($unsigned(reg2235[(3'h7):(3'h7)])) + (!{{reg978,
                          reg1050,
                          wire924},
                      $unsigned(reg2221)})) : reg959);
              reg2285 <= reg1046;
              reg2286 <= reg933[(2'h3):(1'h1)];
              reg2287 <= $signed((~&($unsigned(reg2232[(5'h17):(1'h1)]) ?
                  reg2228 : $signed($unsigned(reg1372)))));
            end
          else
            begin
              reg2281 <= $signed((reg1370 ?
                  {($signed(reg2223) > (^~reg1005)),
                      ($unsigned(wire925) >= $unsigned(reg2270)),
                      reg979[(2'h2):(1'h1)]} : {$signed((reg931 ?
                          reg2270 : reg1370))}));
              reg2284 = (7'h4d);
              reg2285 <= (+reg1002);
              reg2288 = wire2260;
              reg2289 = ($unsigned((($unsigned(reg944) ?
                      $signed(reg972) : reg1372[(4'ha):(4'ha)]) + reg963)) ?
                  (8'hbe) : $unsigned($unsigned(((~reg2223) ?
                      (~^reg959) : $signed((7'h58))))));
              reg2290 <= $unsigned($signed(reg1375));
              reg2291 <= (7'h42);
            end
          if ($unsigned(($unsigned((~&(~^(7'h4d)))) | reg2217)))
            begin
              reg2292 <= $unsigned(reg1009);
              reg2293 <= reg1344;
            end
          else
            begin
              reg2294 = {$signed($signed((reg2199 << $unsigned(reg943)))),
                  (($signed(reg1335[(4'he):(2'h2)]) || ((reg981 ?
                      reg2199 : (7'h57)) <= reg2209)) >> reg1020[(4'he):(2'h2)]),
                  $unsigned($unsigned(({reg981,
                      reg1020,
                      reg2291} < (~^(8'ha8)))))};
              reg2295 = $signed($unsigned((reg2255 ?
                  (reg2213 == $unsigned(reg1333)) : forvar2265)));
              reg2296 <= reg955;
              reg2297 <= ({({((7'h4e) ^ reg2292),
                      (8'ha1)} >= wire2260)} >= $unsigned($unsigned($signed((+reg976)))));
              reg2298 <= ({({$signed(reg1023),
                      reg2248[(3'h7):(3'h6)],
                      reg1347[(3'h7):(1'h1)]} << ($signed(reg2269) ?
                      reg957[(4'hd):(3'h5)] : (reg1020 ~^ (7'h4c)))),
                  ($unsigned(wire2195) * (&(reg1369 & wire925)))} || (^~(-reg2266)));
            end
          for (forvar2299 = (1'h0); (forvar2299 < (3'h5)); forvar2299 = (forvar2299 + (1'h1)))
            begin
              reg2300 = $unsigned({$unsigned(reg1054[(3'h4):(1'h0)]),
                  (!($unsigned(reg2266) * ((8'h9c) ^ (7'h4e))))});
              reg2301 <= forvar2265;
              reg2302 <= (((+reg1355[(5'h11):(4'he)]) ?
                  (reg2203[(2'h3):(1'h1)] ?
                      (8'hbc) : (&$signed(reg2273))) : $signed(((&(8'hbb)) ?
                      reg2203 : (~^(7'h47))))) ^ $unsigned(reg2286));
              reg2303 = $unsigned($unsigned($unsigned(($signed(reg936) >= $unsigned(reg2248)))));
              reg2304 <= (~&reg982[(5'h10):(2'h2)]);
            end
        end
      else
        begin
          reg2265 <= (|$signed(reg2275[(2'h2):(2'h2)]));
          for (forvar2266 = (1'h0); (forvar2266 < (3'h6)); forvar2266 = (forvar2266 + (1'h1)))
            begin
              reg2267 <= $signed((8'hb5));
              reg2272 = $signed(reg1036);
              reg2273 <= forvar2265[(1'h0):(1'h0)];
              reg2274 <= reg1372;
            end
          for (forvar2275 = (1'h0); (forvar2275 < (2'h2)); forvar2275 = (forvar2275 + (1'h1)))
            begin
              reg2276 <= $signed($signed(reg2264));
              reg2279 <= {{reg2228[(1'h0):(1'h0)],
                      reg2273,
                      reg932[(1'h1):(1'h1)]}};
              reg2281 <= reg2246[(3'h6):(1'h1)];
              reg2282 <= $signed($signed($signed(((reg1009 >> reg1057) ?
                  (+reg1351) : $signed(reg2246)))));
              reg2284 = {(reg1345[(4'hc):(2'h3)] > (((reg1046 ?
                          (8'ha8) : reg1373) <<< (reg2289 ^~ reg2209)) ?
                      $signed(reg996[(4'hd):(3'h4)]) : $signed($signed(reg931)))),
                  (8'haa)};
              reg2288 = (reg1359 ?
                  $unsigned(reg2270[(4'hf):(1'h1)]) : wire928[(4'he):(4'hd)]);
            end
          reg2290 <= ({$unsigned($unsigned((reg955 ? reg996 : (8'hba)))),
                  ((~^$unsigned(reg1375)) << $unsigned((reg1346 ?
                      (7'h42) : reg2242))),
                  (8'hb4)} ?
              reg2225[(4'h8):(3'h6)] : reg981[(2'h3):(1'h0)]);
          if (((^~(~^$unsigned(reg994))) ?
              reg2246[(4'hb):(3'h7)] : reg2301[(5'h16):(2'h3)]))
            begin
              reg2294 = ($signed(wire2260[(3'h7):(3'h7)]) ?
                  ((reg1370 ? reg1353 : (^~$unsigned(reg1346))) ?
                      ((~|$signed(reg996)) ~^ ((reg2292 >= reg2268) <<< (wire1013 ?
                          reg2215 : (8'ha1)))) : $unsigned(reg989[(4'h9):(1'h1)])) : $unsigned(reg2215));
              reg2295 = ((reg1005 & (reg970 ?
                  reg2302[(4'hb):(3'h4)] : ($unsigned(wire2260) >>> forvar2266))) && $signed((^~(reg2266[(3'h4):(2'h2)] ?
                  (reg978 ? reg931 : wire1770) : reg2272))));
              reg2299 = reg1020[(3'h5):(2'h2)];
              reg2300 = ({$signed($unsigned(((8'had) + reg1054)))} && $unsigned(reg1373[(4'hb):(4'h8)]));
              reg2303 = reg1346[(3'h7):(3'h6)];
            end
          else
            begin
              reg2294 = $unsigned((($signed($signed(reg955)) ?
                  reg976 : $signed((reg986 && reg997))) != reg2234[(1'h1):(1'h1)]));
              reg2296 <= $unsigned(reg1346[(2'h3):(1'h0)]);
              reg2297 <= reg989;
              reg2298 <= ($signed(reg1365[(4'ha):(1'h0)]) ?
                  ((($unsigned(reg2255) ?
                      $signed(reg2222) : (reg2271 ?
                          reg1052 : reg2294)) || (~^(reg970 ?
                      reg2286 : reg2216))) <= (forvar2299 ?
                      $unsigned((^~reg2273)) : (!{reg2296,
                          reg1351,
                          reg2293}))) : ((-reg1339) ?
                      $signed($unsigned(reg2234[(1'h0):(1'h0)])) : {$unsigned(reg1009)}));
              reg2301 <= reg1346[(2'h2):(1'h0)];
            end
          if (($signed(reg1338) ?
              (reg2301[(5'h10):(4'h9)] > wire928) : {{$signed(reg2272[(2'h3):(2'h3)])},
                  (!reg2223)}))
            begin
              reg2305 = ({((reg2290[(3'h6):(1'h0)] < $unsigned(reg1044)) * $signed($signed(reg1352))),
                      (reg1050 ? reg1371 : reg961[(2'h3):(2'h3)]),
                      ($unsigned($signed((7'h48))) & ($signed(reg1374) * $unsigned(reg2224)))} ?
                  reg2294[(4'he):(3'h5)] : reg959[(5'h19):(4'h9)]);
            end
          else
            begin
              reg2304 <= $signed(($unsigned((^reg985)) * reg2255));
              reg2306 <= $unsigned($signed((~|(~|(wire926 ^ (7'h57))))));
              reg2307 <= ($unsigned(reg2304[(5'h17):(3'h4)]) <<< $signed($unsigned({$signed(reg2276),
                  (reg2290 && reg2280),
                  (reg1052 ? reg2274 : reg2234)})));
              reg2308 = reg2292;
              reg2309 <= $unsigned(reg2263);
              reg2310 = $unsigned(reg2225[(5'h1b):(4'h9)]);
            end
        end
      if ($signed(wire1013))
        begin
          if (({(reg1046[(3'h4):(1'h1)] ?
                  ($unsigned(reg1355) ?
                      $signed(reg1375) : reg982) : $signed($signed((8'h9e))))} > $unsigned(reg2209[(4'hd):(3'h4)])))
            begin
              reg2311 = (|{(7'h4f),
                  $signed($signed((reg2290 ? reg1353 : reg2291)))});
              reg2312 <= {$unsigned({(+(reg1005 >>> wire1013))}),
                  reg995,
                  reg1335[(4'hf):(4'hf)]};
              reg2313 <= $unsigned((^~(reg2216 ?
                  reg945[(1'h1):(1'h1)] : $unsigned(reg1002[(2'h3):(1'h0)]))));
              reg2314 = reg2225;
              reg2315 <= reg1001[(5'h15):(5'h15)];
              reg2316 <= (~^(8'hb0));
            end
          else
            begin
              reg2311 = (reg2263 | (reg2282[(5'h1e):(5'h13)] ?
                  reg2278[(4'hc):(3'h5)] : $signed($signed((|reg1343)))));
              reg2314 = $unsigned(($unsigned({reg940[(4'h9):(3'h6)]}) ?
                  reg1362 : wire928));
              reg2315 <= ($unsigned((($unsigned(reg2232) ?
                      forvar2299 : (~(8'hba))) ?
                  (~|reg2215) : (7'h4c))) | (^(+(&(!reg1054)))));
            end
        end
      else
        begin
          if (reg2268)
            begin
              reg2311 = $signed(($unsigned((&(8'hba))) ?
                  wire1770 : (($unsigned(reg931) ?
                      reg1052 : $signed(reg985)) | (~|(~&reg2297)))));
            end
          else
            begin
              reg2311 = $unsigned($signed(reg2298[(4'ha):(1'h0)]));
              reg2312 <= reg2307;
              reg2314 = reg2299;
            end
          reg2317 = $signed($unsigned(reg1001));
        end
      if (reg2296)
        begin
          reg2318 = reg1050[(4'ha):(4'h9)];
        end
      else
        begin
          reg2318 = $unsigned(reg991);
          if ($unsigned($signed($unsigned($signed((reg2311 ?
              reg1349 : reg2270))))))
            begin
              reg2319 <= ($signed(($signed((!reg2283)) ?
                      ((reg2203 ?
                          reg1001 : reg1335) ^ (reg985 * reg2308)) : reg1352)) ?
                  ({(+$unsigned(reg996)),
                          ((~&reg1355) ?
                              $signed(reg2301) : $unsigned(forvar2266)),
                          (!reg1346[(2'h2):(2'h2)])} ?
                      reg2230 : reg1009) : (!$unsigned(reg997[(2'h3):(2'h2)])));
              reg2320 <= reg2221[(4'he):(4'hb)];
              reg2321 <= reg2277[(5'h16):(3'h5)];
              reg2322 = ((~reg2199) ?
                  $unsigned(($unsigned($unsigned(reg2261)) ?
                      $unsigned((reg966 > reg2316)) : reg995[(3'h5):(1'h0)])) : $signed((~|(&wire2195[(3'h5):(3'h5)]))));
              reg2323 <= {($unsigned($unsigned($unsigned(reg995))) << $unsigned(((reg1009 ?
                      reg976 : forvar2266) <<< (reg1374 ? reg2312 : reg2247)))),
                  $unsigned(reg944[(2'h2):(1'h1)])};
              reg2324 = (+$unsigned(reg2310[(3'h4):(3'h4)]));
            end
          else
            begin
              reg2319 <= ((-({((8'hb5) ? wire1772 : reg1355),
                  (~&wire1772)} < ((reg1036 ? reg1052 : reg2234) ?
                  $unsigned(reg2221) : reg989[(4'h9):(4'h9)]))) == reg1009[(1'h1):(1'h1)]);
              reg2322 = $signed($signed(reg2305[(2'h3):(1'h1)]));
              reg2324 = reg2269[(1'h1):(1'h0)];
              reg2325 = ((reg970 ?
                  reg982[(4'hd):(2'h3)] : (~&{(reg931 ?
                          reg2303 : reg1338)})) <= $signed((^~$signed($unsigned(reg2313)))));
              reg2326 = reg972;
              reg2327 <= reg2294;
            end
          reg2328 <= (~(reg2295[(1'h1):(1'h1)] ?
              $signed({(reg2268 ? reg2294 : reg945)}) : (|reg2292)));
          if (reg2324[(5'h12):(4'hf)])
            begin
              reg2329 <= reg2283[(4'hf):(4'hd)];
              reg2330 = $unsigned($unsigned((-({reg986} ?
                  (!(8'hb3)) : reg1347[(4'hd):(1'h0)]))));
              reg2331 <= ({(($signed(wire924) <= $signed(reg1005)) ^ (reg2203 ?
                          $signed(reg962) : (~|(8'hbc))))} ?
                  reg1344[(5'h16):(3'h7)] : $signed($unsigned((~&$signed(reg1370)))));
              reg2332 = ((+reg1001) >> ($unsigned(reg991[(1'h1):(1'h1)]) ?
                  (7'h4d) : $signed((~(reg2328 ? (8'hb7) : reg1023)))));
              reg2333 = (wire2260[(2'h3):(2'h2)] == (&(!reg985[(5'h12):(2'h3)])));
            end
          else
            begin
              reg2330 = (({$unsigned($unsigned(reg2223)),
                      reg2321} & {$unsigned($unsigned(reg2292))}) ?
                  reg1365 : $unsigned(reg2286));
              reg2331 <= (8'ha8);
              reg2332 = {reg2255,
                  (($signed(((7'h50) - wire2260)) >> ((|reg2305) | $signed(reg2255))) * ((8'haa) ?
                      reg2317[(4'h9):(4'h8)] : ($signed((7'h42)) ?
                          (forvar2265 ^~ reg2310) : (reg981 > reg2286)))),
                  (reg2281[(5'h19):(4'hb)] < ($signed((^~reg2306)) ?
                      ((reg2216 >>> reg2322) ?
                          {(7'h51),
                              reg1369} : $unsigned(reg2263)) : $signed((reg2261 ?
                          (7'h48) : (8'hba)))))};
              reg2333 = ((reg981[(3'h4):(1'h1)] & reg1371) & $signed(reg997[(4'hf):(3'h4)]));
              reg2334 = $signed(((-($signed(reg2271) ?
                      $unsigned(reg2300) : $unsigned((7'h50)))) ?
                  (8'hba) : (~|$signed($signed(reg2292)))));
              reg2335 = $signed((~^(~&{$signed(reg2234),
                  reg936[(4'hd):(4'hc)]})));
              reg2336 <= (&(~{reg970[(4'h8):(2'h3)], reg1046}));
            end
        end
    end
  assign wire2337 = {{((reg1043[(2'h3):(2'h3)] & reg1339) ?
                                $signed($unsigned(reg1374)) : (reg1372 ?
                                    reg2216[(5'h18):(4'h8)] : (reg1351 ?
                                        reg1369 : reg985))),
                            $unsigned((reg1345 ?
                                (reg976 ?
                                    reg1025 : reg941) : $signed((8'hbf)))),
                            $signed(($signed(reg2279) << $signed(reg1335)))}};
  assign wire2338 = $unsigned($signed((~^{$unsigned(reg2290), (-reg2287)})));
  assign wire2339 = reg2302;
  always
    @(posedge clk) begin
      reg2340 <= (~&{(~^$unsigned((-reg2304))),
          (reg2234[(4'h9):(1'h0)] ? $signed(reg2203) : {$signed(wire924)}),
          reg2309});
    end
  always
    @(posedge clk) begin
      if (reg2320[(4'hd):(3'h5)])
        begin
          for (forvar2341 = (1'h0); (forvar2341 < (3'h4)); forvar2341 = (forvar2341 + (1'h1)))
            begin
              reg2342 <= reg2327[(1'h0):(1'h0)];
              reg2343 = {reg994[(4'ha):(1'h1)],
                  ($unsigned((~(+reg1050))) ?
                      ((~^reg2313) ?
                          $unsigned(reg1346[(1'h0):(1'h0)]) : wire928[(5'h11):(4'hc)]) : reg1338[(4'h8):(3'h5)]),
                  (~^reg2296)};
              reg2344 <= $unsigned($signed((~^$unsigned((~|(7'h56))))));
              reg2345 <= reg2291;
              reg2346 = (reg2221[(5'h12):(4'hb)] ?
                  {$signed(((reg1347 + reg956) || (reg2286 ~^ reg1345))),
                      reg996[(4'hf):(4'h8)]} : ((reg1036 > (7'h4f)) ?
                      {((reg2286 ?
                              reg2221 : reg1353) ^~ $signed(reg997))} : (reg1057 == reg2281)));
              reg2347 <= $signed(({reg2270[(4'ha):(4'ha)],
                      (~$signed(reg2321)),
                      $signed(reg2343[(5'h10):(3'h4)])} ?
                  $signed(reg2290) : $unsigned({reg2342[(3'h4):(2'h2)],
                      (^reg957),
                      (^reg2270)})));
              reg2348 = reg2282;
            end
          if (reg1001[(5'h17):(3'h4)])
            begin
              reg2349 <= reg2292[(4'hb):(4'h9)];
              reg2350 = $signed(($unsigned((reg2344[(5'h19):(5'h11)] ?
                  $signed(reg959) : (reg932 <= reg2306))) > ({{(7'h56),
                      wire2338},
                  (reg2346 ^~ wire925),
                  (reg2285 ? reg1333 : (8'haf))} != (7'h54))));
              reg2351 <= $signed(reg963);
              reg2352 = (~&reg1036[(4'h9):(1'h0)]);
              reg2353 <= $unsigned({$signed(reg2265)});
            end
          else
            begin
              reg2349 <= reg2216;
              reg2350 = {reg2319[(2'h2):(1'h0)], $unsigned(reg1057)};
              reg2352 = reg2264[(2'h3):(1'h1)];
              reg2353 <= $signed($signed(((~^(~^reg2246)) ^ (reg941 - wire927))));
              reg2354 = wire928;
            end
        end
      else
        begin
          reg2341 <= {(({$unsigned(reg1046), reg2296} ?
                      (8'ha3) : ((+reg1349) ?
                          {reg2285, reg995} : (reg1050 > reg1372))) ?
                  {$unsigned((reg931 > reg2352))} : $unsigned({{reg2199},
                      (~^reg2213)})),
              reg2343[(1'h1):(1'h0)]};
        end
      reg2355 = (~^reg2350);
      if ($unsigned(reg2247[(3'h5):(1'h1)]))
        begin
          reg2356 <= ((reg2265 >= (8'h9c)) ?
              $signed($unsigned(reg940)) : (!{reg2266}));
          if ((~($signed($signed((reg1347 ?
              reg2232 : wire927))) * {{$signed(reg2279),
                  (reg2336 ? reg2217 : (7'h47))}})))
            begin
              reg2357 <= reg991;
              reg2358 <= reg1346[(4'h8):(3'h7)];
              reg2359 <= $signed($signed(wire2337));
              reg2360 <= $unsigned((~|reg940[(4'he):(2'h3)]));
              reg2361 = (reg2346 ?
                  {$signed(((reg2286 != reg995) * (reg1371 >> (7'h55))))} : (&$signed($unsigned((reg1373 - forvar2341)))));
            end
          else
            begin
              reg2357 <= $signed(($signed(reg1052) > wire2339[(2'h2):(1'h1)]));
              reg2361 = ($unsigned($signed($signed((reg2350 ?
                      (7'h58) : reg1054)))) ?
                  reg1355[(1'h0):(1'h0)] : ((wire928[(2'h3):(1'h1)] ?
                          ((reg988 ? reg1352 : reg964) ?
                              reg2323 : {reg1036}) : $unsigned((reg2209 ?
                              reg955 : reg2213))) ?
                      (((reg943 ? reg2230 : reg2336) <<< ((8'hbe) ?
                              reg2343 : (8'hb7))) ?
                          ($unsigned(reg1353) ?
                              ((7'h40) ~^ reg1036) : $signed(wire1013)) : reg1339[(4'ha):(3'h5)]) : (((^~reg979) <= reg1020[(3'h5):(1'h0)]) ?
                          $unsigned({(7'h49),
                              reg1054}) : $unsigned($unsigned(reg943)))));
              reg2362 <= ((|$signed({reg972,
                  $signed(reg2279)})) >= (~^reg2271[(4'h8):(2'h2)]));
              reg2363 <= $unsigned(reg1359);
            end
          for (forvar2364 = (1'h0); (forvar2364 < (1'h1)); forvar2364 = (forvar2364 + (1'h1)))
            begin
              reg2365 = (((7'h47) ?
                      reg976[(4'hc):(4'h9)] : {(~^$signed(reg978)),
                          $unsigned($signed(reg994))}) ?
                  $signed((reg956 ?
                      $unsigned((7'h56)) : ((~reg2316) & reg2273))) : (!$signed(reg955)));
            end
          for (forvar2366 = (1'h0); (forvar2366 < (2'h3)); forvar2366 = (forvar2366 + (1'h1)))
            begin
              reg2367 <= ($signed(reg981[(3'h4):(1'h0)]) ?
                  (({reg2271, (reg997 ? (8'hbb) : (8'hbb))} ?
                      $signed({reg2315,
                          reg1005}) : $signed(reg1351)) || ((reg2358 ?
                      $signed(reg2365) : $unsigned(reg2336)) || reg1345)) : (reg1357 + (({reg2270,
                          (7'h48)} ?
                      (&reg940) : $signed(reg1365)) <<< $unsigned({reg2360,
                      (8'h9e),
                      reg2350}))));
              reg2368 <= $unsigned($unsigned((^$unsigned($unsigned((8'ha1))))));
              reg2369 = $unsigned(((reg2279[(2'h3):(1'h0)] ?
                      $signed(((7'h46) ?
                          reg2263 : (7'h52))) : reg2356[(3'h4):(2'h3)]) ?
                  $unsigned((reg2255 < ((8'hb2) ?
                      reg2228 : reg956))) : reg964[(1'h0):(1'h0)]));
              reg2370 = reg2203[(2'h2):(1'h1)];
              reg2371 = ((7'h56) + forvar2366);
              reg2372 = ((~reg985) ^ (&$unsigned(((reg1001 ?
                  reg2263 : reg2371) && (~(8'had))))));
            end
          for (forvar2373 = (1'h0); (forvar2373 < (3'h4)); forvar2373 = (forvar2373 + (1'h1)))
            begin
              reg2374 = ((7'h43) <<< {$unsigned(((reg1372 ^~ reg943) ^~ (8'hba)))});
              reg2375 = ($unsigned(reg994[(1'h1):(1'h0)]) ?
                  reg1353 : $unsigned($signed($signed($signed(reg2235)))));
              reg2376 = {forvar2341[(5'h1b):(4'h8)]};
            end
          for (forvar2377 = (1'h0); (forvar2377 < (2'h3)); forvar2377 = (forvar2377 + (1'h1)))
            begin
              reg2378 <= reg2235[(4'ha):(4'h8)];
              reg2379 = $unsigned({$signed((8'had))});
              reg2380 <= (reg1362 ~^ $unsigned((reg2344 << reg2292)));
              reg2381 <= (-$signed((($unsigned((8'ha2)) ^~ ((8'haa) ?
                  reg2357 : reg2222)) << (reg1005 * (|reg1352)))));
              reg2382 <= (~^$signed((7'h40)));
              reg2383 <= ((|(8'haf)) << reg2222);
              reg2384 = (^~((reg2209 <<< ((-reg2304) | $unsigned(reg2342))) >> (8'hb1)));
            end
          if (((reg2344[(5'h11):(4'hb)] ?
              (~&reg2362[(3'h4):(2'h3)]) : (~reg991[(2'h2):(2'h2)])) >> $unsigned(($signed((reg2298 && reg2367)) ?
              reg1339[(2'h3):(2'h2)] : $unsigned($unsigned((8'hba)))))))
            begin
              reg2385 <= $unsigned((8'ha9));
            end
          else
            begin
              reg2386 = ((!(~&reg2319)) & ({{$signed(reg2313), reg1373},
                      reg970[(2'h2):(1'h1)]} ?
                  {$signed(reg2323[(1'h1):(1'h0)]),
                      (reg2312 << reg1346),
                      (!$signed(reg2362))} : $signed({$unsigned(reg972),
                      (reg2281 <= reg936),
                      (reg2290 ? reg961 : reg1344)})));
              reg2387 <= (|(~&reg2368[(1'h1):(1'h0)]));
              reg2388 <= ({(((reg1355 ^~ reg961) ?
                          $signed((7'h4b)) : reg2376) <= reg2247)} ?
                  ((+reg988[(1'h1):(1'h1)]) ?
                      reg2283 : {{reg2328,
                              $unsigned((7'h4c))}}) : $signed(reg1020));
              reg2389 <= wire926;
              reg2390 <= reg933[(1'h0):(1'h0)];
              reg2391 <= (reg2375 ?
                  (($signed({reg1023, (8'had)}) ?
                      reg997 : $signed(reg2388)) >>> reg1057) : $signed({(^~reg970),
                      {$signed(reg1010), $signed(reg2276), $signed(reg2343)}}));
            end
        end
      else
        begin
          reg2361 = ((+(((reg2376 ?
                      reg2276 : reg1044) < reg1338[(4'h8):(2'h3)]) ?
                  $signed($signed(forvar2364)) : ((reg2286 * reg2341) >>> (forvar2373 ?
                      (8'hab) : reg2222)))) ?
              reg1370 : $signed((^~($signed(reg2282) ?
                  (+reg2276) : (~&(7'h4e))))));
        end
      if (reg994[(4'h9):(4'h8)])
        begin
          for (forvar2392 = (1'h0); (forvar2392 < (3'h4)); forvar2392 = (forvar2392 + (1'h1)))
            begin
              reg2393 = (reg2342[(3'h4):(3'h4)] ?
                  ($signed(reg2283) & ($unsigned((|(8'hbe))) || wire1327)) : $signed(reg1352));
              reg2394 <= ($signed(({{reg1054, (7'h52), reg996},
                      $signed((8'hbb)),
                      $unsigned(forvar2392)} >> {$unsigned(reg2353),
                      (reg2313 ? reg2393 : (8'hbb)),
                      ((7'h4d) ? reg945 : (7'h43))})) ?
                  ({($signed(reg2327) <= reg932[(4'h9):(3'h4)]),
                          {(reg2390 ? reg1005 : reg2266),
                              $unsigned(reg2276),
                              reg2368}} ?
                      ({reg2327,
                          (reg1347 ?
                              reg2371 : reg2382)} - reg2381[(3'h5):(3'h4)]) : $unsigned({{reg2391,
                              reg940,
                              reg2381},
                          (reg2359 < (8'ha3))})) : (+wire2339));
              reg2395 = reg1355[(4'hd):(4'hc)];
              reg2396 <= $signed((^(|((reg2375 <= wire924) || ((7'h4a) | wire2339)))));
              reg2397 <= (reg2268[(1'h1):(1'h0)] ?
                  ($unsigned(reg2297[(4'hd):(4'h9)]) ?
                      ((reg966 ~^ reg2203[(2'h3):(2'h2)]) ?
                          reg2359[(1'h1):(1'h1)] : $signed($unsigned(reg1023))) : reg1025[(4'hf):(1'h1)]) : (reg1054 ?
                      reg2255 : $unsigned((~&wire928))));
              reg2398 <= $signed($signed(reg964[(1'h1):(1'h1)]));
            end
          for (forvar2399 = (1'h0); (forvar2399 < (1'h1)); forvar2399 = (forvar2399 + (1'h1)))
            begin
              reg2400 = reg2344;
            end
          reg2401 <= reg2384;
          for (forvar2402 = (1'h0); (forvar2402 < (3'h4)); forvar2402 = (forvar2402 + (1'h1)))
            begin
              reg2403 = (+reg2216[(4'he):(2'h2)]);
              reg2404 <= {(~^$signed($unsigned(reg941))),
                  forvar2399[(2'h2):(1'h0)],
                  (($signed({reg2286}) ^~ (+wire1013[(5'h15):(5'h10)])) ?
                      ({reg1357[(4'hc):(4'h9)],
                          {reg1044},
                          (^reg2372)} <= $signed((~|reg944))) : reg1023)};
              reg2405 <= (^$signed((8'haa)));
              reg2406 = ((^~(((~^reg2276) <= $signed((7'h43))) ?
                      $signed((wire926 > reg2323)) : (reg2321 << reg2217[(5'h14):(1'h0)]))) ?
                  ($unsigned((7'h44)) * ((((7'h42) ~^ reg1362) << reg2343) ?
                      (&$unsigned(reg964)) : ((~&reg2306) ?
                          $signed(reg1009) : $signed(reg2286)))) : reg2319[(2'h3):(1'h1)]);
            end
          reg2407 = $signed(((~^{(~^reg1365), $unsigned(reg982)}) * reg1338));
          for (forvar2408 = (1'h0); (forvar2408 < (1'h0)); forvar2408 = (forvar2408 + (1'h1)))
            begin
              reg2409 = (8'ha2);
              reg2410 = ($signed($signed(reg2393[(1'h0):(1'h0)])) ?
                  ((8'ha5) ? reg1043 : forvar2408) : reg2286);
              reg2411 <= ($unsigned({$signed($signed(reg2316))}) ?
                  reg1357[(3'h4):(2'h2)] : (+($signed({reg961, reg981}) ?
                      reg2359 : {((7'h43) < reg1352), (reg940 & reg988)})));
              reg2412 = reg2320[(3'h7):(1'h0)];
              reg2413 <= reg2266[(5'h10):(3'h6)];
            end
          reg2414 = (-reg2365);
        end
      else
        begin
          for (forvar2392 = (1'h0); (forvar2392 < (3'h4)); forvar2392 = (forvar2392 + (1'h1)))
            begin
              reg2394 <= (($signed((reg2246[(3'h7):(3'h5)] <<< $unsigned((7'h4c)))) <<< ((reg2232 == reg2279) != $signed($signed(reg2319)))) ?
                  ((reg1052 ^ ((reg2376 ? reg2371 : (8'h9e)) >>> {reg1344})) ?
                      (^((reg2359 ? wire924 : reg1371) ?
                          wire928 : (8'h9e))) : (~&(8'ha1))) : (+reg2356[(4'h9):(4'h8)]));
              reg2395 = reg944[(2'h2):(1'h0)];
              reg2396 <= reg933[(2'h2):(1'h1)];
              reg2399 = {(&({reg2378[(4'hc):(4'hb)]} ~^ ($unsigned(reg970) * (reg1349 - reg989)))),
                  ((reg955 | reg2336) <= $signed({reg2225[(5'h1a):(5'h15)],
                      $signed(reg2400),
                      (reg2301 ? reg964 : reg2389)}))};
            end
          for (forvar2400 = (1'h0); (forvar2400 < (2'h2)); forvar2400 = (forvar2400 + (1'h1)))
            begin
              reg2402 = (+(8'hab));
              reg2403 = $unsigned((7'h40));
              reg2406 = ((reg1043[(3'h4):(3'h4)] ^~ $unsigned($unsigned(reg940[(2'h3):(2'h3)]))) >= {$signed(reg936[(1'h1):(1'h0)]),
                  {$unsigned((|reg2248))},
                  $signed(($unsigned(reg1351) == $unsigned(reg2232)))});
              reg2407 = ($signed(reg1355[(5'h14):(1'h1)]) ?
                  $unsigned($signed($signed(reg2406[(2'h2):(1'h0)]))) : ({(8'haa)} ?
                      $signed(reg2281[(5'h10):(1'h1)]) : ((7'h45) ^ reg2302)));
              reg2408 = ($unsigned(($unsigned({reg2304}) ?
                      {$signed(reg2351),
                          {(8'hae), reg2293, reg956},
                          {reg2396}} : $signed(forvar2373[(4'hf):(2'h3)]))) ?
                  (|(+(reg1345 ?
                      (|reg1047) : $unsigned((8'hbb))))) : $unsigned((&(!reg970))));
              reg2409 = reg936;
              reg2411 <= ((~|(~^$signed((8'h9e)))) || {reg2248[(3'h6):(2'h3)],
                  $signed((reg982 ?
                      (reg2302 ? reg2349 : reg936) : (reg2360 | reg2390))),
                  reg2329[(2'h2):(2'h2)]});
            end
          if (((&($signed($signed((8'ha6))) >>> $signed((reg2390 ?
              reg1345 : reg970)))) <<< reg985[(5'h17):(3'h4)]))
            begin
              reg2412 = wire2339[(2'h2):(1'h1)];
              reg2414 = (-((^~(|reg2304)) == (|wire2339)));
              reg2415 <= ((($signed((~&reg966)) | (reg2307[(1'h0):(1'h0)] ?
                      (reg2202 ?
                          reg2202 : (7'h54)) : reg2360[(5'h16):(5'h12)])) ?
                  (!$signed($signed(reg2412))) : (reg1352[(3'h5):(3'h4)] ?
                      ($signed(reg2342) ?
                          {(7'h46), reg1339} : {reg2287,
                              reg2242,
                              reg988}) : ($signed((7'h45)) ^ ((8'hbc) >= reg943)))) >> {reg2372,
                  $unsigned((7'h46))});
              reg2416 = (|((((wire924 ? reg2359 : reg2271) ?
                      (^reg1043) : (reg2279 ? (8'ha8) : wire2260)) ?
                  (7'h47) : $unsigned($signed((7'h41)))) ^~ $unsigned(($unsigned(reg2225) ?
                  (7'h43) : reg2232))));
              reg2417 = ((8'ha5) >> reg2283);
              reg2418 <= (+(reg963[(3'h4):(1'h0)] << $unsigned($signed((~&reg2397)))));
            end
          else
            begin
              reg2413 <= reg2387[(1'h1):(1'h1)];
              reg2415 <= $signed($unsigned((reg2255[(2'h2):(1'h1)] ?
                  ((7'h46) ? reg961 : (reg952 ? (7'h52) : reg1359)) : reg959)));
              reg2416 = (~^reg2306[(5'h17):(1'h1)]);
              reg2417 = ((~($unsigned($signed(reg2293)) <<< $unsigned(((8'h9f) ?
                      reg2298 : reg2413)))) ?
                  $unsigned($unsigned((~$unsigned(wire926)))) : ((reg2209 ?
                      (((7'h54) ?
                          (8'hb7) : reg1338) << $unsigned(reg2341)) : (+(-wire928))) ^~ $signed(reg2307[(1'h0):(1'h0)])));
              reg2418 <= {{(8'ha1)},
                  (reg1375 >= reg2383[(4'he):(4'hc)]),
                  ($signed(reg1346) ?
                      (reg2213[(3'h4):(2'h2)] >>> reg2224) : $unsigned(reg957))};
            end
          reg2419 <= $unsigned(($signed(reg1052) ?
              (|$signed(reg2235)) : ((~|{(8'hbd), reg2216, reg2403}) ?
                  {{reg2352, forvar2366, reg1351},
                      (|reg2418),
                      (7'h54)} : (reg2418[(2'h2):(2'h2)] ?
                      $unsigned(reg1359) : reg2279[(3'h6):(2'h2)]))));
          for (forvar2420 = (1'h0); (forvar2420 < (3'h4)); forvar2420 = (forvar2420 + (1'h1)))
            begin
              reg2421 <= $unsigned(reg2395);
              reg2422 = $signed(reg2267);
              reg2423 <= (7'h52);
              reg2424 = reg2343;
              reg2425 <= $unsigned($signed(((forvar2366 ?
                  (-(8'hb0)) : (^~reg2419)) != (reg1362[(5'h1b):(5'h15)] < $unsigned(reg1370)))));
              reg2426 = (($unsigned(reg933) ?
                  reg2395 : (~&$unsigned((^(8'h9d))))) <<< ($unsigned((8'ha5)) ?
                  $unsigned(($signed(reg2228) ?
                      reg2355 : $unsigned((8'ha8)))) : forvar2366[(3'h4):(2'h3)]));
              reg2427 <= ($signed((forvar2364 + (((8'hbd) ?
                  reg2379 : reg981) <= wire927))) < $unsigned({reg2387,
                  reg1046[(1'h1):(1'h0)]}));
            end
          reg2428 <= reg2400[(2'h2):(1'h1)];
          reg2429 <= ((($signed($unsigned(reg2370)) - $unsigned($signed(reg2400))) == $unsigned($unsigned(reg2319[(1'h1):(1'h1)]))) >>> (wire2337[(1'h0):(1'h0)] << reg2343[(4'hd):(3'h7)]));
        end
      reg2430 <= ($signed((^$signed((^~reg2349)))) <= $unsigned((-reg963[(3'h7):(2'h3)])));
      if ($unsigned($signed(forvar2377[(1'h0):(1'h0)])))
        begin
          if ((reg1347[(3'h6):(3'h4)] != reg2397))
            begin
              reg2431 = reg2290[(3'h4):(1'h1)];
              reg2432 <= $signed((reg2323 >> $signed((7'h4e))));
              reg2433 <= {(reg2404 ?
                      $signed(reg2372) : ((~{reg2357}) ?
                          $signed({reg1347, reg2400, reg964}) : (8'hbe)))};
              reg2434 = $signed((7'h43));
              reg2435 <= $signed(reg2328);
            end
          else
            begin
              reg2431 = wire927[(5'h18):(4'hc)];
              reg2434 = reg961;
            end
          if ({($unsigned((reg1009[(4'h8):(3'h7)] * reg2389)) * ($signed((-reg1047)) <<< (-$unsigned(reg2354)))),
              reg2422[(4'hf):(4'he)],
              $signed((8'hbd))})
            begin
              reg2436 <= ((|(!((reg2394 ? reg2301 : wire2339) ?
                      reg1355 : {reg978, reg2235, forvar2408}))) ?
                  reg2268 : ((({reg2293, reg2312} && reg2414[(4'hf):(4'hc)]) ?
                      (-(reg1005 == reg957)) : (reg2320 ?
                          reg2386 : $unsigned(reg2217))) | reg994));
            end
          else
            begin
              reg2436 <= {reg2367};
              reg2437 = $unsigned(reg2230);
              reg2438 <= reg2405[(2'h3):(2'h2)];
              reg2439 <= reg995;
            end
          reg2440 <= ($signed((((reg962 ?
              reg2406 : wire1770) < {(8'hbb)}) ^ reg2312[(2'h2):(2'h2)])) ^ (reg2358[(3'h6):(3'h5)] ?
              $unsigned(reg1355[(3'h6):(1'h1)]) : $unsigned(reg2302)));
          reg2441 = {(^{$signed((8'hbc))})};
          reg2442 = $signed({$signed((^(wire2195 ? (7'h4c) : reg1005)))});
          if ({(~&(&reg2407[(5'h10):(2'h2)])),
              reg2216,
              ((8'ha9) | (reg2349[(1'h1):(1'h0)] ?
                  {$unsigned(reg2228),
                      {forvar2377,
                          reg2369,
                          reg955}} : (&reg2269[(1'h1):(1'h0)])))})
            begin
              reg2443 = (((|((+reg2255) ?
                  wire926[(4'h8):(2'h2)] : (^~(8'h9c)))) | (7'h4d)) - $signed((($unsigned(reg2390) ~^ (&reg1335)) + $signed((reg2224 != (8'hb9))))));
              reg2444 = (^($unsigned((reg1339 ?
                      forvar2377[(4'hb):(2'h3)] : $signed(reg2395))) ?
                  forvar2400[(5'h14):(4'h8)] : reg2412[(5'h1d):(4'hc)]));
              reg2445 = wire1770;
              reg2446 = (8'haf);
              reg2447 <= $signed(reg940);
              reg2448 <= $signed((8'ha4));
              reg2449 <= (|$unsigned(((reg2341 ?
                  (forvar2392 * (8'hbd)) : $unsigned((7'h43))) * $signed({reg1365,
                  reg1333,
                  reg2421}))));
            end
          else
            begin
              reg2443 = $unsigned((8'hb0));
              reg2444 = $unsigned($signed(reg2283[(3'h4):(1'h0)]));
              reg2447 <= $signed((!($unsigned((reg1343 ? reg1052 : reg2351)) ?
                  ((reg2381 ?
                      forvar2402 : reg2379) <= $unsigned(reg2418)) : ((reg2402 ?
                      reg2397 : reg1043) & (reg2348 ? (7'h52) : reg2215)))));
              reg2450 = (~&reg2447);
              reg2451 <= ($signed(((^~reg2328[(4'hb):(3'h7)]) <= (((7'h54) ?
                      reg2440 : reg2406) || (reg2367 ? reg1345 : reg2403)))) ?
                  reg2438[(5'h12):(3'h7)] : (reg2411[(4'h8):(3'h5)] | {(|(^reg2345)),
                      ((reg2393 ? reg2202 : reg1370) < reg2291),
                      ((reg2379 ? reg1346 : reg1057) ?
                          {reg2209,
                              reg2426,
                              reg2222} : reg2437[(2'h3):(1'h0)])}));
              reg2452 <= ((($signed((~reg931)) ~^ reg2383[(5'h10):(1'h1)]) <= $signed($signed(reg2388))) >>> {$signed(reg1362)});
              reg2453 <= $signed({reg2449,
                  {(((7'h41) ? reg1002 : reg2221) ?
                          (reg1369 ^ reg1046) : reg2435)},
                  (~|{wire928[(4'hd):(3'h4)]})});
            end
        end
      else
        begin
          reg2431 = reg932;
          reg2434 = ($unsigned(reg2437) ? (8'ha0) : $signed(reg988));
          if ((7'h49))
            begin
              reg2435 <= (&reg2450);
              reg2437 = (+$unsigned(reg995[(3'h4):(3'h4)]));
              reg2438 <= (-(reg2292[(4'hb):(3'h6)] >>> reg1339[(3'h5):(2'h2)]));
              reg2441 = $signed(((^{reg1005}) >> $unsigned(($unsigned(reg2355) << reg990[(4'hb):(3'h7)]))));
            end
          else
            begin
              reg2435 <= reg1023;
              reg2436 <= reg2202;
              reg2437 = $signed(reg2352[(1'h1):(1'h0)]);
              reg2441 = (reg2397[(5'h16):(2'h3)] <<< forvar2400[(4'he):(3'h6)]);
              reg2447 <= (!reg1020[(5'h11):(4'hd)]);
              reg2450 = (+reg933[(2'h3):(1'h0)]);
              reg2451 <= ($unsigned(reg2342) ?
                  $signed((reg970[(3'h7):(3'h6)] < reg2437)) : (((forvar2420[(4'hb):(3'h4)] <<< $signed(forvar2392)) ?
                      $unsigned($signed(reg2248)) : ((reg2279 << (7'h41)) >> $signed(reg2432))) & reg1359[(5'h13):(3'h7)]));
            end
          reg2454 = ($unsigned($unsigned((reg964[(2'h2):(1'h0)] ?
                  reg2419[(4'hf):(4'he)] : $unsigned(reg2399)))) ?
              (8'ha8) : (reg2409 ?
                  $unsigned((7'h50)) : (((^reg2276) ?
                          $signed((8'hb1)) : $signed(reg1052)) ?
                      (~^$signed(reg988)) : ((reg2307 ^~ reg2342) ?
                          {reg2342, reg952, (8'ha7)} : (forvar2408 ?
                              reg2388 : wire1013)))));
          reg2455 <= (reg1375[(3'h4):(1'h0)] > (-reg2271[(4'hd):(1'h0)]));
          if ($signed(reg1347[(3'h5):(1'h0)]))
            begin
              reg2456 <= $signed($signed((reg1359[(2'h3):(1'h1)] * $signed($signed(reg963)))));
              reg2457 <= (7'h45);
              reg2458 = $signed({reg1002[(4'h9):(3'h5)],
                  $signed(reg2306[(3'h7):(1'h1)])});
              reg2459 = ($unsigned({forvar2408,
                      $signed((reg952 >>> reg2389))}) ?
                  (~&{{((8'hb9) | reg2404), reg936}, reg963}) : (8'hb2));
            end
          else
            begin
              reg2458 = reg2451[(2'h3):(2'h3)];
              reg2460 <= reg2329[(3'h4):(2'h2)];
              reg2461 <= (^$unsigned((($unsigned(reg2355) != $unsigned(reg2228)) ?
                  {reg957[(4'h8):(3'h6)],
                      $signed(reg2230)} : reg1374[(4'he):(4'hb)])));
              reg2462 = $signed({reg1351[(4'he):(2'h2)],
                  ($signed((~|wire1770)) >= (((7'h58) ?
                      reg2438 : reg2428) >> reg2430[(4'h8):(3'h7)]))});
              reg2463 = forvar2373;
              reg2464 = $signed(reg2434[(2'h3):(1'h1)]);
              reg2465 = (^~reg2353[(3'h6):(2'h3)]);
            end
          reg2466 = $unsigned(((~($signed(reg2271) ~^ $signed(reg1362))) ?
              ($signed($signed(reg1044)) >>> ((~^reg989) ?
                  (7'h51) : (reg2403 && reg2234))) : $signed((7'h53))));
        end
    end
  module2467 #() modinst2805 (wire2804, clk, reg2293, reg976, reg2301, wire924, reg2291);
  always
    @(posedge clk) begin
      reg2806 <= $signed({reg2329});
      for (forvar2807 = (1'h0); (forvar2807 < (3'h5)); forvar2807 = (forvar2807 + (1'h1)))
        begin
          for (forvar2808 = (1'h0); (forvar2808 < (3'h4)); forvar2808 = (forvar2808 + (1'h1)))
            begin
              reg2809 <= $unsigned(reg1005);
              reg2810 <= (((~($signed(reg957) ?
                          wire2260[(3'h4):(2'h2)] : reg2307)) ?
                      reg2349 : $signed((7'h43))) ?
                  reg2340[(3'h7):(3'h7)] : (+wire1013[(3'h6):(1'h0)]));
              reg2811 <= ($unsigned((~reg2246[(4'hf):(4'h8)])) || $signed(reg2225[(5'h1c):(5'h19)]));
              reg2812 <= ((&$signed((~&(~reg2368)))) ?
                  (+(~^$unsigned((~wire2804)))) : (&((&(8'hbd)) & reg2457)));
              reg2813 = (7'h42);
              reg2814 <= $signed(($unsigned(reg2216[(4'he):(4'h8)]) << wire1772));
            end
          for (forvar2815 = (1'h0); (forvar2815 < (2'h3)); forvar2815 = (forvar2815 + (1'h1)))
            begin
              reg2816 <= (|reg2341);
            end
          reg2817 = reg936;
          reg2818 = reg985[(1'h0):(1'h0)];
          for (forvar2819 = (1'h0); (forvar2819 < (3'h5)); forvar2819 = (forvar2819 + (1'h1)))
            begin
              reg2820 = reg996[(2'h2):(1'h1)];
              reg2821 = (reg1357 ?
                  ($unsigned(wire924) ?
                      ($unsigned(reg2433[(4'ha):(2'h3)]) ?
                          reg2440 : $signed(reg2423)) : ((-reg2419) ~^ (8'haf))) : $unsigned(reg941));
              reg2822 <= {$signed((~^reg2455[(1'h1):(1'h0)]))};
              reg2823 <= $signed($signed((^~$unsigned(reg2321[(3'h7):(2'h3)]))));
              reg2824 = ($unsigned(reg2266[(3'h5):(3'h5)]) > wire2339);
              reg2825 = reg952[(1'h1):(1'h0)];
              reg2826 <= $signed(((^~reg2383[(5'h14):(4'h8)]) ?
                  (+(((8'haa) ^ reg2453) ?
                      {reg2433,
                          reg2427,
                          reg2309} : (~^wire2337))) : reg2309[(2'h3):(1'h1)]));
            end
          for (forvar2827 = (1'h0); (forvar2827 < (3'h5)); forvar2827 = (forvar2827 + (1'h1)))
            begin
              reg2828 <= {{reg2232}};
              reg2829 <= (~|$unsigned($signed({reg963, (8'hac)})));
              reg2830 = reg2360;
              reg2831 = (reg1347 ?
                  $signed($unsigned($unsigned(reg1043))) : (((&reg2383[(5'h19):(3'h5)]) ?
                          ((reg989 == reg2461) != (~wire926)) : reg997[(5'h13):(4'h8)]) ?
                      $signed(((reg2429 ? reg2223 : reg955) ?
                          forvar2808[(4'ha):(4'h8)] : (^~reg2404))) : $signed({(+reg2306),
                          reg2276,
                          (reg2267 ? reg2383 : reg2432)})));
              reg2832 = $signed($signed((^((reg2209 < wire1770) + $unsigned(reg1023)))));
            end
          if (forvar2815)
            begin
              reg2833 = ((reg1351 ?
                      $signed(((reg1025 < reg2380) ?
                          reg1346 : reg2316)) : $signed(reg2817)) ?
                  (reg1375[(4'h8):(1'h0)] ?
                      reg1333 : (reg2831[(2'h3):(2'h2)] ?
                          reg2217 : (-$unsigned(reg2832)))) : $signed($unsigned(reg1050)));
            end
          else
            begin
              reg2833 = (~(~reg959));
              reg2834 = $unsigned(reg1351[(4'hc):(1'h0)]);
              reg2835 <= $unsigned($signed((($unsigned(wire926) ?
                      (|reg2456) : (reg2816 * reg2398)) ?
                  reg2358 : wire2804)));
              reg2836 = reg1335;
              reg2837 = $signed(($unsigned($unsigned(((8'hb3) || reg2829))) > {{{reg1351,
                          reg2255},
                      (reg1344 ^ reg2298),
                      reg2390[(3'h7):(3'h5)]},
                  $unsigned({reg989, reg991, reg1046}),
                  $unsigned(reg997)}));
              reg2838 = reg2423[(3'h5):(3'h4)];
              reg2839 = reg1357;
            end
        end
      reg2840 = (-(^~(({reg1344, reg1344, reg2274} ?
          reg1335[(1'h0):(1'h0)] : (reg943 & reg979)) | (reg2398 ?
          (reg2274 * reg2831) : (~|reg2315)))));
      if ($unsigned($signed((+((^~reg1333) ^~ $signed(reg2396))))))
        begin
          reg2841 = (reg2298 >> ($unsigned($unsigned(reg978[(5'h1b):(1'h1)])) && (((-wire1013) <<< (reg2269 ?
              (8'ha3) : reg2302)) ^~ $unsigned(reg1335))));
          if ($unsigned((-reg1369)))
            begin
              reg2842 <= $signed($unsigned((^$unsigned({reg2223}))));
              reg2843 = $signed(reg2342);
              reg2844 = reg2306[(5'h14):(3'h7)];
              reg2845 <= ($unsigned(reg2825[(5'h10):(4'ha)]) ^~ (~|$signed(reg2833[(3'h7):(2'h3)])));
              reg2846 <= $unsigned($unsigned($unsigned($unsigned(reg988))));
              reg2847 = $unsigned($unsigned({$signed(((8'hbf) ?
                      reg2216 : reg2323)),
                  (reg2453 <<< {reg1050}),
                  $unsigned(((8'hb4) - reg2357))}));
            end
          else
            begin
              reg2842 <= ($signed(({$signed(reg2816)} || reg2390)) ?
                  ($unsigned((~|((8'h9c) ? reg2845 : reg1369))) ?
                      (&$signed((reg2296 != (8'ha7)))) : $unsigned($signed($signed(reg2451)))) : $signed((({reg2383,
                      reg2828} - ((7'h51) ^ reg2282)) || (reg2246[(3'h4):(3'h4)] || reg2385))));
              reg2843 = reg2415[(1'h1):(1'h0)];
              reg2845 <= reg2391[(4'hd):(4'ha)];
              reg2846 <= $unsigned(((((reg2222 ? reg1043 : (8'hb3)) ?
                      $signed((8'ha1)) : (reg2316 ?
                          reg1349 : reg1353)) < $unsigned({reg2440})) ?
                  $signed(((^~reg1346) ?
                      $unsigned(reg1370) : (reg2396 ?
                          reg2836 : reg2320))) : $unsigned({$unsigned((7'h40)),
                      reg2398[(4'h9):(4'h8)]})));
              reg2848 <= {{reg2297,
                      $signed({(~&reg1369)}),
                      {$unsigned(reg2812),
                          ((reg2199 <<< reg2359) ?
                              $signed(reg2209) : $unsigned(reg2269)),
                          reg2301[(4'h8):(3'h4)]}},
                  ((($unsigned(reg2290) ?
                          {(8'hae),
                              (7'h44)} : $unsigned((8'hae))) || $signed($signed(reg2296))) ?
                      reg2215 : $signed(($unsigned(wire1013) ?
                          (|reg986) : (reg995 ? reg2279 : reg2368)))),
                  (~(+reg1343[(2'h3):(2'h3)]))};
              reg2849 = (reg2447[(5'h12):(4'hc)] == reg2307[(2'h2):(2'h2)]);
            end
          for (forvar2850 = (1'h0); (forvar2850 < (3'h4)); forvar2850 = (forvar2850 + (1'h1)))
            begin
              reg2851 <= ((reg964 ?
                      ((-(^~reg1001)) ?
                          $signed((reg1338 ^ reg2222)) : $signed((wire928 << reg2271))) : reg1346) ?
                  (forvar2807[(2'h3):(2'h2)] <= (8'ha2)) : ($unsigned($signed((8'h9d))) ~^ ((reg2421 || (reg2818 ?
                      (7'h46) : reg1374)) == reg2228)));
              reg2852 = ((!reg2448[(3'h4):(2'h2)]) * reg2296);
              reg2853 <= reg2359;
              reg2854 <= (~^$unsigned($unsigned((!reg2823))));
              reg2855 = reg2387[(1'h0):(1'h0)];
              reg2856 = $signed({(((~&reg2432) ?
                          $unsigned(reg2415) : $unsigned(reg945)) ?
                      wire926[(1'h0):(1'h0)] : (|$unsigned(reg2270)))});
              reg2857 = {$unsigned(reg2433[(3'h5):(2'h2)]), reg2831, (7'h55)};
            end
        end
      else
        begin
          reg2841 = ((~|reg2306) <= $unsigned((^(|{reg1054}))));
          reg2843 = $signed((7'h46));
          reg2844 = (~(+reg2224));
        end
      reg2858 = ((((^~(+reg2323)) ?
          (!$unsigned(forvar2819)) : (^~reg2306)) ~^ {$unsigned((^reg2817))}) <<< (((~|$signed((7'h56))) ?
          reg2362 : $unsigned(reg936)) >> reg2285));
    end
  always
    @(posedge clk) begin
      if (reg2438[(5'h16):(5'h16)])
        begin
          if (reg981)
            begin
              reg2859 = (8'h9c);
              reg2860 = reg2248;
              reg2861 <= $unsigned(reg2271[(3'h5):(2'h2)]);
              reg2862 <= (~&$signed(reg2435));
              reg2863 <= (reg995[(2'h2):(1'h0)] ?
                  reg955 : (^$unsigned(((reg2427 ?
                      reg988 : reg2854) || $signed(reg2267)))));
              reg2864 <= (^~(reg979[(2'h3):(2'h2)] < (!(&{reg2427}))));
            end
          else
            begin
              reg2859 = (~&reg941);
              reg2860 = reg2862;
              reg2861 <= reg2438[(5'h10):(4'h9)];
              reg2862 <= reg1057[(3'h7):(3'h4)];
            end
          reg2865 <= reg941;
          if ((8'hb5))
            begin
              reg2866 <= (|$signed($unsigned(((^~reg2266) ?
                  (7'h4f) : (7'h41)))));
              reg2867 <= reg2286[(2'h3):(1'h1)];
              reg2868 = {(~($unsigned((reg2279 ? reg2292 : reg2449)) ?
                      (&(wire928 && (8'had))) : reg986))};
              reg2869 = ($signed(reg2868[(3'h7):(1'h0)]) ^ (&$unsigned(reg2209[(4'he):(3'h4)])));
            end
          else
            begin
              reg2868 = reg2867;
              reg2870 <= {$unsigned(((~(!reg2228)) ?
                      {(reg2264 ? reg2281 : reg991),
                          (reg1036 <= reg2387)} : reg957)),
                  $signed($signed(($signed(reg2246) ?
                      $signed(reg2267) : (^reg2202)))),
                  (!reg1343[(3'h5):(1'h1)])};
            end
        end
      else
        begin
          reg2859 = $unsigned($unsigned((reg1050[(4'hf):(3'h4)] > (reg2232[(5'h11):(3'h6)] ?
              ((7'h55) & reg2217) : (reg961 ? reg2265 : reg982)))));
          for (forvar2860 = (1'h0); (forvar2860 < (3'h5)); forvar2860 = (forvar2860 + (1'h1)))
            begin
              reg2868 = ((reg2435 | (&reg2814[(4'he):(4'hd)])) < (|$signed(reg2394)));
              reg2870 <= reg2405[(5'h10):(4'h8)];
              reg2871 = ($unsigned({reg2430,
                      {$unsigned(reg2279),
                          (reg2341 ? reg1036 : (7'h42)),
                          $unsigned(reg959)},
                      $signed(reg2342)}) ?
                  ((((|(7'h47)) ?
                              reg1025[(5'h14):(1'h1)] : (reg2217 >= reg1047)) ?
                          reg2228[(4'hb):(3'h4)] : reg2356[(3'h7):(3'h7)]) ?
                      ($signed((reg1047 != reg2411)) && ($unsigned(reg931) == $unsigned(reg2449))) : ((~&(reg2387 ?
                              reg2287 : wire1013)) ?
                          reg2286[(5'h11):(3'h7)] : $unsigned((reg1010 << reg2221)))) : ((((reg2415 >>> reg2404) ~^ $signed(reg1002)) || $unsigned((reg2869 ?
                      reg941 : reg1344))) ^ (reg2413 ?
                      {$unsigned(reg2232), (!reg2429)} : $unsigned((reg991 ?
                          reg1338 : (8'hba))))));
              reg2872 <= $signed(reg1054);
            end
          reg2873 <= ((reg2865 ?
              (reg2203 ?
                  (~&{reg990, (7'h56)}) : (~(7'h4a))) : ({(reg1050 == reg2449),
                      (reg2389 < reg996)} ?
                  ((reg2336 || reg2202) >>> (reg2826 ?
                      reg2296 : (8'hbb))) : ($unsigned(reg2328) << (reg985 ?
                      reg2315 : reg2429)))) != $signed((+reg988)));
          if (reg2329[(3'h4):(3'h4)])
            begin
              reg2874 <= reg2453[(5'h15):(4'hf)];
              reg2875 = reg1044;
              reg2876 = reg2307;
            end
          else
            begin
              reg2874 <= (!reg2872);
              reg2875 = $signed(reg2331[(5'h13):(4'h9)]);
              reg2876 = ({reg2812[(5'h12):(4'hf)]} ?
                  {(reg1347 == $unsigned(reg2297[(4'h9):(1'h0)])),
                      ((~^(reg2439 == reg2861)) ?
                          ((reg2283 ^~ wire2804) ?
                              reg2381 : reg1351[(3'h5):(3'h4)]) : {(~|(7'h4d)),
                              $signed(reg2452),
                              $unsigned(reg2810)})} : reg2854);
              reg2877 <= reg2453[(1'h0):(1'h0)];
              reg2878 <= ($unsigned(($unsigned((reg2221 ?
                      forvar2860 : reg1371)) ^~ {$signed((8'hbe)),
                      $unsigned(reg2423)})) ?
                  reg2285 : {$unsigned($signed((~|reg2347))),
                      ((reg2320[(5'h10):(4'ha)] ~^ reg1371[(2'h3):(1'h0)]) ?
                          reg964 : $signed(reg989[(1'h1):(1'h0)]))});
              reg2879 <= reg2866[(3'h7):(3'h5)];
            end
          reg2880 = ((-(~(+$signed(reg2851)))) * (reg2209 | (+$unsigned(reg2810[(5'h17):(2'h3)]))));
          reg2881 <= (^(reg1351[(4'hb):(4'ha)] < (reg2859 != reg985[(4'h9):(3'h4)])));
          for (forvar2882 = (1'h0); (forvar2882 < (2'h3)); forvar2882 = (forvar2882 + (1'h1)))
            begin
              reg2883 = reg2863[(4'hc):(2'h2)];
              reg2884 = $signed(reg994);
            end
        end
      if ((~{(((+reg2457) >= (reg985 ? reg2363 : reg2309)) ?
              (~$signed(reg978)) : (~(reg2865 ? wire2804 : reg2224))),
          forvar2860[(5'h16):(2'h2)],
          $signed($signed(reg2304))}))
        begin
          reg2885 = ($unsigned($unsigned((reg2319 ?
                  ((7'h4b) >>> forvar2882) : $unsigned(reg2809)))) ?
              ($unsigned($unsigned($signed((8'hbd)))) ?
                  $unsigned(reg2447[(4'h9):(1'h0)]) : (&reg2877[(4'h8):(2'h3)])) : $signed((+reg990[(4'ha):(1'h1)])));
          for (forvar2886 = (1'h0); (forvar2886 < (1'h0)); forvar2886 = (forvar2886 + (1'h1)))
            begin
              reg2887 <= reg2872;
              reg2888 <= $unsigned(reg2846);
              reg2889 = forvar2882;
              reg2890 = (($unsigned(reg2342[(3'h4):(1'h0)]) >> (((reg1347 <<< reg2880) ?
                  (reg2853 >>> reg2439) : (reg2845 ?
                      reg1010 : reg2223)) << $signed($unsigned(forvar2886)))) ^ ((~&{reg962,
                  (|reg2274)}) || (8'ha4)));
              reg2891 <= reg2877[(5'h11):(4'he)];
            end
          if ($unsigned((|$unsigned(((~|reg986) ?
              (reg2439 ? reg959 : reg2814) : reg2298[(1'h0):(1'h0)])))))
            begin
              reg2892 = $signed((reg2380 ?
                  ($signed(reg966) ?
                      reg2381 : (8'hb1)) : (reg2865[(2'h3):(1'h0)] ?
                      $unsigned($signed((8'ha0))) : reg2331)));
              reg2893 <= $signed((&($signed({reg1370,
                  reg2266}) && ($unsigned(reg1005) ?
                  $signed(reg2341) : reg2884[(1'h0):(1'h0)]))));
              reg2894 <= (~^$unsigned((~&((reg994 || reg2862) ?
                  reg2353[(1'h1):(1'h0)] : (reg2890 | reg2888)))));
              reg2895 <= ((reg2269 ?
                  reg2321 : ($unsigned(reg2865) ?
                      (((7'h56) ?
                          (8'ha2) : reg2853) > (reg982 >= reg1353)) : (reg2290[(4'h9):(2'h2)] - (7'h41)))) >= {($unsigned(reg961[(3'h7):(3'h4)]) ?
                      $signed((reg2223 ?
                          reg961 : reg2342)) : $unsigned((&reg957))),
                  (reg2341 ?
                      $signed($signed((8'hb1))) : (&(reg2388 ?
                          reg961 : reg1054)))});
            end
          else
            begin
              reg2892 = reg2230;
              reg2896 = ($signed(((reg2387[(5'h11):(3'h7)] ^~ reg2247) ?
                  $unsigned($signed(reg1338)) : reg2382)) && $signed(($signed($unsigned(reg2890)) ?
                  reg2347 : {((7'h56) ? reg2319 : (8'ha4))})));
              reg2897 <= reg2273;
            end
        end
      else
        begin
          for (forvar2885 = (1'h0); (forvar2885 < (1'h0)); forvar2885 = (forvar2885 + (1'h1)))
            begin
              reg2886 = (^(((!(+reg2814)) ?
                  ((reg2851 ^~ reg2320) ?
                      (reg1373 >= reg2453) : (~&reg2401)) : reg1036) - ({reg1005[(4'ha):(4'h9)],
                  reg1370[(3'h4):(1'h0)]} < reg1001[(2'h2):(2'h2)])));
              reg2887 <= (($signed($unsigned($signed((7'h4e)))) <<< reg1057[(4'ha):(4'ha)]) ?
                  (|({$unsigned(reg2296)} ?
                      (^~((8'h9e) + (8'ha5))) : ((reg978 ?
                          reg991 : reg2822) < (~|reg2302)))) : $unsigned((~|reg1025[(4'ha):(3'h7)])));
              reg2889 = $unsigned($signed({(8'ha3),
                  (~$signed(reg2423)),
                  ({reg2427, reg2358, reg2880} ^ (reg2265 ?
                      reg2826 : reg2362))}));
              reg2890 = (((($signed((8'hbb)) & reg2353) < $unsigned({reg2224})) * (7'h49)) * (!(reg1359 ?
                  $signed(((7'h4b) <<< reg2345)) : (^~{(7'h43),
                      reg2209,
                      reg2418}))));
              reg2891 <= ((reg2893 ?
                      $signed((-(!reg2394))) : {(reg2886[(4'he):(4'h8)] ?
                              (reg2848 >> reg2861) : ((7'h45) << reg995)),
                          (reg2894 >= (reg2224 || reg2427))}) ?
                  (({(^(7'h55))} ?
                      ((reg2449 ?
                          reg2276 : reg2889) + (-reg985)) : reg2460[(3'h5):(1'h0)]) >> (reg943[(3'h4):(1'h0)] ?
                      (8'ha2) : (reg2877[(3'h6):(1'h1)] ?
                          reg961[(4'h9):(4'h8)] : (wire1327 ?
                              reg2887 : reg2247)))) : {reg2274});
              reg2893 <= (7'h4e);
            end
          for (forvar2894 = (1'h0); (forvar2894 < (3'h4)); forvar2894 = (forvar2894 + (1'h1)))
            begin
              reg2895 <= {(|reg2853), (~reg982[(4'hb):(4'hb)]), (~&(7'h4b))};
              reg2896 = {({$unsigned($signed(reg2870)),
                      reg2267[(2'h2):(1'h1)]} || $unsigned(reg1353[(1'h1):(1'h0)]))};
              reg2898 = (reg2810 + (!$signed($signed($signed(reg2810)))));
              reg2899 <= $unsigned((~&reg979[(1'h1):(1'h0)]));
            end
          if ($unsigned(($signed((reg2345[(2'h3):(2'h2)] + reg2356)) & ((|{reg1374,
                  reg2385,
                  reg955}) ?
              (!{reg945}) : ({(7'h41)} ? (+reg2823) : (reg2382 >> reg1046))))))
            begin
              reg2900 = $signed($unsigned($unsigned(wire2338)));
              reg2901 = (($signed((((7'h4f) ?
                  (7'h47) : reg2321) + (reg2822 >>> reg1054))) || $unsigned(reg2835)) <<< $unsigned((^~((reg2427 < (8'h9c)) ^ (reg997 ?
                  (7'h43) : reg2895)))));
              reg2902 <= $unsigned($unsigned((reg2221 ?
                  reg933 : (|$signed(reg2421)))));
            end
          else
            begin
              reg2902 <= reg2826;
              reg2903 = $signed($unsigned({reg936, reg2439[(4'he):(4'hc)]}));
              reg2904 = $signed(((($signed(reg2461) ?
                      (reg2427 + reg2323) : wire926) && $signed((wire1013 ?
                      reg1343 : reg2881))) ?
                  (reg2292[(2'h3):(1'h0)] > ($unsigned(reg985) ?
                      reg2835[(4'h8):(1'h1)] : ((7'h4e) ?
                          reg2274 : reg2854))) : reg2829));
              reg2905 <= (!reg2336);
              reg2906 = reg2893[(4'hc):(4'ha)];
              reg2907 <= (^~((((reg2307 ?
                          reg2886 : reg966) << $unsigned((8'ha8))) ?
                      reg1370 : $unsigned(reg2874[(3'h7):(3'h5)])) ?
                  (reg2263 ?
                      (~|$unsigned(reg2319)) : $signed($signed(reg1343))) : (^reg2452)));
            end
          if ((8'ha4))
            begin
              reg2908 = reg2263[(5'h12):(4'ha)];
              reg2909 <= reg989;
              reg2910 = (((8'hbe) ?
                      ($signed(reg2230[(3'h4):(1'h0)]) + ({reg994} && (7'h51))) : $unsigned(((reg2902 ^~ reg1343) != $signed(reg2363)))) ?
                  wire2195[(1'h1):(1'h0)] : ((&(|(reg986 ? reg996 : (7'h53)))) ?
                      $signed((|{reg2889,
                          wire924})) : $unsigned($unsigned((forvar2882 ?
                          (8'hab) : reg1362)))));
            end
          else
            begin
              reg2908 = (!$signed(reg2264));
            end
        end
      reg2911 <= (((!$unsigned((7'h41))) == $unsigned((~$signed(reg2404)))) | $signed((({reg1036,
              reg972} != (^reg2870)) ?
          $signed(((7'h51) ?
              reg2885 : reg1345)) : $unsigned($signed(reg1344)))));
      for (forvar2912 = (1'h0); (forvar2912 < (2'h3)); forvar2912 = (forvar2912 + (1'h1)))
        begin
          if (reg2383)
            begin
              reg2913 <= reg2904;
              reg2914 = wire2260;
            end
          else
            begin
              reg2914 = ({((reg970[(1'h0):(1'h0)] ?
                          reg2449 : (reg2881 >>> (7'h47))) ?
                      (~&$unsigned(reg2336)) : reg2291),
                  (($unsigned((8'hba)) >> (reg1043 < reg2296)) ^~ reg1043),
                  (7'h4c)} >> (~&$signed(reg2320[(5'h11):(4'hc)])));
              reg2915 <= ((+reg1369) >> ($unsigned(reg2910) >> (!((reg932 ?
                      reg1044 : reg981) ?
                  ((8'hba) && reg2835) : $unsigned(reg2224)))));
              reg2916 <= (wire927[(4'h9):(2'h3)] ^~ (reg2255[(5'h1b):(2'h3)] ?
                  $unsigned(reg988) : ((reg2846[(4'hd):(3'h4)] == (reg1362 || reg1355)) - $unsigned(((8'hbb) ?
                      reg2903 : reg2868)))));
              reg2917 = {(&reg1002[(5'h14):(4'ha)]),
                  $unsigned(reg2307[(2'h2):(1'h1)]),
                  reg1370};
            end
          reg2918 <= (reg2903[(4'hd):(2'h2)] ?
              reg2286 : ((~|reg936[(1'h0):(1'h0)]) <<< ((reg2391[(5'h15):(1'h0)] * reg2222[(3'h6):(3'h4)]) >= ((reg2363 ?
                  reg2286 : reg2842) != $unsigned(reg2285)))));
          if (($signed(reg2217[(2'h2):(1'h1)]) * reg2321[(4'hd):(3'h5)]))
            begin
              reg2919 <= $signed({(~^{$unsigned((7'h43))}),
                  {((^reg2826) ? (~reg2907) : $signed(reg2360))},
                  {$unsigned($unsigned(reg2302)), (!$signed(reg2331))}});
            end
          else
            begin
              reg2919 <= reg2873;
              reg2920 = (8'hb8);
            end
          if ($signed({((~|$signed(reg2865)) ~^ ((reg2235 <= (8'ha4)) != (-reg989)))}))
            begin
              reg2921 = reg1355[(3'h7):(1'h0)];
              reg2922 = $unsigned((($unsigned((reg2230 ~^ wire2804)) ?
                      reg2263[(5'h11):(2'h2)] : reg1020[(5'h13):(2'h2)]) ?
                  reg2809 : reg2359));
              reg2923 = $unsigned((~&$unsigned((^(reg1001 ?
                  wire1772 : (8'haf))))));
            end
          else
            begin
              reg2924 <= {{reg2433[(4'hb):(3'h4)]},
                  reg2273[(4'ha):(3'h7)],
                  (~&reg2271[(2'h2):(1'h0)])};
              reg2925 = $unsigned(reg2432[(3'h5):(3'h5)]);
              reg2926 <= (forvar2885 << ($unsigned(($signed(reg2874) >= reg1043)) >= $signed(((!reg943) > (reg1044 || reg1351)))));
              reg2927 = $unsigned((reg994 ?
                  reg1333 : (reg940[(4'hd):(3'h4)] << (~reg2461))));
            end
          reg2928 <= (($signed(($unsigned(reg2296) | (reg2363 > reg2347))) <= reg2279[(3'h5):(1'h0)]) ?
              (-(&{(reg2898 << reg2413),
                  $signed(reg2264)})) : (reg1338[(4'h8):(4'h8)] == (($unsigned(reg2835) ?
                      $signed(wire2260) : reg2421[(2'h3):(2'h3)]) ?
                  $signed((reg1343 ?
                      reg2809 : reg1005)) : (reg2267 == (8'haf)))));
        end
      for (forvar2929 = (1'h0); (forvar2929 < (3'h4)); forvar2929 = (forvar2929 + (1'h1)))
        begin
          reg2930 = reg957[(5'h11):(1'h0)];
        end
      reg2931 = $signed((~&reg982[(2'h2):(1'h1)]));
    end
  always
    @(posedge clk) begin
      if (({((|reg2429[(2'h2):(2'h2)]) || ($signed(reg2341) ?
              (reg2440 - reg2315) : (reg2223 ? reg2842 : (8'ha7)))),
          {reg2873}} * (8'hbc)))
        begin
          if ((~$signed(($signed((reg2894 >> reg2810)) != (7'h56)))))
            begin
              reg2932 <= (&$signed({(~^(7'h45))}));
              reg2933 = $signed((reg2228[(4'hb):(3'h4)] ?
                  (!((reg1372 ?
                      reg2419 : (7'h49)) != reg2323)) : $signed(reg2209)));
              reg2934 = $signed($unsigned(reg1043[(2'h3):(2'h3)]));
              reg2935 <= $signed({(($unsigned(reg2307) + $signed(reg2874)) ?
                      ((reg2877 ? reg2911 : reg2398) ?
                          ((7'h51) >= reg978) : $signed(reg2826)) : $unsigned((wire928 & reg2265)))});
            end
          else
            begin
              reg2933 = (($signed((~^(reg2447 ? reg2302 : reg2269))) ?
                  ((~((8'hb1) << reg2202)) << reg994[(1'h0):(1'h0)]) : {((reg997 + reg2323) << (8'h9e)),
                      reg964}) || $unsigned($unsigned(((reg1355 ?
                      reg2934 : reg2867) ?
                  $signed((8'hbb)) : (reg2919 ? reg944 : reg2909)))));
              reg2934 = ({(&(8'had)),
                      (-reg2290),
                      (reg2413[(1'h0):(1'h0)] || ((reg2438 >> reg2866) ?
                          $unsigned(reg952) : $signed(reg2297)))} ?
                  ({($signed((8'hb5)) + reg985[(3'h7):(1'h1)]),
                      reg2286[(3'h6):(3'h4)]} >= $unsigned($signed(reg2230[(5'h10):(2'h2)]))) : $unsigned($signed(((reg2279 >> reg2449) || {reg2202,
                      (8'ha5),
                      reg1043}))));
              reg2935 <= reg2438;
              reg2936 <= (~&({((reg1375 ?
                          reg2224 : (8'hb3)) ~^ $unsigned(reg2916)),
                      $signed((reg2287 == reg2329)),
                      reg2918} ?
                  $unsigned((+reg2870)) : ((+(8'hbb)) ?
                      $signed((reg2870 ? reg2199 : (7'h41))) : (^reg966))));
            end
          if ((reg1036[(4'ha):(4'ha)] ?
              $signed(($signed((reg2307 < reg2319)) ~^ reg1338[(3'h7):(1'h1)])) : (wire1327[(5'h10):(4'h8)] ?
                  $signed(reg2926[(2'h2):(1'h0)]) : (~|reg2389[(3'h5):(3'h4)]))))
            begin
              reg2937 = (^~(reg1355[(1'h0):(1'h0)] ~^ (reg2292[(4'h8):(3'h5)] ?
                  reg932[(1'h1):(1'h0)] : reg2842[(4'hc):(2'h2)])));
              reg2938 = reg2897[(3'h5):(1'h0)];
              reg2939 = ((&((7'h53) <= $signed($signed((8'hb3))))) - reg1357);
              reg2940 = (^~$signed($unsigned(((8'hbc) <<< reg2360))));
              reg2941 = {reg1057[(4'hc):(3'h7)], reg1374[(4'hd):(1'h0)]};
              reg2942 <= $signed(reg2309[(2'h2):(2'h2)]);
            end
          else
            begin
              reg2937 = ($signed(($unsigned({reg2881}) ?
                  $signed((reg2315 <<< (7'h44))) : {(&reg1043),
                      $signed((8'haf)),
                      $unsigned(reg2447)})) || ($signed(reg959[(5'h1b):(4'ha)]) ?
                  (^(~reg991)) : reg2248[(4'hf):(4'he)]));
              reg2942 <= reg2309;
              reg2943 = $unsigned((reg2320[(4'h8):(4'h8)] ?
                  (-(wire1327[(5'h13):(4'h9)] ?
                      {reg1353,
                          reg955,
                          wire928} : reg1338[(1'h1):(1'h1)])) : (8'haf)));
              reg2944 = {(^$unsigned(reg2419[(5'h19):(5'h17)])),
                  ($signed(({reg1009} ?
                          (reg978 ? reg2457 : reg941) : (reg2902 ?
                              (7'h58) : (8'hb6)))) ?
                      $signed($signed(reg2845)) : {reg2263,
                          (((8'had) >>> reg985) ? reg2199 : (~|(8'ha4))),
                          ($unsigned(reg2296) ?
                              (reg2368 != reg2928) : $signed(reg2225))}),
                  (|(reg2242 ?
                      (^$signed(reg989)) : {(^reg991),
                          {(7'h53), reg2902},
                          reg1372[(2'h3):(1'h1)]}))};
              reg2945 = (reg2453 ?
                  reg2822 : (~(($unsigned(reg2433) ?
                      (reg2297 * reg2887) : (-reg2940)) >> reg1345)));
              reg2946 <= $unsigned(($unsigned((^~{reg2389})) + reg2826));
            end
          reg2947 <= reg2234;
          for (forvar2948 = (1'h0); (forvar2948 < (1'h1)); forvar2948 = (forvar2948 + (1'h1)))
            begin
              reg2949 = ({$unsigned(reg997[(2'h3):(2'h2)]),
                      $unsigned((~reg2897[(5'h10):(3'h4)])),
                      reg2273[(4'he):(1'h0)]} ?
                  (~^$unsigned($signed($unsigned((8'h9f))))) : {((~&(reg2418 ?
                          reg2285 : reg2224)) <= ((reg2297 * reg988) ^~ $signed(reg2867))),
                      $signed({(-reg1355)}),
                      ($signed(((7'h47) >= (7'h52))) << $signed(wire928))});
              reg2950 = ((~|((~|(reg1343 ?
                      reg2268 : reg2865)) >>> reg1359[(5'h12):(4'hd)])) ?
                  (&reg1044) : (~^$signed($unsigned((^reg978)))));
              reg2951 <= $signed($unsigned((reg2439[(5'h19):(5'h11)] - ($unsigned(reg2950) << $signed(reg2853)))));
              reg2952 = (8'hb7);
              reg2953 <= $signed((!$unsigned(((+reg1339) || (reg2228 + reg2235)))));
            end
          reg2954 <= {$signed({$unsigned(((7'h50) - reg1023)),
                  $unsigned((reg2909 ? reg2877 : reg997)),
                  ($signed((8'ha9)) ? (reg994 ? (8'had) : reg2861) : reg2276)}),
              ((((reg2274 ? reg972 : reg985) && $unsigned(reg995)) == (reg2405 ?
                  $signed((8'h9e)) : reg2418[(1'h1):(1'h1)])) ^ $unsigned(((~^reg956) ?
                  (wire925 ? reg2854 : reg2247) : reg1057))),
              $signed((($unsigned(reg978) & $unsigned(reg2405)) ?
                  reg2281[(1'h1):(1'h0)] : $unsigned($signed(reg2202))))};
          reg2955 <= {(+(^((reg2405 != reg2223) ?
                  (^reg941) : reg2814[(1'h0):(1'h0)]))),
              $unsigned($signed(($unsigned(reg2234) >> $signed(reg2230))))};
        end
      else
        begin
          reg2933 = $signed(reg2398[(4'hb):(4'h9)]);
        end
      for (forvar2956 = (1'h0); (forvar2956 < (3'h5)); forvar2956 = (forvar2956 + (1'h1)))
        begin
          if ((|$unsigned($signed(reg2282[(4'h8):(3'h6)]))))
            begin
              reg2957 = {$unsigned((~&(-$signed(reg2359)))),
                  (((~$unsigned(reg955)) ?
                      ($signed(reg2320) ?
                          $signed(reg2378) : (reg2357 ?
                              reg1375 : (8'hba))) : reg2228[(5'h11):(4'he)]) || reg2293[(4'hb):(3'h6)])};
              reg2958 <= (|$signed($unsigned(reg2342[(2'h2):(2'h2)])));
              reg2959 = ((($unsigned((+reg944)) ?
                      (reg2428 ?
                          (reg2228 ?
                              (8'hac) : reg2265) : (reg2439 >> (8'had))) : (7'h57)) ^ $signed(({reg2304,
                      (7'h4e)} | (~reg2913)))) ?
                  ((&($unsigned((8'hb6)) >> $signed(reg931))) ?
                      reg2878[(2'h3):(1'h1)] : (~&({reg979, reg2404} ?
                          (wire2804 < (8'ha8)) : (reg2891 >= (8'ha5))))) : $signed($unsigned((reg1010 ?
                      $unsigned(reg961) : reg1372))));
              reg2960 <= reg2321;
              reg2961 <= $signed($signed($unsigned((wire1327[(3'h6):(3'h6)] ?
                  (reg970 * reg2959) : reg2230))));
              reg2962 <= (!reg2419[(1'h0):(1'h0)]);
            end
          else
            begin
              reg2957 = reg2213[(3'h4):(1'h1)];
              reg2959 = reg2296;
              reg2960 <= ($unsigned($signed(reg2421)) ?
                  ({reg2873} & ($unsigned((-reg2909)) ?
                      {(reg2907 ?
                              reg2806 : reg2344)} : $unsigned((~reg2283)))) : reg2382[(4'he):(2'h3)]);
              reg2961 <= $signed(reg2309[(1'h0):(1'h0)]);
            end
          reg2963 = $unsigned(reg2268[(5'h11):(4'hb)]);
          reg2964 <= reg2394[(4'hb):(3'h4)];
          reg2965 = (wire924[(2'h3):(2'h3)] - (~&$unsigned(reg2301[(5'h10):(4'hc)])));
          reg2966 <= {{($unsigned($unsigned(reg1333)) >= reg2315[(1'h0):(1'h0)]),
                  $unsigned({(!reg2907),
                      $unsigned((7'h4d)),
                      (reg2835 ? reg995 : reg1052)}),
                  reg2385}};
          for (forvar2967 = (1'h0); (forvar2967 < (2'h3)); forvar2967 = (forvar2967 + (1'h1)))
            begin
              reg2968 <= ((~|((reg2235[(4'hc):(2'h3)] ?
                  reg2401 : wire2804) < $signed($unsigned(reg2965)))) + ((^reg1338[(3'h4):(2'h2)]) ?
                  reg1343 : ((7'h40) * reg2954[(4'hd):(3'h7)])));
              reg2969 = $signed(((^~$unsigned($signed(reg2285))) ?
                  reg2811[(5'h1d):(5'h1b)] : (-$signed(reg2203))));
              reg2970 = ({(({reg2947, reg1349, reg2430} ?
                      $unsigned(reg2425) : (reg2307 < reg1005)) - reg2853),
                  $signed((reg2301 ?
                      reg2268 : $unsigned(reg2949)))} != reg2235[(5'h12):(3'h4)]);
              reg2971 <= reg2290;
              reg2972 <= reg970[(3'h6):(1'h0)];
              reg2973 <= ((!reg2281[(5'h16):(1'h1)]) ^~ (7'h45));
            end
          if ($unsigned(($unsigned(($unsigned(reg2455) < $signed(reg2263))) <= (8'hba))))
            begin
              reg2974 <= {reg2826,
                  ((((reg2268 ? reg2307 : reg972) ^~ $unsigned(reg2347)) ?
                          (reg1375 <= reg2264[(4'hf):(4'hd)]) : reg1373[(2'h3):(1'h1)]) ?
                      reg2822 : (~reg2344))};
            end
          else
            begin
              reg2975 = (~(~&$signed({$signed(reg2342),
                  (reg990 ? reg2945 : reg956),
                  ((8'hbf) ? reg2312 : reg2811)})));
              reg2976 = $unsigned((!$signed({(reg2312 <= (7'h4e)),
                  reg2242[(4'hc):(3'h6)]})));
              reg2977 <= reg2234;
              reg2978 = (~^$unsigned(reg1001));
              reg2979 <= reg2413;
              reg2980 = reg2428[(1'h0):(1'h0)];
            end
        end
      for (forvar2981 = (1'h0); (forvar2981 < (3'h6)); forvar2981 = (forvar2981 + (1'h1)))
        begin
          reg2982 <= $unsigned($unsigned($unsigned(((-(7'h47)) <= {reg2429,
              reg989,
              (7'h48)}))));
          reg2983 <= $unsigned((~^(&(reg2440 ?
              $signed(reg1374) : (reg2224 < reg2934)))));
          reg2984 <= reg2388[(3'h5):(2'h3)];
          if (($signed(reg2835[(3'h4):(1'h0)]) ?
              $unsigned(reg932[(2'h2):(1'h0)]) : {{$signed((8'haf)),
                      $signed(reg2452[(3'h6):(1'h1)])},
                  (8'hbd),
                  ({(reg2440 >>> reg2312)} <= reg1057[(4'hc):(3'h5)])}))
            begin
              reg2985 = $signed({$signed(reg2461[(5'h1c):(5'h15)]),
                  {$signed((reg2894 ? reg2248 : reg2389)),
                      reg940[(4'h9):(3'h7)],
                      {$signed(reg1057)}},
                  $unsigned($unsigned((&reg2810)))});
              reg2986 = $unsigned({$unsigned(reg2816[(1'h1):(1'h0)])});
            end
          else
            begin
              reg2987 <= $signed((wire926[(2'h3):(2'h3)] > ((reg2360[(5'h14):(2'h2)] << $signed(reg2842)) >>> reg2358)));
              reg2988 = (+reg933);
              reg2989 = reg979[(1'h0):(1'h0)];
              reg2990 <= ($unsigned((reg2881 ?
                      $signed(reg2356[(4'ha):(1'h0)]) : reg1371)) ?
                  (7'h50) : ((~|$unsigned($unsigned(reg2958))) && {(7'h48),
                      (7'h45)}));
              reg2991 <= ({(&(&(^reg963))), reg2899[(5'h17):(1'h1)]} ?
                  ($unsigned($signed((wire2260 ?
                      reg2961 : reg2864))) && (~|{$signed(reg1052),
                      (reg2897 ? reg2359 : reg1043)})) : reg2937);
              reg2992 <= reg2816;
            end
          for (forvar2993 = (1'h0); (forvar2993 < (1'h1)); forvar2993 = (forvar2993 + (1'h1)))
            begin
              reg2994 = ((reg2320[(2'h3):(2'h2)] * (~^($signed(reg932) > $signed((7'h57))))) >>> reg1333);
              reg2995 <= reg2448[(4'hd):(4'h8)];
            end
        end
      reg2996 <= ((reg2230[(5'h10):(1'h1)] || ($unsigned(reg2271) ?
              ($signed(reg2425) ?
                  reg2986 : ((7'h46) >= reg996)) : $unsigned($signed(reg1374)))) ?
          (reg933 != (reg2891 & reg1349)) : $signed((|forvar2948)));
      for (forvar2997 = (1'h0); (forvar2997 < (3'h4)); forvar2997 = (forvar2997 + (1'h1)))
        begin
          reg2998 = $unsigned((($signed(reg1333) == (^{reg2457})) ?
              (^~$signed((-reg2423))) : $unsigned(((reg2281 ?
                      wire926 : reg2344) ?
                  (~reg2822) : $unsigned(reg2881)))));
          for (forvar2999 = (1'h0); (forvar2999 < (1'h1)); forvar2999 = (forvar2999 + (1'h1)))
            begin
              reg3000 = ({(^(8'hac)),
                  (|($unsigned(reg1372) ~^ $unsigned(reg1351))),
                  reg2864} <<< reg2907[(3'h4):(1'h1)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg3001 = reg1373;
      reg3002 <= reg2439[(5'h12):(4'h9)];
      reg3003 = $signed($unsigned($unsigned(reg2991)));
      reg3004 <= reg2891[(2'h3):(1'h0)];
      if ($signed(wire2337[(3'h4):(1'h0)]))
        begin
          for (forvar3005 = (1'h0); (forvar3005 < (1'h0)); forvar3005 = (forvar3005 + (1'h1)))
            begin
              reg3006 = (reg2854 != reg2873);
              reg3007 = $unsigned(reg2336);
            end
        end
      else
        begin
          reg3005 = ($unsigned(((^~{reg1351, reg2461, reg2951}) ?
                  $unsigned((|reg979)) : $signed(reg997[(2'h2):(1'h1)]))) ?
              ($unsigned(reg2851) ?
                  reg2421[(2'h3):(1'h0)] : reg1054) : reg3007);
          for (forvar3006 = (1'h0); (forvar3006 < (2'h2)); forvar3006 = (forvar3006 + (1'h1)))
            begin
              reg3008 <= reg2222;
              reg3009 = (($signed((reg2419 ^ reg2862[(5'h11):(4'ha)])) ?
                      reg1353[(2'h3):(1'h1)] : $unsigned($unsigned((reg1345 ?
                          reg2356 : reg2347)))) ?
                  (~^reg2396) : $signed($signed(((!reg2360) ?
                      (8'hb1) : reg952[(4'h9):(3'h7)]))));
              reg3010 <= reg2328[(3'h7):(3'h6)];
              reg3011 <= reg2893[(5'h10):(3'h7)];
              reg3012 = (reg1346[(2'h2):(2'h2)] ?
                  $unsigned(((reg1010[(2'h2):(1'h0)] - reg2874) ?
                      reg2268[(5'h13):(4'h9)] : reg2811[(5'h10):(4'h9)])) : (reg2344 ^ (~^$signed((reg3005 + (7'h56))))));
              reg3013 = reg2924;
            end
          reg3014 <= $signed(($signed(reg2447[(5'h15):(3'h5)]) < (&(+$unsigned((8'hb6))))));
          for (forvar3015 = (1'h0); (forvar3015 < (3'h6)); forvar3015 = (forvar3015 + (1'h1)))
            begin
              reg3016 <= reg944[(2'h2):(2'h2)];
              reg3017 <= ({($unsigned((7'h42)) + wire927),
                  $unsigned($unsigned((wire1327 ? reg2316 : reg2453))),
                  reg3004} | $unsigned($unsigned($unsigned((reg3005 ^ reg2363)))));
              reg3018 = reg2897;
              reg3019 = reg2282[(5'h1a):(5'h15)];
              reg3020 <= {$unsigned($unsigned($unsigned((reg3010 ?
                      reg2306 : reg2810)))),
                  $unsigned((((^~reg2248) ^~ $signed(reg2312)) == reg2349))};
              reg3021 = ({(8'h9d)} ?
                  reg2344[(3'h4):(2'h3)] : ((&reg2432[(4'ha):(4'h9)]) ?
                      (reg1002[(3'h5):(2'h2)] ?
                          $signed($signed(reg2814)) : (+(|reg1052))) : (reg2926 ^ ($signed(reg2992) ?
                          $unsigned(reg2264) : $unsigned(reg2971)))));
              reg3022 = $signed({((~&reg2387) + reg2893),
                  {$signed((|wire2339)),
                      reg2954[(1'h1):(1'h1)],
                      ((reg2996 ~^ reg1359) ?
                          (reg2319 - (7'h4f)) : (reg2356 ^ (7'h47)))}});
            end
          for (forvar3023 = (1'h0); (forvar3023 < (3'h6)); forvar3023 = (forvar3023 + (1'h1)))
            begin
              reg3024 <= (~|$unsigned((forvar3006[(2'h3):(1'h0)] | (((7'h54) ?
                  (8'hac) : reg2276) ^ (~^reg2216)))));
              reg3025 = $unsigned($signed({({reg2829, reg1044, reg2331} ?
                      (+reg2879) : (reg3003 ? reg933 : reg2415)),
                  {(reg2960 ? reg2336 : reg2902),
                      ((7'h45) ? (7'h46) : reg2283),
                      reg2456},
                  $signed($signed(reg2991))}));
            end
        end
    end
  always
    @(posedge clk) begin
      reg3026 <= reg2887[(5'h17):(2'h2)];
      if ({($signed({(&reg981),
                  reg1036[(5'h17):(5'h15)],
                  (reg2413 ? wire2338 : reg2992)}) ?
              (8'hb2) : (reg2996[(5'h13):(3'h7)] >= (8'hac))),
          (reg1344 ~^ reg931[(1'h0):(1'h0)])})
        begin
          reg3027 <= (reg2380[(1'h0):(1'h0)] >> (-reg943));
          reg3028 = reg2292[(3'h4):(2'h2)];
          reg3029 = ((reg2276[(4'ha):(4'h9)] <= ($signed(reg2911[(5'h13):(4'h9)]) ~^ reg2863[(5'h1b):(5'h1a)])) ?
              $signed((reg1372 - (!reg2995))) : reg2270);
          reg3030 <= $signed(((reg2983[(5'h16):(3'h6)] ?
                  ((reg1370 <<< reg2895) > (~^reg2216)) : ($signed(reg936) ?
                      $signed((7'h54)) : (^reg2895))) ?
              (~|((&reg2381) & (reg991 >> reg2357))) : $signed($signed(reg2378[(3'h7):(2'h2)]))));
          for (forvar3031 = (1'h0); (forvar3031 < (3'h4)); forvar3031 = (forvar3031 + (1'h1)))
            begin
              reg3032 <= $unsigned(reg2448);
              reg3033 <= $signed($signed(reg2918));
              reg3034 <= reg2848[(5'h15):(4'hc)];
            end
          reg3035 <= reg940;
          reg3036 <= $signed(reg976[(5'h10):(3'h5)]);
        end
      else
        begin
          reg3028 = (~^reg2448[(4'ha):(4'h9)]);
        end
      reg3037 = (7'h46);
      for (forvar3038 = (1'h0); (forvar3038 < (3'h5)); forvar3038 = (forvar3038 + (1'h1)))
        begin
          if ($unsigned(reg2292[(4'hb):(2'h3)]))
            begin
              reg3039 = (((7'h40) ?
                  reg2954 : $unsigned((!$signed(wire1013)))) > ((~($unsigned(reg2290) ?
                  $unsigned(reg933) : (reg2202 ?
                      reg2457 : reg2391))) & {reg2835}));
              reg3040 <= $signed((reg2816[(3'h5):(2'h2)] ?
                  $unsigned($signed(reg2291)) : ($unsigned(((7'h58) - reg955)) ?
                      $unsigned($unsigned(reg2453)) : $signed(reg3010))));
              reg3041 = (((reg2302[(1'h0):(1'h0)] ?
                  ($unsigned(reg2955) & {(8'hbc),
                      reg2436,
                      (8'ha3)}) : (8'hb1)) == (~(^(reg2983 ?
                  reg2297 : reg2358)))) >>> ((~reg1345) ~^ (reg3037 & (reg2425[(3'h4):(2'h3)] > (reg940 <= reg2323)))));
              reg3042 <= ((reg2362[(5'h1a):(5'h12)] == reg2276[(5'h16):(5'h13)]) ?
                  (reg932[(4'hb):(4'hb)] == $signed($unsigned(reg2381))) : ($signed($signed(reg2816[(5'h17):(5'h15)])) ?
                      (reg1036 || (!reg2362[(4'hf):(4'he)])) : {(7'h47),
                          $unsigned({reg2383, wire926})}));
            end
          else
            begin
              reg3039 = $unsigned((((reg1346[(1'h1):(1'h0)] >>> {(7'h50),
                          reg2874}) ?
                      (reg2982[(4'h8):(2'h3)] >= {reg2428,
                          reg2232}) : ((reg2812 ? reg1009 : reg2235) ?
                          (^reg3041) : {reg2270, (7'h4d)})) ?
                  (&($unsigned(reg2306) ?
                      $signed(reg2987) : $unsigned(reg2977))) : (-$unsigned((reg2270 ?
                      reg2327 : reg2398)))));
            end
        end
      reg3043 <= (((&((reg2958 && reg2382) ?
          (-reg936) : $signed(reg2461))) <<< wire1772) ~^ reg991[(1'h1):(1'h1)]);
      if (($unsigned(((+$signed((8'hba))) ?
              reg2907[(4'he):(3'h4)] : ((reg2864 >> reg2341) | {reg2864}))) ?
          reg2968[(4'ha):(1'h0)] : ((8'hb4) ?
              {(reg2269[(1'h1):(1'h1)] ^ reg2342),
                  reg2425} : reg2301[(3'h6):(3'h6)])))
        begin
          reg3044 <= (~|$signed($unsigned(((7'h4c) ?
              $signed(reg2962) : $signed((8'hb5))))));
          reg3045 <= wire924;
          reg3046 = $unsigned($signed($signed(reg2814[(5'h13):(5'h13)])));
        end
      else
        begin
          for (forvar3044 = (1'h0); (forvar3044 < (1'h0)); forvar3044 = (forvar3044 + (1'h1)))
            begin
              reg3046 = ((reg3027[(5'h12):(4'h9)] ?
                      {reg2983[(5'h18):(4'h9)]} : ((!(^(8'hb7))) >= reg1351[(4'hd):(4'hd)])) ?
                  (&reg2928) : reg2449[(2'h2):(2'h2)]);
              reg3047 = $unsigned($unsigned((reg3017[(4'hf):(1'h0)] ?
                  reg2285[(3'h7):(1'h0)] : reg3044[(2'h3):(1'h0)])));
              reg3048 <= $unsigned(reg2953[(4'h8):(1'h0)]);
            end
          reg3049 <= reg2425[(3'h4):(2'h2)];
          for (forvar3050 = (1'h0); (forvar3050 < (3'h6)); forvar3050 = (forvar3050 + (1'h1)))
            begin
              reg3051 <= ($signed($unsigned(wire2195[(4'h9):(1'h0)])) << $unsigned(reg2329[(3'h5):(3'h4)]));
              reg3052 = (~^forvar3044);
              reg3053 = reg1351[(4'he):(2'h2)];
              reg3054 <= reg2263;
              reg3055 <= reg1047;
              reg3056 = (~|(($signed((|reg2872)) >> (-$signed(reg2331))) ?
                  (reg3051[(1'h0):(1'h0)] || reg959) : $unsigned($unsigned($signed(reg2301)))));
            end
        end
      if (reg2990[(3'h7):(1'h0)])
        begin
          for (forvar3057 = (1'h0); (forvar3057 < (2'h3)); forvar3057 = (forvar3057 + (1'h1)))
            begin
              reg3058 <= reg2230[(2'h2):(1'h0)];
              reg3059 <= (((^~reg2809) * ($signed($unsigned((7'h48))) ?
                  (^~reg2947) : reg2396[(3'h6):(1'h0)])) >= $unsigned((^reg2360)));
            end
        end
      else
        begin
          for (forvar3057 = (1'h0); (forvar3057 < (3'h4)); forvar3057 = (forvar3057 + (1'h1)))
            begin
              reg3060 = (~^(+$unsigned((+reg2438))));
              reg3061 = $unsigned($unsigned((reg2255[(5'h1c):(2'h3)] >> $signed(reg2293[(3'h6):(2'h3)]))));
            end
          reg3062 <= ($signed(wire2339[(1'h0):(1'h0)]) > reg2447[(5'h15):(2'h3)]);
          reg3063 = reg2853[(2'h2):(1'h1)];
        end
    end
  module1773 #() modinst3065 (.wire1778(reg976), .wire1776(wire2337), .y(wire3064), .wire1774(reg3058), .wire1777(reg2990), .wire1775(reg2984), .clk(clk));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module71
#(parameter param843 = ({(~|(((8'hb0) <<< (7'h58)) ? ((7'h4a) * (8'ha5)) : ((8'hb5) == (8'h9e))))} ? {(|({(8'ha6), (7'h4a)} ? ((7'h55) == (7'h50)) : ((8'hb0) | (8'hb8)))), (^~(((7'h57) ? (8'ha3) : (8'hb9)) ? ((7'h47) && (8'ha0)) : (~&(8'hbb)))), {(~&(^~(7'h4b)))}} : {{(((8'h9f) <= (8'hb8)) <= (&(7'h40))), (8'hbb), (((7'h41) ? (8'h9f) : (7'h50)) ? ((8'ha5) ^~ (8'hb8)) : ((8'hb6) ? (7'h48) : (7'h4e)))}}))
(y, clk, wire77, wire76, wire75, wire74, wire73, wire72);
  output wire [(32'h1c04):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire77;
  input wire [(2'h2):(1'h0)] wire76;
  input wire signed [(4'hf):(1'h0)] wire75;
  input wire signed [(3'h4):(1'h0)] wire74;
  input wire signed [(2'h3):(1'h0)] wire73;
  input wire [(5'h11):(1'h0)] wire72;
  wire [(5'h16):(1'h0)] wire842;
  wire [(4'hb):(1'h0)] wire840;
  wire signed [(5'h1c):(1'h0)] wire730;
  wire signed [(4'he):(1'h0)] wire683;
  wire [(5'h16):(1'h0)] wire241;
  wire signed [(5'h1d):(1'h0)] wire240;
  wire signed [(4'hc):(1'h0)] wire164;
  wire [(4'hf):(1'h0)] wire163;
  wire [(3'h7):(1'h0)] wire79;
  wire [(4'hd):(1'h0)] wire78;
  reg signed [(2'h3):(1'h0)] reg841 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg837 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg836 = (1'h0);
  reg [(4'ha):(1'h0)] reg835 = (1'h0);
  reg [(5'h12):(1'h0)] reg833 = (1'h0);
  reg [(5'h14):(1'h0)] reg827 = (1'h0);
  reg [(4'h8):(1'h0)] reg825 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg824 = (1'h0);
  reg [(3'h6):(1'h0)] reg822 = (1'h0);
  reg [(3'h5):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg818 = (1'h0);
  reg [(4'hf):(1'h0)] reg814 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg813 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg811 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg809 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg808 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg807 = (1'h0);
  reg [(5'h17):(1'h0)] reg806 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg805 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg803 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg802 = (1'h0);
  reg [(2'h3):(1'h0)] reg800 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg799 = (1'h0);
  reg [(5'h17):(1'h0)] reg793 = (1'h0);
  reg [(2'h3):(1'h0)] reg791 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg784 = (1'h0);
  reg [(4'he):(1'h0)] reg783 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg782 = (1'h0);
  reg [(4'hb):(1'h0)] reg781 = (1'h0);
  reg [(2'h3):(1'h0)] reg776 = (1'h0);
  reg [(3'h6):(1'h0)] reg775 = (1'h0);
  reg [(5'h19):(1'h0)] reg773 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg772 = (1'h0);
  reg [(5'h17):(1'h0)] reg771 = (1'h0);
  reg [(5'h15):(1'h0)] reg770 = (1'h0);
  reg [(4'hd):(1'h0)] reg768 = (1'h0);
  reg [(5'h1e):(1'h0)] reg764 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg763 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg757 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg756 = (1'h0);
  reg [(5'h17):(1'h0)] reg746 = (1'h0);
  reg [(2'h2):(1'h0)] reg743 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg742 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg741 = (1'h0);
  reg [(3'h4):(1'h0)] reg740 = (1'h0);
  reg [(4'he):(1'h0)] reg737 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg735 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg728 = (1'h0);
  reg [(4'hc):(1'h0)] reg727 = (1'h0);
  reg [(4'hb):(1'h0)] reg724 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg723 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg719 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg718 = (1'h0);
  reg [(5'h1b):(1'h0)] reg716 = (1'h0);
  reg [(4'h8):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg714 = (1'h0);
  reg [(5'h16):(1'h0)] reg711 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg708 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg705 = (1'h0);
  reg [(5'h17):(1'h0)] reg701 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg699 = (1'h0);
  reg [(5'h12):(1'h0)] reg687 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg696 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg695 = (1'h0);
  reg [(5'h12):(1'h0)] reg692 = (1'h0);
  reg [(5'h11):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg90 = (1'h0);
  reg [(5'h12):(1'h0)] reg98 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg102 = (1'h0);
  reg [(5'h16):(1'h0)] reg104 = (1'h0);
  reg [(5'h10):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg111 = (1'h0);
  reg [(5'h1f):(1'h0)] reg113 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg115 = (1'h0);
  reg [(5'h18):(1'h0)] reg117 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg121 = (1'h0);
  reg [(5'h1c):(1'h0)] reg125 = (1'h0);
  reg [(5'h14):(1'h0)] reg129 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg130 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg133 = (1'h0);
  reg [(4'hc):(1'h0)] reg134 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg135 = (1'h0);
  reg [(2'h3):(1'h0)] reg136 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg141 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg142 = (1'h0);
  reg [(5'h14):(1'h0)] reg145 = (1'h0);
  reg [(3'h7):(1'h0)] reg151 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg152 = (1'h0);
  reg [(5'h1b):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg162 = (1'h0);
  reg [(5'h1a):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg167 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg168 = (1'h0);
  reg [(5'h16):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg182 = (1'h0);
  reg [(5'h19):(1'h0)] reg186 = (1'h0);
  reg [(4'hc):(1'h0)] reg191 = (1'h0);
  reg [(5'h1d):(1'h0)] reg178 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg194 = (1'h0);
  reg [(5'h15):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg200 = (1'h0);
  reg [(2'h2):(1'h0)] reg201 = (1'h0);
  reg [(4'h9):(1'h0)] reg204 = (1'h0);
  reg [(5'h14):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg206 = (1'h0);
  reg [(5'h13):(1'h0)] reg209 = (1'h0);
  reg [(4'h9):(1'h0)] reg210 = (1'h0);
  reg [(5'h12):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg218 = (1'h0);
  reg [(5'h1e):(1'h0)] reg219 = (1'h0);
  reg [(5'h11):(1'h0)] reg222 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg227 = (1'h0);
  reg [(2'h3):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg232 = (1'h0);
  reg [(4'hb):(1'h0)] reg233 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg234 = (1'h0);
  reg [(5'h12):(1'h0)] reg239 = (1'h0);
  reg [(4'h9):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg251 = (1'h0);
  reg [(5'h15):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg255 = (1'h0);
  reg [(4'hf):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg257 = (1'h0);
  reg [(3'h5):(1'h0)] reg258 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg263 = (1'h0);
  reg signed [(4'he):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg266 = (1'h0);
  reg [(3'h4):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg269 = (1'h0);
  reg [(4'hf):(1'h0)] reg270 = (1'h0);
  reg [(2'h2):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg275 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg276 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg279 = (1'h0);
  reg [(4'h9):(1'h0)] reg281 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg283 = (1'h0);
  reg [(4'he):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg291 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg293 = (1'h0);
  reg [(5'h16):(1'h0)] reg295 = (1'h0);
  reg [(2'h2):(1'h0)] reg296 = (1'h0);
  reg [(4'hd):(1'h0)] reg299 = (1'h0);
  reg [(5'h10):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg304 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg307 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg311 = (1'h0);
  reg [(4'hf):(1'h0)] reg312 = (1'h0);
  reg [(5'h10):(1'h0)] reg313 = (1'h0);
  reg [(5'h18):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg315 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg320 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg321 = (1'h0);
  reg [(4'h9):(1'h0)] reg322 = (1'h0);
  reg [(4'h8):(1'h0)] reg324 = (1'h0);
  reg [(4'ha):(1'h0)] reg325 = (1'h0);
  reg [(5'h14):(1'h0)] reg839 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg838 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg834 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg832 = (1'h0);
  reg [(5'h15):(1'h0)] reg831 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg830 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg829 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg828 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar826 = (1'h0);
  reg [(5'h12):(1'h0)] forvar823 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg821 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg820 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar817 = (1'h0);
  reg [(5'h13):(1'h0)] reg816 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg815 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg812 = (1'h0);
  reg [(3'h4):(1'h0)] forvar810 = (1'h0);
  reg [(5'h10):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar801 = (1'h0);
  reg [(4'h9):(1'h0)] reg798 = (1'h0);
  reg [(5'h19):(1'h0)] reg797 = (1'h0);
  reg [(5'h11):(1'h0)] reg796 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg795 = (1'h0);
  reg [(4'ha):(1'h0)] reg794 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg792 = (1'h0);
  reg [(4'hb):(1'h0)] forvar790 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg789 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg788 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg787 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg786 = (1'h0);
  reg [(5'h16):(1'h0)] reg785 = (1'h0);
  reg [(2'h2):(1'h0)] reg779 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg780 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar779 = (1'h0);
  reg [(5'h1d):(1'h0)] reg778 = (1'h0);
  reg [(5'h18):(1'h0)] reg777 = (1'h0);
  reg [(4'ha):(1'h0)] reg774 = (1'h0);
  reg [(4'h9):(1'h0)] reg769 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg766 = (1'h0);
  reg [(5'h17):(1'h0)] reg765 = (1'h0);
  reg [(5'h1f):(1'h0)] reg762 = (1'h0);
  reg [(5'h12):(1'h0)] reg761 = (1'h0);
  reg [(5'h19):(1'h0)] forvar760 = (1'h0);
  reg [(4'hb):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg758 = (1'h0);
  reg [(4'hc):(1'h0)] reg755 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg754 = (1'h0);
  reg [(4'hf):(1'h0)] reg753 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar752 = (1'h0);
  reg [(5'h16):(1'h0)] reg751 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg750 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg749 = (1'h0);
  reg [(4'hc):(1'h0)] reg748 = (1'h0);
  reg [(5'h13):(1'h0)] reg747 = (1'h0);
  reg [(2'h3):(1'h0)] reg745 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg744 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg739 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg738 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg736 = (1'h0);
  reg [(5'h11):(1'h0)] reg734 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg733 = (1'h0);
  reg [(5'h1b):(1'h0)] reg732 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar731 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg729 = (1'h0);
  reg [(5'h13):(1'h0)] reg726 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg725 = (1'h0);
  reg [(4'h8):(1'h0)] reg722 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar721 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg720 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar715 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar700 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg717 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg713 = (1'h0);
  reg [(3'h7):(1'h0)] reg712 = (1'h0);
  reg [(3'h5):(1'h0)] reg709 = (1'h0);
  reg [(3'h4):(1'h0)] reg707 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg706 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg704 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg702 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg700 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg698 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg697 = (1'h0);
  reg [(5'h1e):(1'h0)] reg694 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg693 = (1'h0);
  reg [(5'h1c):(1'h0)] reg691 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg690 = (1'h0);
  reg [(5'h1a):(1'h0)] reg689 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg688 = (1'h0);
  reg [(5'h17):(1'h0)] forvar687 = (1'h0);
  reg [(5'h16):(1'h0)] reg685 = (1'h0);
  reg [(5'h19):(1'h0)] reg323 = (1'h0);
  reg [(5'h17):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg318 = (1'h0);
  reg [(3'h7):(1'h0)] reg317 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar316 = (1'h0);
  reg [(3'h5):(1'h0)] forvar302 = (1'h0);
  reg [(4'h8):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar296 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg309 = (1'h0);
  reg [(5'h1f):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg306 = (1'h0);
  reg [(2'h3):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar301 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg300 = (1'h0);
  reg [(5'h1c):(1'h0)] reg298 = (1'h0);
  reg [(5'h1b):(1'h0)] reg297 = (1'h0);
  reg [(5'h1b):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg292 = (1'h0);
  reg [(5'h19):(1'h0)] reg290 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg289 = (1'h0);
  reg [(5'h12):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg286 = (1'h0);
  reg [(3'h4):(1'h0)] forvar285 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg284 = (1'h0);
  reg [(2'h2):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg280 = (1'h0);
  reg [(5'h1d):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg267 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar261 = (1'h0);
  reg [(3'h4):(1'h0)] reg259 = (1'h0);
  reg [(5'h11):(1'h0)] forvar254 = (1'h0);
  reg [(5'h16):(1'h0)] forvar242 = (1'h0);
  reg [(5'h19):(1'h0)] reg265 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar259 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg252 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg250 = (1'h0);
  reg [(5'h1d):(1'h0)] reg249 = (1'h0);
  reg [(4'ha):(1'h0)] reg247 = (1'h0);
  reg [(2'h3):(1'h0)] reg246 = (1'h0);
  reg [(5'h1f):(1'h0)] reg245 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg244 = (1'h0);
  reg [(4'hc):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg242 = (1'h0);
  reg [(4'ha):(1'h0)] reg238 = (1'h0);
  reg [(5'h1d):(1'h0)] reg237 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg236 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg231 = (1'h0);
  reg [(5'h19):(1'h0)] forvar230 = (1'h0);
  reg [(5'h18):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar224 = (1'h0);
  reg [(5'h1e):(1'h0)] reg223 = (1'h0);
  reg [(3'h7):(1'h0)] forvar221 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg220 = (1'h0);
  reg [(5'h12):(1'h0)] reg216 = (1'h0);
  reg [(5'h14):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar212 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg208 = (1'h0);
  reg [(5'h15):(1'h0)] reg207 = (1'h0);
  reg [(5'h1f):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg198 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg197 = (1'h0);
  reg [(3'h5):(1'h0)] reg196 = (1'h0);
  reg [(4'he):(1'h0)] reg193 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg190 = (1'h0);
  reg [(5'h17):(1'h0)] reg189 = (1'h0);
  reg [(4'hb):(1'h0)] reg188 = (1'h0);
  reg [(5'h11):(1'h0)] reg187 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg185 = (1'h0);
  reg [(3'h4):(1'h0)] forvar184 = (1'h0);
  reg [(4'he):(1'h0)] reg183 = (1'h0);
  reg [(4'he):(1'h0)] reg180 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar178 = (1'h0);
  reg [(5'h17):(1'h0)] reg176 = (1'h0);
  reg [(5'h16):(1'h0)] reg174 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar173 = (1'h0);
  reg [(5'h10):(1'h0)] reg172 = (1'h0);
  reg [(5'h19):(1'h0)] reg170 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar166 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg161 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg159 = (1'h0);
  reg [(3'h7):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg156 = (1'h0);
  reg [(5'h1a):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar154 = (1'h0);
  reg [(5'h16):(1'h0)] reg153 = (1'h0);
  reg [(4'ha):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar149 = (1'h0);
  reg [(5'h1c):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg148 = (1'h0);
  reg [(5'h1d):(1'h0)] reg147 = (1'h0);
  reg [(5'h17):(1'h0)] forvar146 = (1'h0);
  reg [(3'h7):(1'h0)] reg144 = (1'h0);
  reg [(3'h6):(1'h0)] reg143 = (1'h0);
  reg [(5'h1e):(1'h0)] reg140 = (1'h0);
  reg [(5'h15):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg138 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg137 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg131 = (1'h0);
  reg [(4'he):(1'h0)] reg128 = (1'h0);
  reg [(4'hf):(1'h0)] forvar127 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg126 = (1'h0);
  reg [(5'h19):(1'h0)] reg124 = (1'h0);
  reg [(5'h1f):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg122 = (1'h0);
  reg [(3'h5):(1'h0)] reg119 = (1'h0);
  reg [(5'h1f):(1'h0)] reg118 = (1'h0);
  reg [(5'h19):(1'h0)] forvar116 = (1'h0);
  reg [(4'hf):(1'h0)] reg99 = (1'h0);
  reg [(5'h18):(1'h0)] forvar98 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg112 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg110 = (1'h0);
  reg [(4'h9):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg106 = (1'h0);
  reg [(5'h1c):(1'h0)] reg105 = (1'h0);
  reg [(4'hb):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg101 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg100 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar99 = (1'h0);
  reg [(4'ha):(1'h0)] reg97 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg96 = (1'h0);
  reg [(3'h5):(1'h0)] reg95 = (1'h0);
  reg [(5'h17):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg93 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg92 = (1'h0);
  reg [(3'h4):(1'h0)] reg91 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg87 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg86 = (1'h0);
  reg [(4'h9):(1'h0)] forvar85 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg82 = (1'h0);
  reg [(5'h18):(1'h0)] forvar81 = (1'h0);
  reg [(5'h10):(1'h0)] forvar80 = (1'h0);
  assign y = {wire842,
                 wire840,
                 wire730,
                 wire683,
                 wire241,
                 wire240,
                 wire164,
                 wire163,
                 wire79,
                 wire78,
                 reg841,
                 reg837,
                 reg836,
                 reg835,
                 reg833,
                 reg827,
                 reg825,
                 reg824,
                 reg822,
                 reg819,
                 reg818,
                 reg814,
                 reg813,
                 reg811,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg803,
                 reg802,
                 reg800,
                 reg799,
                 reg793,
                 reg791,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 reg776,
                 reg775,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 reg768,
                 reg764,
                 reg763,
                 reg757,
                 reg756,
                 reg746,
                 reg743,
                 reg742,
                 reg741,
                 reg740,
                 reg737,
                 reg735,
                 reg728,
                 reg727,
                 reg724,
                 reg723,
                 reg719,
                 reg718,
                 reg716,
                 reg715,
                 reg714,
                 reg711,
                 reg710,
                 reg708,
                 reg705,
                 reg701,
                 reg699,
                 reg687,
                 reg696,
                 reg695,
                 reg692,
                 reg686,
                 reg83,
                 reg89,
                 reg90,
                 reg98,
                 reg102,
                 reg104,
                 reg108,
                 reg111,
                 reg113,
                 reg115,
                 reg117,
                 reg120,
                 reg121,
                 reg125,
                 reg129,
                 reg130,
                 reg132,
                 reg133,
                 reg134,
                 reg135,
                 reg136,
                 reg141,
                 reg142,
                 reg145,
                 reg151,
                 reg152,
                 reg158,
                 reg162,
                 reg165,
                 reg167,
                 reg168,
                 reg169,
                 reg171,
                 reg175,
                 reg177,
                 reg181,
                 reg182,
                 reg186,
                 reg191,
                 reg178,
                 reg194,
                 reg195,
                 reg200,
                 reg201,
                 reg204,
                 reg205,
                 reg206,
                 reg209,
                 reg210,
                 reg213,
                 reg217,
                 reg218,
                 reg219,
                 reg222,
                 reg227,
                 reg228,
                 reg232,
                 reg233,
                 reg234,
                 reg239,
                 reg248,
                 reg251,
                 reg253,
                 reg254,
                 reg255,
                 reg256,
                 reg257,
                 reg258,
                 reg260,
                 reg261,
                 reg262,
                 reg263,
                 reg264,
                 reg266,
                 reg268,
                 reg269,
                 reg270,
                 reg274,
                 reg275,
                 reg276,
                 reg278,
                 reg279,
                 reg281,
                 reg283,
                 reg288,
                 reg291,
                 reg293,
                 reg295,
                 reg296,
                 reg299,
                 reg302,
                 reg304,
                 reg305,
                 reg307,
                 reg310,
                 reg311,
                 reg312,
                 reg313,
                 reg314,
                 reg315,
                 reg320,
                 reg321,
                 reg322,
                 reg324,
                 reg325,
                 reg839,
                 reg838,
                 reg834,
                 reg832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 forvar826,
                 forvar823,
                 reg821,
                 reg820,
                 forvar817,
                 reg816,
                 reg815,
                 reg812,
                 forvar810,
                 reg804,
                 forvar801,
                 reg798,
                 reg797,
                 reg796,
                 reg795,
                 reg794,
                 reg792,
                 forvar790,
                 reg789,
                 reg788,
                 reg787,
                 reg786,
                 reg785,
                 reg779,
                 reg780,
                 forvar779,
                 reg778,
                 reg777,
                 reg774,
                 reg769,
                 reg767,
                 reg766,
                 reg765,
                 reg762,
                 reg761,
                 forvar760,
                 reg759,
                 reg758,
                 reg755,
                 reg754,
                 reg753,
                 forvar752,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg747,
                 reg745,
                 reg744,
                 reg739,
                 reg738,
                 reg736,
                 reg734,
                 reg733,
                 reg732,
                 forvar731,
                 reg729,
                 reg726,
                 reg725,
                 reg722,
                 forvar721,
                 reg720,
                 forvar715,
                 forvar700,
                 reg717,
                 reg713,
                 reg712,
                 reg709,
                 reg707,
                 reg706,
                 reg704,
                 reg703,
                 reg702,
                 reg700,
                 reg698,
                 reg697,
                 reg694,
                 reg693,
                 reg691,
                 reg690,
                 reg689,
                 reg688,
                 forvar687,
                 reg685,
                 reg323,
                 reg319,
                 reg318,
                 reg317,
                 forvar316,
                 forvar302,
                 reg301,
                 forvar296,
                 reg309,
                 reg308,
                 reg306,
                 reg303,
                 forvar301,
                 reg300,
                 reg298,
                 reg297,
                 reg294,
                 reg292,
                 reg290,
                 reg289,
                 reg287,
                 reg286,
                 forvar285,
                 reg284,
                 reg282,
                 reg280,
                 reg277,
                 reg273,
                 reg272,
                 reg271,
                 reg267,
                 forvar261,
                 reg259,
                 forvar254,
                 forvar242,
                 reg265,
                 forvar259,
                 reg252,
                 reg250,
                 reg249,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg231,
                 forvar230,
                 reg229,
                 reg226,
                 reg225,
                 forvar224,
                 reg223,
                 forvar221,
                 reg220,
                 reg216,
                 reg215,
                 reg214,
                 forvar212,
                 reg211,
                 reg208,
                 reg207,
                 reg203,
                 reg202,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg193,
                 reg192,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg185,
                 forvar184,
                 reg183,
                 reg180,
                 reg179,
                 forvar178,
                 reg176,
                 reg174,
                 forvar173,
                 reg172,
                 reg170,
                 forvar166,
                 reg161,
                 reg160,
                 reg159,
                 reg157,
                 reg156,
                 reg155,
                 forvar154,
                 reg153,
                 reg150,
                 forvar149,
                 reg146,
                 reg148,
                 reg147,
                 forvar146,
                 reg144,
                 reg143,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg131,
                 reg128,
                 forvar127,
                 reg126,
                 reg124,
                 reg123,
                 reg122,
                 reg119,
                 reg118,
                 forvar116,
                 reg99,
                 forvar98,
                 reg114,
                 reg112,
                 reg110,
                 reg109,
                 reg107,
                 reg106,
                 reg105,
                 reg103,
                 reg101,
                 reg100,
                 forvar99,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg88,
                 reg87,
                 reg86,
                 forvar85,
                 reg84,
                 reg82,
                 forvar81,
                 forvar80,
                 (1'h0)};
  assign wire78 = ({$signed($signed((wire74 >= (8'hab)))),
                      $signed($unsigned(wire72[(4'hf):(4'ha)]))} < wire76[(2'h2):(2'h2)]);
  assign wire79 = (wire78 ?
                      (wire77[(3'h4):(2'h3)] ?
                          (((wire78 ? wire74 : wire78) ?
                              $signed(wire72) : $unsigned(wire76)) ^~ (wire75[(3'h5):(1'h1)] - (wire72 ?
                              wire72 : wire77))) : (wire74[(3'h4):(2'h3)] ?
                              ({wire73,
                                  wire72} & ((8'hb5) + wire77)) : wire75)) : wire72[(5'h10):(3'h6)]);
  always
    @(posedge clk) begin
      for (forvar80 = (1'h0); (forvar80 < (2'h3)); forvar80 = (forvar80 + (1'h1)))
        begin
          for (forvar81 = (1'h0); (forvar81 < (1'h1)); forvar81 = (forvar81 + (1'h1)))
            begin
              reg82 = (($signed($unsigned(wire78)) ?
                  (~|{(wire75 ?
                          wire78 : wire74)}) : (((~^wire75) || wire79) >= ((^~wire78) ?
                      wire79 : wire72))) >> {$signed($signed((wire72 << wire78)))});
              reg83 <= ((7'h56) > ($unsigned($signed(forvar81[(3'h5):(2'h2)])) ?
                  forvar80[(3'h7):(3'h5)] : wire78));
            end
          reg84 = ($signed((wire77 <= wire76)) ?
              (7'h58) : $unsigned($unsigned($signed(reg83[(1'h0):(1'h0)]))));
          for (forvar85 = (1'h0); (forvar85 < (3'h5)); forvar85 = (forvar85 + (1'h1)))
            begin
              reg86 = $unsigned((reg82[(4'hc):(2'h3)] < {{(forvar85 && forvar80),
                      wire78[(4'h9):(3'h5)]}}));
              reg87 = $signed(($unsigned(wire73[(1'h0):(1'h0)]) ^~ ($unsigned(reg83[(5'h14):(4'h8)]) >>> {wire72[(3'h7):(3'h5)],
                  (wire77 ? forvar85 : (7'h4e))})));
              reg88 = (($signed((&(forvar85 ?
                  wire76 : (7'h53)))) ~^ $signed($signed($unsigned(wire73)))) & reg84[(4'hb):(3'h6)]);
              reg89 <= $signed(wire78);
              reg90 <= $unsigned({$signed($unsigned(reg87))});
              reg91 = $signed((((((7'h48) - wire77) - (wire78 ?
                      wire75 : (8'ha7))) > (8'hbd)) ?
                  reg89 : $signed(wire79)));
            end
          reg92 = (wire72[(3'h6):(3'h6)] ?
              $signed(reg84) : wire72[(4'he):(1'h1)]);
          reg93 = reg87[(3'h6):(3'h5)];
          reg94 = $signed($signed((!((wire76 ? reg92 : reg84) ?
              wire73 : (-wire76)))));
          reg95 = (-$signed($unsigned($unsigned((wire72 > wire78)))));
        end
      reg96 = {($unsigned($signed((reg86 ?
              wire74 : reg95))) < {wire74[(3'h4):(1'h0)],
              (-(wire75 ~^ reg84)),
              ((reg90 << reg84) ? reg93[(3'h5):(3'h5)] : $signed(wire72))}),
          wire79[(3'h7):(3'h7)]};
      reg97 = $signed($unsigned($signed((|(reg82 ? (7'h41) : wire76)))));
      if ((8'hab))
        begin
          reg98 <= (~&($unsigned($unsigned((reg90 - reg91))) == {($unsigned(reg88) || (forvar80 > wire76)),
              $unsigned((|wire72)),
              reg83}));
          for (forvar99 = (1'h0); (forvar99 < (1'h0)); forvar99 = (forvar99 + (1'h1)))
            begin
              reg100 = (~&($signed(reg94[(4'hd):(3'h4)]) ?
                  $unsigned(reg89) : {$signed((&reg87)),
                      $unsigned((~|wire79))}));
              reg101 = (^~{(reg84[(5'h12):(3'h6)] ?
                      $unsigned(forvar80) : wire73),
                  (($unsigned(reg95) ? reg90[(2'h3):(2'h3)] : reg87) ?
                      (~&reg86) : (!wire77))});
              reg102 <= forvar99;
              reg103 = (&{((reg87[(3'h7):(3'h5)] ? reg92 : (wire72 >= reg86)) ?
                      wire78[(3'h5):(1'h0)] : ($signed(reg97) ?
                          $unsigned(forvar80) : reg88[(4'h8):(2'h3)])),
                  forvar81[(5'h10):(5'h10)],
                  (~&($unsigned(wire73) ? (|reg90) : reg93[(3'h5):(2'h3)]))});
              reg104 <= reg103;
              reg105 = ((&$signed($signed(((8'ha7) >= reg102)))) || ($signed($signed((forvar99 > reg83))) ?
                  ((~|reg82) <= (^~$unsigned(forvar81))) : (-$signed((7'h49)))));
            end
          reg106 = (forvar85[(3'h6):(1'h0)] ?
              ((((reg87 ? reg105 : reg93) ?
                  $unsigned((8'h9d)) : $unsigned(forvar85)) & reg93[(5'h12):(4'he)]) || (wire72[(3'h6):(2'h2)] || (reg105[(5'h15):(4'hc)] ^ (^~reg98)))) : ($unsigned((reg96[(3'h5):(1'h1)] ?
                      (wire73 - reg87) : (-wire77))) ?
                  $unsigned(reg104) : $signed(((~&reg83) ?
                      ((8'hbb) ? wire78 : reg87) : ((8'h9f) ?
                          wire79 : reg90)))));
          if ({(^~wire76), reg100[(1'h1):(1'h0)]})
            begin
              reg107 = {{$unsigned($signed($signed(forvar81))), (8'hbc)}};
              reg108 <= $signed(reg107);
              reg109 = reg105;
              reg110 = (~|reg109[(2'h3):(1'h1)]);
              reg111 <= $unsigned(reg106);
            end
          else
            begin
              reg107 = (~&(~^wire77));
              reg108 <= (($signed((reg106[(3'h7):(1'h1)] ^ wire77)) ^ $signed(reg87[(4'ha):(3'h5)])) ^~ $signed((reg96[(4'hb):(4'ha)] == reg82[(3'h7):(3'h4)])));
              reg109 = reg104[(3'h7):(3'h5)];
              reg111 <= $signed($unsigned(wire79));
              reg112 = reg86;
              reg113 <= forvar99[(1'h1):(1'h0)];
              reg114 = reg101;
            end
          reg115 <= $unsigned($unsigned($signed(({reg87,
              (7'h47)} | (|reg102)))));
        end
      else
        begin
          for (forvar98 = (1'h0); (forvar98 < (3'h4)); forvar98 = (forvar98 + (1'h1)))
            begin
              reg99 = forvar80;
              reg100 = ((reg86 && $signed((reg105[(4'h8):(1'h1)] ?
                  (!wire78) : {(8'hac),
                      wire74,
                      reg95}))) >>> $unsigned({$signed((^~reg112)),
                  (~reg114),
                  $unsigned((+(8'hb3)))}));
              reg102 <= reg114[(4'hf):(3'h5)];
              reg103 = (forvar80 ^ $unsigned(wire75[(4'hd):(4'hc)]));
              reg104 <= $signed(forvar85[(1'h0):(1'h0)]);
            end
          reg108 <= $unsigned(reg87);
        end
      for (forvar116 = (1'h0); (forvar116 < (2'h3)); forvar116 = (forvar116 + (1'h1)))
        begin
          if ($signed(reg108))
            begin
              reg117 <= (+(|wire76[(1'h1):(1'h0)]));
              reg118 = reg107;
              reg119 = wire76[(2'h2):(2'h2)];
              reg120 <= ((&$unsigned($signed($signed(forvar85)))) + (~wire73));
              reg121 <= $unsigned($unsigned($unsigned($unsigned((8'hae)))));
            end
          else
            begin
              reg118 = {(($signed($signed(reg87)) ?
                      ($signed(wire77) ?
                          (~^wire72) : reg90) : ($unsigned((7'h57)) ?
                          reg88 : $signed(reg117))) >> {wire72[(5'h11):(4'h9)]}),
                  (^~({(reg101 ? (8'hac) : forvar99),
                      (reg91 + forvar98)} << $unsigned((~&reg109)))),
                  (reg94[(5'h11):(2'h3)] ?
                      ((reg83[(5'h19):(2'h2)] >>> (8'hb8)) && reg100[(3'h7):(3'h6)]) : (+(reg109 ?
                          $unsigned(reg120) : {reg94, reg109})))};
              reg119 = reg98[(4'ha):(4'ha)];
              reg122 = (reg83 ?
                  (8'hb4) : $signed($unsigned($unsigned((reg91 ?
                      (7'h52) : reg87)))));
              reg123 = reg96;
            end
          if ((reg117 ? (&reg92) : $signed(reg87[(4'hd):(4'hb)])))
            begin
              reg124 = {reg89[(5'h10):(3'h7)]};
              reg125 <= ((reg94 >>> ((-wire78) < ($unsigned(reg96) <= reg105[(5'h1a):(3'h7)]))) <= (8'h9d));
              reg126 = $signed((^~(8'haa)));
            end
          else
            begin
              reg124 = wire79[(2'h3):(1'h0)];
            end
        end
      for (forvar127 = (1'h0); (forvar127 < (1'h0)); forvar127 = (forvar127 + (1'h1)))
        begin
          if (($signed($unsigned(wire73)) ?
              $signed(forvar99) : $signed($unsigned($unsigned((wire79 ?
                  reg113 : reg124))))))
            begin
              reg128 = reg121[(2'h2):(2'h2)];
              reg129 <= $unsigned(((+{$signed(reg119)}) <<< reg117[(5'h10):(4'h9)]));
              reg130 <= ($unsigned($signed(($unsigned(reg112) < (&wire79)))) | $unsigned($signed($unsigned($signed((7'h47))))));
              reg131 = reg122[(5'h10):(4'he)];
              reg132 <= reg92;
              reg133 <= wire74;
            end
          else
            begin
              reg128 = $unsigned((8'hb0));
              reg129 <= $unsigned({$signed((reg130[(3'h4):(3'h4)] - reg121[(5'h16):(2'h2)])),
                  $signed((wire79 | $unsigned(forvar116)))});
              reg131 = ((~reg92) ?
                  ((($signed((8'hac)) & (reg92 + reg86)) ?
                      ($unsigned((8'had)) ?
                          ((7'h4a) << reg120) : $unsigned(reg119)) : $unsigned((wire77 || reg120))) > $signed(reg88)) : reg125);
              reg132 <= (~|reg126);
              reg133 <= $signed(reg109);
            end
          reg134 <= {(wire72 ?
                  ({$unsigned(reg83),
                      reg91[(2'h2):(1'h0)]} - $signed((reg91 <<< reg96))) : (reg112[(2'h3):(2'h3)] ?
                      (reg93 ? $unsigned(reg87) : (~^reg113)) : forvar99))};
          reg135 <= ($unsigned($signed((wire77[(4'he):(4'he)] > reg100))) + reg112[(4'hf):(4'hc)]);
          if (($unsigned((($signed((7'h54)) >>> $unsigned(reg133)) > reg130)) ?
              {(^~($unsigned(reg97) ?
                      $unsigned((7'h47)) : (-reg89)))} : ((reg110[(1'h1):(1'h0)] ?
                      (~&(^~forvar98)) : ($signed(reg101) | $signed((8'h9e)))) ?
                  ((~&(^reg120)) ?
                      $signed(reg99[(2'h3):(1'h0)]) : {$signed(reg89)}) : ($signed(reg119[(3'h5):(2'h3)]) < $signed($unsigned(reg104))))))
            begin
              reg136 <= (($signed((reg113[(5'h13):(3'h4)] ?
                  wire79[(1'h0):(1'h0)] : $signed(reg92))) & {reg108,
                  (reg130[(3'h5):(2'h3)] ?
                      (wire75 ? reg131 : reg115) : (forvar80 ?
                          forvar116 : forvar85)),
                  $signed($unsigned(wire76))}) || $signed(wire77[(1'h0):(1'h0)]));
              reg137 = reg136[(2'h3):(2'h3)];
              reg138 = (((7'h42) ?
                  (($signed(reg130) ?
                      {reg109} : reg107) >= (&(reg132 * reg95))) : (reg129 - {reg102[(3'h6):(2'h2)]})) * reg108[(4'ha):(1'h0)]);
              reg139 = wire75;
              reg140 = ($signed((reg114 - (reg89 ?
                      $signed(reg110) : reg89[(4'he):(4'ha)]))) ?
                  reg93 : (8'hb8));
              reg141 <= reg113[(4'hc):(4'hc)];
            end
          else
            begin
              reg137 = $signed((~(-forvar98[(5'h15):(5'h15)])));
              reg138 = reg129;
              reg139 = ((~&(reg83[(4'hc):(3'h4)] & wire79)) ?
                  reg104 : reg119[(1'h0):(1'h0)]);
              reg141 <= $unsigned($unsigned(reg100));
              reg142 <= $signed(((~$unsigned((reg90 | (7'h47)))) < (reg89[(2'h3):(1'h1)] ~^ (^(reg126 ?
                  reg95 : (8'hb1))))));
              reg143 = {reg96[(2'h3):(1'h0)]};
              reg144 = ($signed(wire75[(3'h4):(1'h0)]) ^ ((reg97[(3'h5):(3'h5)] <= reg107[(5'h10):(4'h8)]) ?
                  $signed(($unsigned(reg123) ?
                      $signed(reg121) : (reg135 == (8'hbd)))) : $unsigned($unsigned($signed((8'ha9))))));
            end
        end
      reg145 <= (~$signed((wire76 <= ($signed((7'h57)) <<< $signed(reg123)))));
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned({(8'hae)})))
        begin
          for (forvar146 = (1'h0); (forvar146 < (3'h4)); forvar146 = (forvar146 + (1'h1)))
            begin
              reg147 = $unsigned({(7'h46)});
            end
          reg148 = $signed(reg136);
        end
      else
        begin
          reg146 = $unsigned((|(($signed(reg145) ?
                  (+reg108) : $unsigned(wire73)) ?
              (~^reg145[(3'h5):(1'h0)]) : $unsigned((reg133 >= wire73)))));
        end
      for (forvar149 = (1'h0); (forvar149 < (1'h0)); forvar149 = (forvar149 + (1'h1)))
        begin
          reg150 = reg142;
          reg151 <= {(|(^~reg132[(4'hb):(1'h0)])),
              $unsigned($unsigned(((|(7'h4f)) ? $unsigned(reg129) : reg148)))};
          reg152 <= forvar146;
          reg153 = reg117[(4'h8):(2'h3)];
        end
      for (forvar154 = (1'h0); (forvar154 < (3'h4)); forvar154 = (forvar154 + (1'h1)))
        begin
          if ((($unsigned(($signed((7'h43)) ? (-reg104) : (^~reg113))) ?
              $unsigned((~&reg141[(2'h2):(1'h1)])) : ((reg133[(5'h15):(4'hd)] < (reg130 ?
                      reg132 : reg120)) ?
                  ((-(8'h9f)) ^~ (+wire76)) : wire72)) < (~^$unsigned(reg148))))
            begin
              reg155 = reg141[(1'h1):(1'h1)];
              reg156 = (wire73 ?
                  {($signed((reg89 ? wire73 : reg98)) ?
                          (^(wire78 | (8'hb2))) : (^~(wire75 != (7'h50))))} : reg125[(5'h1a):(4'hb)]);
              reg157 = reg153[(5'h10):(1'h0)];
            end
          else
            begin
              reg158 <= (+((wire72[(3'h5):(2'h3)] >>> wire72[(3'h7):(3'h6)]) || (({reg111} <<< (8'hb2)) ?
                  $signed(reg89) : reg113[(2'h3):(2'h2)])));
            end
          reg159 = reg111;
        end
      reg160 = $signed($signed(reg102[(5'h18):(4'hc)]));
      reg161 = ($unsigned((8'haf)) || $unsigned((^reg111[(4'hb):(4'h8)])));
      reg162 <= reg125[(2'h2):(1'h1)];
    end
  assign wire163 = $signed(((reg134[(1'h0):(1'h0)] ?
                           ((reg102 ? wire77 : reg120) ^~ (reg121 ?
                               reg120 : reg113)) : $unsigned(wire78)) ?
                       $unsigned(reg158[(2'h3):(2'h3)]) : reg142));
  assign wire164 = wire75;
  always
    @(posedge clk) begin
      reg165 <= (wire78 == (|$signed(wire74[(1'h1):(1'h1)])));
      for (forvar166 = (1'h0); (forvar166 < (1'h1)); forvar166 = (forvar166 + (1'h1)))
        begin
          if ($signed({$unsigned(reg111[(4'hd):(4'h9)]),
              (7'h4d),
              {$signed((wire79 != reg135))}}))
            begin
              reg167 <= ($unsigned((-$unsigned((|(8'hb1))))) ?
                  (|$unsigned((^{reg136, reg113}))) : reg133[(4'hb):(3'h5)]);
            end
          else
            begin
              reg167 <= (!$unsigned(reg108));
              reg168 <= (|$signed((|$signed((reg132 ? (7'h44) : reg129)))));
              reg169 <= (wire73 * ($unsigned($unsigned(wire73)) ?
                  (wire77[(5'h10):(4'hf)] == $unsigned((7'h4e))) : {(reg113[(5'h1b):(5'h14)] ?
                          {wire164, reg117, (8'ha0)} : {wire72, reg136})}));
              reg170 = $signed($signed(wire163[(4'h8):(3'h6)]));
            end
          reg171 <= {(wire163 ?
                  {reg115[(4'h9):(1'h0)],
                      wire76[(2'h2):(1'h0)],
                      ((&reg151) - ((8'h9f) >>> reg134))} : reg135),
              reg98[(4'hc):(3'h7)]};
          reg172 = {(^(^($unsigned(reg102) ? reg133 : $signed(reg83)))),
              wire75[(4'hd):(3'h4)]};
          for (forvar173 = (1'h0); (forvar173 < (1'h1)); forvar173 = (forvar173 + (1'h1)))
            begin
              reg174 = (reg145[(4'hb):(1'h0)] < {$unsigned(reg120[(3'h7):(3'h5)]),
                  reg132[(3'h4):(3'h4)]});
            end
          if ({(~&$signed(((reg174 ^~ wire77) ?
                  reg132 : reg134[(3'h5):(2'h3)]))),
              ($signed({$signed((8'haa))}) ?
                  reg136 : $signed((!(reg111 && reg174)))),
              wire76})
            begin
              reg175 <= (($unsigned($signed(reg132[(3'h6):(3'h4)])) >>> ($signed(wire163[(1'h1):(1'h1)]) ?
                  $unsigned(wire79[(3'h5):(2'h2)]) : $signed((!(8'ha2))))) >> reg111[(5'h13):(5'h10)]);
              reg176 = $unsigned(reg162);
              reg177 <= (($unsigned(reg132[(4'h8):(2'h2)]) - $signed(((&wire72) ?
                  (reg171 <<< reg169) : (reg174 || reg111)))) != (~|reg121[(4'h8):(2'h3)]));
            end
          else
            begin
              reg175 <= reg176[(4'hf):(3'h7)];
              reg176 = $signed(reg142[(3'h7):(3'h4)]);
            end
        end
      if ($signed((~^reg158[(4'hd):(1'h0)])))
        begin
          for (forvar178 = (1'h0); (forvar178 < (1'h1)); forvar178 = (forvar178 + (1'h1)))
            begin
              reg179 = ((7'h51) || reg169[(4'h8):(4'h8)]);
            end
          reg180 = $signed({$unsigned($unsigned((reg170 ? reg83 : reg158))),
              {(+reg158[(4'hd):(2'h2)])},
              ($signed($unsigned(reg111)) ?
                  $unsigned(reg111) : $unsigned($unsigned(reg136)))});
          if ((~|reg145))
            begin
              reg181 <= reg168[(3'h4):(2'h3)];
              reg182 <= ((~$unsigned($unsigned((|reg165)))) ?
                  (7'h55) : $signed((reg102 ? {(8'hbb)} : reg120)));
            end
          else
            begin
              reg183 = $unsigned((&(|(7'h46))));
            end
          for (forvar184 = (1'h0); (forvar184 < (1'h0)); forvar184 = (forvar184 + (1'h1)))
            begin
              reg185 = $unsigned($signed((reg168 < $signed($unsigned(reg176)))));
              reg186 <= {((!(~&$unsigned(reg117))) ?
                      $unsigned((~(8'hbc))) : $unsigned(wire77)),
                  (^~reg89)};
            end
          if (wire73)
            begin
              reg187 = ($signed({$signed((^~reg120))}) ?
                  $signed(wire73[(2'h3):(1'h0)]) : (7'h4d));
              reg188 = (~{{$unsigned((^reg145)), (^(^forvar173)), (8'hab)},
                  $signed((forvar178 ? wire163[(4'he):(4'he)] : (+(8'hbc)))),
                  $unsigned(($unsigned((7'h44)) && (|reg142)))});
              reg189 = $signed((($unsigned($unsigned((7'h45))) ~^ $unsigned((reg129 ~^ (7'h4f)))) <<< $signed({$signed(reg111),
                  (reg174 ? wire75 : reg142),
                  wire74[(2'h3):(1'h0)]})));
              reg190 = $signed($unsigned(({$unsigned(reg169)} ^ {reg141,
                  (wire74 ? reg83 : reg170),
                  $signed(reg189)})));
              reg191 <= ((({(wire73 ? forvar178 : wire73), $unsigned((8'hac))} ?
                      (reg167 <= (wire74 ? reg190 : reg167)) : $signed((reg167 ?
                          wire72 : reg158))) ?
                  ($unsigned($signed(wire73)) ?
                      ({reg104, reg186} ?
                          $unsigned((7'h47)) : ((8'hb6) * (7'h53))) : reg83) : $signed((((7'h50) ~^ reg174) >>> (+reg89)))) <= (~|$signed((reg174[(3'h6):(1'h0)] ^~ (+reg132)))));
            end
          else
            begin
              reg191 <= ((-reg90[(4'h9):(4'h8)]) ?
                  reg90 : ((^((reg111 ? reg167 : reg188) ?
                      (reg129 == reg190) : reg90[(4'hd):(4'ha)])) ~^ $unsigned(((reg181 || reg170) >>> (7'h48)))));
            end
        end
      else
        begin
          reg178 <= (+((^$unsigned(reg136[(1'h0):(1'h0)])) && $unsigned($unsigned(reg179))));
          reg179 = {(~^$unsigned((reg182[(5'h10):(4'hf)] >= reg179[(2'h3):(2'h2)]))),
              $unsigned({(reg141 != {reg130})}),
              $unsigned($unsigned(reg188[(4'hb):(2'h2)]))};
        end
      if (((&(((&forvar173) != forvar178[(5'h12):(3'h7)]) > ($unsigned(reg121) ?
          reg135[(4'ha):(2'h3)] : (reg151 ? reg186 : forvar184)))) <<< wire74))
        begin
          if (reg176[(4'he):(4'hb)])
            begin
              reg192 = $signed(((reg134[(4'h9):(3'h6)] ?
                  wire73 : $unsigned((reg176 - reg142))) >>> ($signed((reg121 ~^ (7'h4a))) ~^ reg179)));
              reg193 = (({$signed((wire79 - reg135)),
                  $signed(wire75)} - reg135[(4'he):(4'ha)]) != (reg165[(3'h6):(3'h6)] << {$signed({reg171,
                      reg141})}));
              reg194 <= reg133;
              reg195 <= $signed(reg186);
              reg196 = reg132[(4'h8):(2'h2)];
            end
          else
            begin
              reg192 = {reg165, forvar178, forvar184[(2'h2):(2'h2)]};
              reg193 = $unsigned(reg189);
              reg194 <= reg104;
            end
          reg197 = (|((~reg170[(5'h15):(4'hb)]) ?
              wire72 : $unsigned(reg176[(5'h12):(2'h2)])));
          if ((^~$signed((|((reg188 ? (8'hbc) : reg196) ?
              forvar166 : $signed(reg189))))))
            begin
              reg198 = $unsigned({(8'h9e),
                  $signed(((~^reg183) ?
                      (reg194 ? reg180 : (8'hb9)) : $unsigned(reg178))),
                  $unsigned((forvar173[(1'h1):(1'h0)] ?
                      reg134 : $unsigned(wire73)))});
              reg199 = reg104[(4'h8):(1'h1)];
              reg200 <= $unsigned({reg196[(3'h4):(3'h4)], $signed(reg121)});
              reg201 <= reg167;
              reg202 = (^~((((~&(8'ha4)) <= $signed(reg152)) ?
                      reg200 : $unsigned(reg113)) ?
                  ($unsigned((reg189 > reg130)) <<< (~|(&reg188))) : reg167[(4'h9):(3'h6)]));
              reg203 = ($signed($signed(reg177)) & wire74);
              reg204 <= (~|$signed(((~&(+reg203)) && $signed(wire74))));
            end
          else
            begin
              reg200 <= ((!reg193) ?
                  (^~reg129) : (reg102[(5'h12):(4'ha)] <= $unsigned({(reg129 ?
                          reg121 : (8'hba)),
                      wire75})));
              reg201 <= {{(reg168 <<< reg90),
                      $unsigned(forvar173),
                      (~^(|(reg108 ? wire77 : reg129)))},
                  reg176,
                  (+$unsigned($unsigned({reg113})))};
              reg202 = (-$unsigned(((^~(^~reg121)) ?
                  (|(forvar173 ?
                      reg134 : reg108)) : ($unsigned(wire75) ~^ ((7'h57) ?
                      reg172 : wire79)))));
              reg203 = $signed(reg182[(4'ha):(3'h4)]);
              reg204 <= {$signed($signed($signed((reg175 ?
                      (8'ha6) : forvar166)))),
                  $signed((reg170[(5'h15):(5'h14)] ^~ (~&$signed(reg111)))),
                  forvar173};
              reg205 <= (~^(~($unsigned((reg177 ? reg191 : reg200)) & reg108)));
              reg206 <= reg204;
            end
          if (($signed($unsigned({(reg117 >>> wire77),
              (^~reg199),
              $signed(reg203)})) ^~ (~|(reg201[(2'h2):(2'h2)] ?
              (8'h9f) : {reg197, reg179, $unsigned(reg169)}))))
            begin
              reg207 = (7'h48);
            end
          else
            begin
              reg207 = ({($unsigned($unsigned(reg194)) >> reg202[(3'h5):(1'h0)]),
                  $unsigned($signed((-wire75))),
                  reg202[(3'h6):(2'h2)]} - {$unsigned((((8'hb4) ?
                          wire79 : reg133) ?
                      $signed(reg205) : (~|reg152))),
                  reg113[(5'h15):(4'h9)],
                  (+(reg169[(5'h12):(5'h12)] == (reg167 << forvar173)))});
              reg208 = (reg125 ?
                  (reg135[(3'h5):(3'h5)] ?
                      $signed(reg186) : ((7'h44) >= {reg125[(4'h9):(1'h0)],
                          reg187[(2'h2):(1'h0)],
                          (8'haa)})) : (+forvar184));
              reg209 <= (reg132 ?
                  $signed($signed(((reg113 >= reg205) ?
                      ((8'hab) >= reg145) : {reg188, (8'hbf)}))) : reg104);
              reg210 <= (!$unsigned($signed(reg167[(4'he):(3'h4)])));
              reg211 = ($signed(($unsigned(reg136[(2'h3):(1'h0)]) ?
                      reg168 : (~|$unsigned(reg108)))) ?
                  {reg204,
                      (reg158[(4'hb):(4'hb)] ?
                          reg129[(2'h3):(2'h2)] : $signed((reg89 != reg168)))} : (~|{(~^reg188),
                      {$signed(reg178),
                          {reg113, reg125, reg205},
                          (wire75 ? (7'h53) : reg89)}}));
            end
          for (forvar212 = (1'h0); (forvar212 < (2'h3)); forvar212 = (forvar212 + (1'h1)))
            begin
              reg213 <= $unsigned(((reg151 ?
                      (wire164[(4'hc):(4'h8)] ?
                          $signed(reg207) : $unsigned((8'ha7))) : ((7'h58) ?
                          $signed(reg125) : reg181[(4'h8):(3'h5)])) ?
                  reg187 : $signed($signed($unsigned(reg172)))));
              reg214 = $unsigned((-((reg120[(3'h4):(1'h0)] << {wire79,
                      wire77}) ?
                  reg206 : (reg208[(3'h4):(1'h0)] ?
                      reg171 : $signed(forvar178)))));
              reg215 = reg132[(4'hb):(1'h0)];
              reg216 = reg120;
              reg217 <= (reg183 ?
                  {$signed($signed($unsigned(reg130))),
                      $unsigned(wire77)} : ((~&((reg198 >= reg130) ?
                          (&reg195) : (forvar184 && reg213))) ?
                      wire78 : $unsigned(({wire75} | (reg132 ?
                          reg135 : reg214)))));
              reg218 <= {(($unsigned($signed(reg162)) ?
                          {wire164,
                              $unsigned(reg145),
                              $unsigned((8'h9d))} : ((|reg187) ?
                              (reg135 ? reg133 : reg206) : (reg194 ?
                                  wire74 : reg168))) ?
                      $signed(((reg175 <= reg201) || reg191)) : ((^~reg205[(1'h1):(1'h1)]) >>> (reg186 ?
                          forvar173[(2'h2):(2'h2)] : wire164)))};
              reg219 <= wire77[(4'hd):(4'hd)];
            end
          reg220 = (forvar212 || reg216[(5'h12):(1'h1)]);
        end
      else
        begin
          reg192 = (reg187 ?
              $signed((~((-reg172) <= reg198))) : (+{$signed(reg168)}));
          if ((^~((~|$signed($unsigned(reg158))) ?
              reg205[(5'h12):(4'h8)] : $unsigned(reg201[(1'h1):(1'h1)]))))
            begin
              reg194 <= $signed(((reg179 ?
                  $unsigned($signed(reg108)) : (8'hbd)) - ((reg208[(3'h7):(3'h4)] ?
                      reg151[(3'h6):(2'h3)] : (reg193 ? reg204 : reg129)) ?
                  (8'h9d) : reg201[(1'h1):(1'h0)])));
              reg196 = ($unsigned($signed(reg121[(4'hd):(3'h5)])) ^~ $unsigned((($unsigned(forvar178) == (reg214 ?
                      reg130 : reg120)) ?
                  (!(-reg197)) : (~^(reg209 ? reg152 : reg170)))));
              reg197 = reg199;
              reg200 <= reg113;
            end
          else
            begin
              reg194 <= (($unsigned($signed(reg218[(4'hb):(3'h6)])) ~^ ($signed((reg136 ?
                          reg151 : reg213)) ?
                      reg187 : reg136[(2'h3):(2'h2)])) ?
                  $unsigned((($signed((8'ha9)) == (reg195 != reg186)) ?
                      $signed((forvar184 ?
                          reg218 : reg182)) : reg181)) : forvar166[(2'h2):(2'h2)]);
              reg196 = reg195[(3'h6):(1'h1)];
              reg197 = ($signed((8'hbd)) ?
                  reg171 : (wire79 ?
                      ($signed(reg115[(1'h0):(1'h0)]) ?
                          ({reg198, reg134, reg201} ?
                              wire72[(4'h8):(3'h7)] : $unsigned(reg136)) : reg181[(5'h1c):(4'hc)]) : $unsigned(({reg174,
                              reg121} ?
                          (|reg209) : {wire164}))));
              reg200 <= reg200[(4'h8):(2'h2)];
            end
        end
      for (forvar221 = (1'h0); (forvar221 < (3'h5)); forvar221 = (forvar221 + (1'h1)))
        begin
          reg222 <= $unsigned($unsigned({$signed(wire72[(4'hf):(4'hf)]),
              (~|(reg174 * reg215))}));
          reg223 = reg129[(5'h12):(5'h12)];
          for (forvar224 = (1'h0); (forvar224 < (2'h3)); forvar224 = (forvar224 + (1'h1)))
            begin
              reg225 = $signed(($signed((~&reg136[(1'h0):(1'h0)])) ?
                  $unsigned($signed($signed((7'h4e)))) : $signed((~|$signed(reg133)))));
              reg226 = (!(~|{{(reg198 ? reg113 : (8'hac)),
                      reg198[(4'h9):(4'h8)],
                      reg172},
                  reg102}));
              reg227 <= $unsigned($signed(wire73));
              reg228 <= $unsigned($signed((reg219[(5'h14):(2'h2)] ?
                  ((forvar212 ?
                      reg102 : reg171) - (wire164 | reg195)) : {reg172,
                      (reg134 < reg125),
                      ((7'h54) <<< (8'haa))})));
              reg229 = {{reg162[(2'h2):(1'h1)],
                      reg142[(2'h3):(1'h1)],
                      $unsigned((~|reg216))}};
            end
          for (forvar230 = (1'h0); (forvar230 < (1'h1)); forvar230 = (forvar230 + (1'h1)))
            begin
              reg231 = ((^~(~|{(~|wire78)})) < reg210[(3'h7):(2'h2)]);
              reg232 <= {(7'h4b),
                  $unsigned((&$unsigned((reg168 * reg220)))),
                  {{reg219[(5'h15):(2'h3)]},
                      $signed($signed($unsigned(reg168))),
                      ($signed($signed(wire73)) ?
                          reg113 : (~^$signed(reg171)))}};
              reg233 <= $signed((7'h40));
            end
          reg234 <= (^reg203);
          reg235 = $unsigned($unsigned((~^reg145[(3'h6):(2'h2)])));
        end
      reg236 = (^(reg151 ?
          (reg199 ?
              $unsigned($unsigned(reg223)) : forvar178[(5'h19):(4'h8)]) : (-(reg227[(2'h2):(2'h2)] ?
              (^reg215) : {reg198, (8'haf), reg165}))));
      reg237 = reg187[(4'h9):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg238 = (+$unsigned($signed((+((7'h4d) ? (8'hba) : reg125)))));
      reg239 <= $signed((8'had));
    end
  assign wire240 = $signed((|wire163));
  assign wire241 = reg201[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      if (reg234[(2'h2):(2'h2)])
        begin
          if ($unsigned(reg217))
            begin
              reg242 = (wire164[(4'h9):(2'h3)] <= (^reg129));
              reg243 = reg129[(1'h0):(1'h0)];
              reg244 = reg233;
              reg245 = ((~&$unsigned(((+(8'hbd)) <= {reg98,
                  reg178}))) >>> wire72);
              reg246 = {($unsigned((!reg142)) ?
                      (reg177[(5'h1d):(4'hb)] << (~&(wire241 * reg244))) : ({(reg142 > (7'h46)),
                          (reg162 >> wire76)} | $signed($unsigned(reg209))))};
              reg247 = {($unsigned((^{reg134})) <<< (reg133 ?
                      $signed((reg111 <<< reg228)) : reg243)),
                  ($signed(reg186[(4'hc):(3'h5)]) ?
                      (~^(~&(reg201 ?
                          reg244 : (7'h40)))) : (-$signed(reg218[(4'h9):(1'h0)]))),
                  (^~$signed((reg191[(3'h5):(3'h4)] == $unsigned(reg132))))};
            end
          else
            begin
              reg242 = {reg111};
              reg243 = (~($unsigned(($unsigned(reg113) ^ $unsigned(reg239))) ?
                  ($signed((reg113 ? reg141 : reg228)) ?
                      $unsigned(reg111[(3'h6):(1'h0)]) : (^{(8'hbf),
                          (8'hb1),
                          (7'h52)})) : (((+reg217) <= reg135) ?
                      {$unsigned(reg195)} : $unsigned((~reg210)))));
              reg248 <= (reg115 ?
                  (reg142 ?
                      {(8'hbc)} : (reg168 ?
                          ((reg178 ?
                              reg233 : (8'ha4)) > (^~(7'h56))) : $signed($signed(reg135)))) : (reg178[(5'h1c):(5'h1a)] ?
                      (|wire164[(3'h6):(1'h1)]) : reg233[(4'hb):(2'h3)]));
              reg249 = $unsigned(reg135[(4'hf):(2'h2)]);
            end
          reg250 = (reg181[(3'h5):(2'h3)] == ((reg83 | reg141[(1'h1):(1'h0)]) ?
              $signed((reg89 == reg171[(3'h4):(2'h3)])) : (((7'h4b) == $unsigned(reg169)) ~^ {reg246[(1'h1):(1'h1)],
                  (reg141 ? reg219 : reg232)})));
          if ($unsigned({reg108}))
            begin
              reg251 <= $signed(reg115);
              reg252 = reg250;
            end
          else
            begin
              reg251 <= (reg194 ?
                  $signed(reg175) : $signed((reg134[(3'h4):(1'h1)] ^ $signed((reg136 ^~ reg227)))));
              reg253 <= (|reg90[(3'h7):(3'h6)]);
              reg254 <= ({$unsigned($signed($unsigned(reg135))), reg222} ?
                  $unsigned($signed(reg239[(4'hc):(3'h4)])) : ($signed((!(reg218 ?
                      wire77 : (7'h53)))) | $signed(reg125[(5'h17):(5'h13)])));
              reg255 <= $unsigned((^reg182));
              reg256 <= reg130[(2'h2):(1'h0)];
            end
          reg257 <= reg205[(3'h4):(3'h4)];
          reg258 <= reg251[(4'hc):(4'hc)];
          for (forvar259 = (1'h0); (forvar259 < (2'h2)); forvar259 = (forvar259 + (1'h1)))
            begin
              reg260 <= $unsigned($unsigned(((~|((8'hab) || (7'h46))) ?
                  $unsigned((reg151 ?
                      wire72 : reg243)) : $unsigned($signed((8'hbc))))));
              reg261 <= $unsigned($unsigned((&reg234)));
              reg262 <= reg201;
              reg263 <= (^~$signed($unsigned(((reg218 ? reg141 : wire75) ?
                  {reg132, reg204, wire241} : $signed(wire72)))));
              reg264 <= (7'h54);
              reg265 = reg258;
              reg266 <= $unsigned($signed(reg165));
            end
        end
      else
        begin
          for (forvar242 = (1'h0); (forvar242 < (2'h2)); forvar242 = (forvar242 + (1'h1)))
            begin
              reg243 = (reg121 ?
                  $unsigned(reg201[(1'h0):(1'h0)]) : (-$signed($unsigned((reg266 & forvar242)))));
              reg248 <= (((^{$unsigned(reg169),
                      ((8'ha4) & reg251),
                      (!(8'hb4))}) && $signed(reg249)) ?
                  $signed($unsigned({{(7'h55), (7'h55)},
                      (~&reg222)})) : (!$signed((reg222[(3'h5):(3'h4)] ?
                      wire164 : reg135))));
              reg249 = ((reg133[(5'h12):(5'h11)] ?
                  $signed($unsigned($unsigned(reg253))) : reg132) || $signed((reg158[(5'h12):(3'h5)] ?
                  {(~&reg244), {reg257, reg261, (7'h44)}} : reg204)));
              reg251 <= (reg245 ?
                  {wire79,
                      {wire76[(2'h2):(1'h1)], reg218}} : {($unsigned(reg151) ?
                          reg108[(3'h7):(2'h2)] : $unsigned({reg175,
                              (8'ha4)}))});
              reg252 = $unsigned(reg233[(2'h2):(2'h2)]);
              reg253 <= ($unsigned((reg254[(5'h15):(5'h14)] || (reg117 ~^ (~|reg158)))) <= ((reg246[(1'h1):(1'h1)] ?
                      $signed((reg255 ?
                          reg178 : reg194)) : wire77[(4'hf):(4'ha)]) ?
                  (~(reg194 ?
                      reg205[(2'h3):(2'h2)] : {(8'hab),
                          wire240})) : $unsigned((reg129 ?
                      reg152[(2'h3):(1'h0)] : {(7'h49), reg125}))));
            end
          for (forvar254 = (1'h0); (forvar254 < (3'h4)); forvar254 = (forvar254 + (1'h1)))
            begin
              reg259 = (reg142 | (^(8'ha1)));
              reg260 <= {$unsigned($signed(($signed((8'h9d)) <<< (reg108 ?
                      reg175 : wire74))))};
            end
          for (forvar261 = (1'h0); (forvar261 < (3'h4)); forvar261 = (forvar261 + (1'h1)))
            begin
              reg265 = reg135[(4'hc):(1'h0)];
            end
        end
      if (($unsigned($signed({(&reg254), reg258, (~reg89)})) <<< reg178))
        begin
          reg267 = reg113;
          if ((reg260 & $unsigned((^~(((7'h56) * reg246) && (reg242 && forvar261))))))
            begin
              reg268 <= ((reg162 ?
                  $unsigned(((reg260 ? reg205 : reg228) ?
                      {reg186} : $unsigned(reg152))) : ({$unsigned(reg181),
                      reg133} - $unsigned($signed((7'h58))))) ^~ ((reg219[(4'ha):(1'h0)] > $unsigned($unsigned(reg251))) + (reg250 ^~ $unsigned(((7'h4d) >= reg113)))));
              reg269 <= (-($signed((~&(7'h43))) ?
                  reg206[(4'hf):(2'h3)] : (reg165 ^ $signed(((7'h43) || reg83)))));
              reg270 <= reg132[(3'h6):(1'h0)];
            end
          else
            begin
              reg271 = reg259[(2'h2):(1'h0)];
              reg272 = $signed(reg104);
              reg273 = reg218[(4'hd):(4'h8)];
              reg274 <= $unsigned($signed($unsigned(reg222)));
              reg275 <= ($signed((!((&reg171) && wire76[(1'h0):(1'h0)]))) << (((^~$unsigned(reg265)) ?
                  (((8'ha8) ?
                      reg168 : reg247) != reg111[(4'hb):(4'ha)]) : $signed($signed((7'h49)))) && reg133));
              reg276 <= $signed(reg89[(4'hd):(3'h6)]);
            end
        end
      else
        begin
          if (reg98[(1'h1):(1'h0)])
            begin
              reg268 <= (~|reg244);
              reg269 <= reg115;
              reg270 <= reg275[(2'h3):(1'h0)];
              reg274 <= {reg254,
                  ($signed(reg121) ?
                      wire163[(4'h8):(3'h7)] : (-((reg234 ? reg191 : reg265) ?
                          reg194 : (reg228 & reg246))))};
              reg277 = $signed($unsigned((~|{(7'h40), $signed(reg158)})));
              reg278 <= (reg232 >= reg239);
            end
          else
            begin
              reg268 <= (((^~reg259) ?
                      $unsigned(($signed((8'hba)) + $unsigned(reg255))) : reg141[(1'h0):(1'h0)]) ?
                  (^~reg219[(3'h6):(2'h3)]) : (~|(((!reg272) ?
                          reg246[(1'h1):(1'h0)] : $signed(reg125)) ?
                      {$unsigned(reg165), $unsigned(reg234)} : ({(8'haa)} ?
                          ((7'h45) ? reg263 : reg209) : $unsigned(reg269)))));
              reg269 <= reg210[(2'h3):(2'h3)];
              reg271 = $signed(reg243[(3'h4):(2'h3)]);
              reg272 = forvar259;
              reg274 <= reg243[(4'ha):(2'h2)];
              reg275 <= (|($unsigned(($signed(reg186) ^ (reg260 ?
                  reg273 : reg115))) && $unsigned(($signed(reg243) >= reg130[(3'h7):(3'h7)]))));
            end
          if (($unsigned({$unsigned((reg259 - reg117)),
                  wire73[(2'h2):(1'h1)]}) ?
              (^$signed(reg261[(4'he):(3'h7)])) : (((~^(reg204 * reg275)) << (~^reg249)) ?
                  ($unsigned($signed(reg178)) && $unsigned($signed(reg177))) : reg213)))
            begin
              reg279 <= (8'hb9);
              reg280 = $unsigned({reg169,
                  (-$signed($unsigned(reg253))),
                  (~^(-reg169[(4'hd):(3'h4)]))});
              reg281 <= $signed(reg243[(3'h5):(2'h2)]);
            end
          else
            begin
              reg280 = reg260[(2'h3):(2'h3)];
              reg282 = $signed(($signed(reg279) > reg277[(4'h8):(3'h6)]));
              reg283 <= ($signed(($unsigned($signed((8'h9e))) <<< $unsigned((~&(7'h47))))) ?
                  (8'ha4) : (^(&(~|(~&reg282)))));
              reg284 = ((|$signed($signed((reg260 ?
                  forvar259 : reg269)))) | ($unsigned($signed(reg257)) >= $signed(($signed(reg252) > $signed((8'had))))));
            end
          for (forvar285 = (1'h0); (forvar285 < (2'h2)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg286 = reg132;
              reg287 = ({(~|$unsigned((~^reg266)))} || {(!(^reg228)), wire72});
              reg288 <= $unsigned((~&$signed(wire72[(3'h7):(2'h2)])));
              reg289 = $signed($signed($unsigned({reg253[(5'h12):(1'h1)],
                  $signed((8'hb6))})));
              reg290 = {reg151[(2'h3):(2'h3)],
                  $unsigned($unsigned($unsigned((~reg264)))),
                  {reg249, (+reg288)}};
            end
          if (({($unsigned($signed(forvar261)) ?
                  $unsigned($signed((7'h4c))) : reg218[(4'he):(3'h7)]),
              (^$unsigned(reg263[(3'h5):(2'h3)]))} - (($signed($signed(reg186)) && reg239) <<< (~((reg204 ?
                  reg167 : (7'h4f)) ?
              {(8'hbf), (8'haf), reg277} : {reg181})))))
            begin
              reg291 <= reg177;
              reg292 = (~&(8'hab));
              reg293 <= $signed($unsigned(reg206));
              reg294 = wire74;
              reg295 <= (-(~^$unsigned(reg210[(4'h9):(1'h1)])));
            end
          else
            begin
              reg292 = $unsigned((reg168[(4'hb):(2'h3)] ?
                  $signed($unsigned($signed((7'h53)))) : {($signed(reg264) + reg152[(1'h0):(1'h0)])}));
            end
        end
      if ((({forvar285[(2'h2):(1'h0)],
          {(reg108 != forvar242),
              (reg279 ? reg152 : wire77),
              $unsigned(reg254)},
          $signed((^~(7'h41)))} ^ ((^~(reg253 ? (7'h57) : reg175)) ?
          ({reg234} ~^ {(8'hba)}) : ($unsigned(reg289) != reg258))) < (-$unsigned(reg259))))
        begin
          reg296 <= (~^reg278);
          reg297 = reg271;
          reg298 = (^~(reg297 ? $signed($signed((8'ha8))) : wire164));
          reg299 <= $unsigned((+(~^{{(8'hb6)}, (-(8'haa))})));
          reg300 = reg178[(5'h1d):(5'h14)];
          for (forvar301 = (1'h0); (forvar301 < (3'h4)); forvar301 = (forvar301 + (1'h1)))
            begin
              reg302 <= $signed((reg252 >>> $unsigned(reg136)));
              reg303 = $unsigned(reg242[(5'h13):(4'ha)]);
              reg304 <= reg205[(4'h9):(3'h7)];
            end
          if (reg274[(2'h2):(2'h2)])
            begin
              reg305 <= (!((&$unsigned(reg250)) ?
                  ($unsigned((reg134 ?
                      reg264 : reg253)) + $unsigned((7'h42))) : ($unsigned((8'hb2)) > $unsigned($signed(reg276)))));
              reg306 = {(reg294[(5'h10):(3'h5)] ?
                      reg158 : (reg134[(4'ha):(2'h3)] == {(^(8'hbe)),
                          $signed(reg270)}))};
              reg307 <= (^~reg133);
              reg308 = $signed(({reg162[(2'h3):(2'h2)]} >> ((^~$unsigned(reg265)) ?
                  $signed(reg303) : (!$unsigned(wire164)))));
              reg309 = reg213;
            end
          else
            begin
              reg305 <= $unsigned({(reg181[(4'hc):(2'h2)] ^ ($signed((7'h42)) ?
                      (reg201 + (8'hb1)) : (reg258 ? reg205 : reg251)))});
              reg306 = $signed((reg217[(2'h3):(2'h3)] ?
                  reg281[(2'h3):(1'h1)] : $signed(reg218[(5'h11):(2'h2)])));
              reg307 <= ({$signed($unsigned(reg268)),
                  $unsigned(($unsigned((7'h4d)) ?
                      (reg201 || reg104) : {reg200}))} ^ {reg218[(2'h3):(2'h3)]});
              reg308 = $signed(reg280);
              reg309 = {$unsigned({(reg260 ?
                          reg219[(4'hc):(3'h7)] : $signed(forvar261)),
                      forvar301}),
                  reg262};
            end
        end
      else
        begin
          for (forvar296 = (1'h0); (forvar296 < (3'h4)); forvar296 = (forvar296 + (1'h1)))
            begin
              reg299 <= $signed(reg261);
              reg300 = reg248;
              reg301 = $signed((reg165 * ((reg248 ?
                      (~wire77) : $unsigned(reg141)) ?
                  ($unsigned(reg83) ?
                      ((8'h9c) <<< reg271) : (reg279 ?
                          reg228 : reg142)) : ({reg245, reg213} & (forvar261 ?
                      reg270 : reg261)))));
            end
          for (forvar302 = (1'h0); (forvar302 < (3'h6)); forvar302 = (forvar302 + (1'h1)))
            begin
              reg304 <= reg290;
              reg305 <= $signed((^reg303[(1'h1):(1'h1)]));
            end
          if (({reg194[(4'hc):(1'h1)],
              $signed($signed({reg117})),
              {(&(reg98 ? forvar302 : reg309))}} && (wire241[(5'h16):(4'he)] ?
              reg228[(1'h1):(1'h0)] : (^reg171[(4'hf):(4'he)]))))
            begin
              reg307 <= reg252;
              reg308 = {((reg309[(2'h3):(1'h1)] || ($signed(reg213) >>> (reg83 ?
                      reg247 : reg130))) < reg255[(2'h2):(2'h2)])};
            end
          else
            begin
              reg307 <= $unsigned($signed($signed($signed((reg191 & reg205)))));
              reg308 = {{(7'h4e),
                      (reg259 ? reg257[(4'hf):(1'h0)] : $unsigned(reg287))}};
            end
          if ((~|$signed((reg308[(5'h17):(2'h2)] < (~$signed(reg260))))))
            begin
              reg310 <= (!$signed($signed(reg108)));
            end
          else
            begin
              reg310 <= (($signed((reg276 > (~|wire78))) != $unsigned($unsigned((!reg182)))) ?
                  {(+((reg120 ? reg298 : reg152) ? (8'hbf) : (~|reg269))),
                      {forvar296,
                          reg302,
                          reg134}} : $signed($signed((~{reg301}))));
              reg311 <= $unsigned($signed((+(~(~(7'h55))))));
              reg312 <= reg279[(3'h7):(3'h4)];
              reg313 <= $unsigned($signed($unsigned($signed(reg108))));
              reg314 <= (-{{((!(8'ha6)) * $signed((8'ha5))), (8'hbe)},
                  ({reg292[(1'h0):(1'h0)]} ?
                      (|{wire72,
                          reg177,
                          reg262}) : $unsigned($unsigned(reg265)))});
              reg315 <= $unsigned(reg129[(4'h8):(2'h3)]);
            end
          for (forvar316 = (1'h0); (forvar316 < (1'h1)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg317 = (reg308[(5'h10):(3'h5)] ?
                  reg213[(4'hc):(3'h5)] : $signed(($unsigned((reg186 ?
                      reg268 : (8'h9e))) - ((-reg129) ?
                      (reg309 ? reg165 : forvar285) : {reg306}))));
              reg318 = (7'h58);
              reg319 = $signed($unsigned($signed(reg295[(4'hf):(1'h1)])));
              reg320 <= (^(+($unsigned(reg281) ?
                  {reg228[(2'h3):(1'h1)],
                      (~(7'h4d)),
                      wire164[(3'h5):(2'h3)]} : reg252[(3'h4):(2'h3)])));
              reg321 <= $signed({$unsigned(((reg263 <<< reg102) & (reg249 ?
                      reg258 : reg277)))});
            end
          if (reg253)
            begin
              reg322 <= (8'ha8);
              reg323 = reg300;
              reg324 <= (|$unsigned($signed((8'haa))));
              reg325 <= reg232;
            end
          else
            begin
              reg323 = forvar316;
            end
        end
    end
  module326 #() modinst684 (wire683, clk, reg111, reg158, reg171, reg191, reg254);
  always
    @(posedge clk) begin
      reg685 = ({{(&wire241[(3'h7):(1'h1)]),
              $unsigned((reg205 ?
                  reg182 : reg233))}} && $signed(((&$unsigned(reg102)) ?
          {((8'h9c) ? reg281 : reg132), $signed(reg83)} : (~&reg158))));
      reg686 <= reg322;
      if ((reg177[(5'h11):(5'h11)] ? reg288 : (7'h45)))
        begin
          for (forvar687 = (1'h0); (forvar687 < (1'h0)); forvar687 = (forvar687 + (1'h1)))
            begin
              reg688 = ($signed($signed((~&(+wire163)))) == $unsigned($signed($unsigned((reg322 < reg151)))));
            end
          if ($signed(reg206[(5'h15):(5'h10)]))
            begin
              reg689 = (|$unsigned((((reg264 ? reg142 : reg248) ?
                      (&reg234) : $signed(reg281)) ?
                  reg686 : $unsigned((reg262 ? (8'hbb) : reg217)))));
              reg690 = reg268;
              reg691 = reg195;
              reg692 <= reg276[(2'h3):(1'h0)];
              reg693 = {($signed(($unsigned(reg141) != (reg182 | reg266))) * (^~(|(reg167 * reg175))))};
              reg694 = (reg195 ?
                  $signed({(!reg175),
                      reg307[(4'ha):(3'h4)],
                      (reg113 >> $unsigned(reg200))}) : ((~(+{(7'h4d),
                      reg293})) && ($unsigned(reg125[(4'he):(4'h8)]) ?
                      reg175 : $unsigned((~(8'hbc))))));
            end
          else
            begin
              reg692 <= $unsigned(($unsigned(reg320) + reg253));
              reg695 <= (~^reg311[(4'hd):(1'h0)]);
              reg696 <= $unsigned($unsigned(($unsigned(reg117) == reg689)));
              reg697 = $signed(((wire79 >> $unsigned(((8'hb4) < (8'h9d)))) ~^ ($unsigned((reg177 ?
                      reg269 : (7'h41))) ?
                  (reg233 * reg694[(1'h0):(1'h0)]) : ($signed((7'h43)) ?
                      (reg302 ? reg270 : wire164) : $unsigned(reg296)))));
            end
        end
      else
        begin
          reg687 <= ($signed((((reg145 ?
                  (8'h9f) : reg219) >> $signed(reg178)) | (&(reg130 ?
                  reg186 : wire74)))) ?
              reg275 : reg186);
        end
      if (reg258)
        begin
          if (reg320[(3'h4):(3'h4)])
            begin
              reg698 = {$unsigned((reg200[(4'h9):(2'h2)] ?
                      {$unsigned(reg299),
                          (reg162 ? reg304 : reg191),
                          (!(8'hb4))} : $unsigned($signed(reg274)))),
                  reg268};
              reg699 <= (($unsigned(($signed(reg234) && $unsigned((8'hb2)))) | (^~(reg186[(1'h0):(1'h0)] < reg311[(4'hb):(3'h4)]))) ?
                  $signed((reg152[(2'h3):(2'h2)] > $signed(reg171))) : $unsigned($unsigned((!(reg305 ^ reg258)))));
              reg700 = {(reg314 >= ($unsigned($unsigned(reg151)) ^~ (~&wire74))),
                  ($signed($signed(reg695[(1'h1):(1'h1)])) ^~ $signed((8'hb1)))};
            end
          else
            begin
              reg699 <= ($signed($signed(reg293)) ?
                  ((~reg288[(4'hd):(2'h2)]) ?
                      (~reg218[(2'h2):(1'h0)]) : $unsigned($signed($unsigned((8'hba))))) : $unsigned((reg288[(3'h7):(3'h5)] - (&(wire79 ?
                      reg169 : reg305)))));
              reg701 <= (|{reg257,
                  ($unsigned(reg206) ? $unsigned($unsigned(reg218)) : reg291),
                  ((wire76 ? reg83[(5'h10):(4'hf)] : reg691) ?
                      ({reg217} - reg152[(2'h3):(2'h2)]) : reg325[(4'h8):(3'h7)])});
              reg702 = (-reg213);
              reg703 = {reg693[(3'h6):(2'h2)],
                  ($unsigned({wire77[(3'h6):(3'h6)],
                      reg162}) < ((reg158[(5'h18):(1'h0)] ?
                      (7'h42) : (reg697 ?
                          reg264 : wire79)) ^ $unsigned((~&reg186))))};
              reg704 = {$signed($unsigned(reg698)),
                  ($unsigned(((reg701 - reg291) ?
                      reg281[(2'h2):(1'h1)] : (reg276 ?
                          reg279 : reg275))) >>> $unsigned({(wire683 ^ reg320),
                      (wire164 ? reg281 : reg178),
                      reg135})),
                  ($signed((^~(~&reg693))) ?
                      $signed(reg696[(2'h2):(1'h0)]) : ({(reg699 ?
                              reg255 : reg322),
                          reg702} <= (^(!reg111))))};
              reg705 <= reg266[(4'h8):(2'h2)];
              reg706 = ((^~$unsigned(reg293[(2'h2):(1'h1)])) ?
                  $signed(reg234) : reg266[(2'h2):(2'h2)]);
            end
          reg707 = $signed({$signed((forvar687 * reg178))});
          if (reg115[(4'h8):(2'h3)])
            begin
              reg708 <= (~(reg692[(3'h5):(1'h1)] ?
                  reg283 : reg213[(4'hd):(3'h4)]));
              reg709 = reg708[(4'hb):(3'h6)];
              reg710 <= $signed((8'hb6));
            end
          else
            begin
              reg708 <= (~&(+forvar687));
            end
          if ({{reg145,
                  $unsigned(reg693[(3'h5):(2'h2)]),
                  (((reg125 ? reg703 : reg233) ?
                      (reg257 ?
                          (8'hb5) : wire163) : reg262[(4'h8):(2'h2)]) * reg703[(2'h3):(1'h0)])},
              reg685[(1'h1):(1'h1)]})
            begin
              reg711 <= (reg283 ^ (7'h4c));
              reg712 = reg130[(3'h4):(1'h1)];
              reg713 = reg686;
              reg714 <= ({(((~reg158) + reg104) <= ($unsigned(reg195) || (~|reg168)))} ?
                  $unsigned($signed(((reg307 ? reg125 : reg692) ?
                      {(7'h4d), reg701} : $unsigned(reg168)))) : reg253);
              reg715 <= {($signed(reg695) ?
                      (~^(~^(~|reg293))) : $unsigned((-reg182[(5'h1e):(4'he)])))};
              reg716 <= ($signed($signed(((reg714 ~^ wire76) + {reg713}))) ^ (reg268 <<< ($unsigned(reg222) ?
                  $unsigned($unsigned(reg169)) : $unsigned(forvar687[(2'h3):(2'h3)]))));
              reg717 = (-($unsigned(reg228) ^ $unsigned(reg257)));
            end
          else
            begin
              reg711 <= $unsigned(wire79[(2'h3):(1'h0)]);
              reg714 <= ({{(~^(7'h4a)),
                          {reg111[(4'he):(1'h1)], reg262, $unsigned(reg307)}},
                      reg713[(2'h3):(1'h1)],
                      reg218[(4'ha):(1'h1)]} ?
                  $unsigned((reg688 ?
                      $signed(reg135) : reg169[(4'h8):(3'h4)])) : $unsigned(reg716[(5'h12):(4'he)]));
              reg717 = ((&$signed({(+(8'hb0)), (8'h9f)})) ?
                  reg310 : (reg111[(4'h9):(3'h6)] << {$signed((wire683 ?
                          (7'h47) : reg121)),
                      {{reg162}, $unsigned((8'ha8)), $signed((7'h42))}}));
            end
          reg718 <= $unsigned($signed({(reg206[(3'h5):(2'h2)] ?
                  (reg696 ^~ reg314) : $signed(reg130)),
              reg305}));
        end
      else
        begin
          reg699 <= $signed((reg260[(4'hb):(1'h1)] >> (((^reg693) || $unsigned(reg134)) || reg299)));
          for (forvar700 = (1'h0); (forvar700 < (2'h3)); forvar700 = (forvar700 + (1'h1)))
            begin
              reg702 = ($signed(($unsigned((&reg255)) ?
                  ($signed(reg693) ?
                      (~reg178) : $signed((8'ha5))) : ((reg305 == reg251) ?
                      (reg311 ?
                          reg219 : (7'h50)) : $signed(reg262)))) << ($unsigned(reg701[(4'ha):(3'h5)]) ?
                  reg145 : (~&$unsigned(reg266[(2'h3):(2'h3)]))));
              reg703 = wire73[(2'h2):(1'h0)];
              reg705 <= wire164[(4'hb):(1'h1)];
              reg706 = reg200[(4'h8):(3'h6)];
              reg708 <= ((^~$signed({(reg703 ? (8'hb5) : reg313)})) ?
                  {({reg217, reg716[(4'hf):(4'hb)]} == reg688),
                      $signed(reg182),
                      (reg321 ?
                          (~$unsigned((7'h56))) : reg694)} : $unsigned(($unsigned((reg702 <= reg325)) ?
                      (wire241 ^~ (8'hb7)) : $unsigned((8'ha8)))));
              reg710 <= $signed((reg261[(5'h11):(4'hf)] ?
                  reg313 : ($signed(forvar700) ^~ ((reg295 >>> (7'h41)) > (+wire241)))));
            end
          reg712 = ($unsigned(reg239[(3'h6):(3'h4)]) ~^ $signed(reg255));
          reg714 <= ((~reg204[(4'h9):(3'h7)]) ?
              {reg158,
                  wire77[(2'h2):(1'h0)],
                  {(+(reg205 ? reg269 : reg117)),
                      $signed($unsigned(reg130)),
                      ((reg186 ?
                          reg703 : reg218) >> reg713)}} : {reg293[(1'h1):(1'h0)],
                  reg713[(3'h7):(2'h2)],
                  wire76});
          for (forvar715 = (1'h0); (forvar715 < (1'h0)); forvar715 = (forvar715 + (1'h1)))
            begin
              reg716 <= $signed($signed((^~$unsigned(reg270))));
              reg718 <= {$signed($signed($unsigned((reg274 ?
                      (8'ha0) : reg321)))),
                  $signed((((forvar687 ^ reg134) ?
                          ((8'hbb) ? reg299 : wire78) : reg278) ?
                      (^~{reg275}) : $unsigned((reg288 ? wire75 : reg89))))};
              reg719 <= (reg275[(1'h0):(1'h0)] ^ wire241);
              reg720 = reg325;
            end
          for (forvar721 = (1'h0); (forvar721 < (3'h5)); forvar721 = (forvar721 + (1'h1)))
            begin
              reg722 = reg254[(2'h2):(1'h0)];
              reg723 <= $signed((!$unsigned(reg251)));
            end
        end
      if (reg102[(5'h17):(3'h7)])
        begin
          reg724 <= ($unsigned(reg108) | $unsigned(reg691[(3'h4):(2'h2)]));
          reg725 = (8'hb1);
          reg726 = $unsigned(($signed($signed((reg283 & reg98))) ?
              ((8'ha7) ^~ reg276[(2'h3):(1'h1)]) : reg715));
        end
      else
        begin
          if ((($signed(reg168[(4'h8):(3'h5)]) ?
              $signed((~^$unsigned((8'h9c)))) : reg689[(3'h4):(1'h1)]) < ($unsigned($signed((8'ha3))) ?
              (^~{$unsigned(reg315),
                  reg687[(5'h10):(4'h8)],
                  {(8'hb1), reg714}}) : ((reg281 ?
                      (reg104 ? reg725 : reg268) : (-reg713)) ?
                  $unsigned(reg312[(4'h9):(4'h9)]) : $unsigned(((7'h4d) ?
                      reg713 : (7'h56)))))))
            begin
              reg724 <= (8'hbf);
              reg725 = (reg288[(3'h7):(1'h1)] ?
                  (|$signed(((~reg263) | (reg134 ?
                      (7'h4d) : reg295)))) : (^~{(&(reg206 ?
                          (8'ha5) : reg253))}));
            end
          else
            begin
              reg724 <= $signed($unsigned(reg312[(4'hb):(4'hb)]));
              reg725 = reg83[(3'h6):(3'h6)];
              reg726 = reg182[(5'h16):(5'h13)];
            end
          reg727 <= ($signed(((+$signed(reg125)) ?
                  ((reg315 != reg705) ?
                      (reg130 > reg313) : reg689[(2'h2):(2'h2)]) : ((reg687 <<< reg283) <<< (reg283 && reg256)))) ?
              $signed({reg291[(3'h6):(3'h6)],
                  reg120[(3'h7):(1'h1)]}) : $unsigned(reg111[(4'hf):(2'h2)]));
          reg728 <= reg191;
          reg729 = (&reg276[(1'h1):(1'h0)]);
        end
    end
  assign wire730 = {$signed((reg209[(4'hc):(4'hc)] ?
                           {reg315, reg276, (~reg232)} : ($unsigned((8'h9c)) ?
                               ((8'hb0) ?
                                   reg314 : reg716) : $unsigned(reg270)))),
                       reg200[(1'h1):(1'h1)]};
  always
    @(posedge clk) begin
      for (forvar731 = (1'h0); (forvar731 < (3'h6)); forvar731 = (forvar731 + (1'h1)))
        begin
          reg732 = $signed(((|reg281) || ($signed((reg89 ? wire730 : reg167)) ?
              (reg132[(3'h7):(3'h6)] ?
                  $signed((7'h52)) : (~reg696)) : reg270)));
          if ({(reg219 ? $unsigned($unsigned($unsigned(reg132))) : (7'h49))})
            begin
              reg733 = $unsigned(($signed(reg113[(4'hd):(3'h4)]) + reg142));
              reg734 = $signed(($signed($unsigned(reg296)) >>> (wire730 ?
                  ((+reg135) ? (+reg152) : (|reg299)) : ((reg239 <<< reg182) ?
                      reg98 : {reg262}))));
              reg735 <= ($signed($signed(($unsigned(reg262) ?
                  (~^reg102) : {reg705,
                      reg251,
                      (7'h52)}))) == $signed($signed($unsigned(reg213))));
              reg736 = ($unsigned(reg254) == $unsigned(reg695));
            end
          else
            begin
              reg735 <= $signed((wire164[(4'hb):(4'hb)] < {$signed(reg735[(1'h0):(1'h0)]),
                  (8'hbb)}));
              reg737 <= $signed($unsigned((reg205[(4'hf):(4'hf)] ?
                  reg83[(5'h12):(5'h10)] : (reg121[(4'hc):(4'hc)] == $unsigned((7'h53))))));
              reg738 = reg213;
              reg739 = (wire77 ?
                  $signed($signed($signed($unsigned((7'h42))))) : (~^$signed(($unsigned(reg304) ^~ (+reg171)))));
              reg740 <= reg204[(3'h5):(1'h0)];
            end
          reg741 <= ($unsigned((!reg310[(1'h1):(1'h0)])) ?
              (~(~&$signed(reg152))) : $unsigned(((reg276[(3'h4):(3'h4)] ?
                  (reg181 ? reg695 : (8'hac)) : ((7'h54) ?
                      (8'hb1) : reg168)) < ((~|reg145) ?
                  (reg133 >= (8'ha6)) : $signed(reg263)))));
          if (reg152[(1'h1):(1'h1)])
            begin
              reg742 <= ({((forvar731[(4'he):(4'ha)] || (reg291 ?
                          (8'hb8) : reg194)) - (~(|reg724))),
                      ({(~^reg701), (reg165 ? wire241 : reg191)} > ((reg134 ?
                              reg260 : reg165) ?
                          $signed(reg283) : $unsigned(reg182)))} ?
                  ($unsigned(reg699[(5'h15):(3'h7)]) ^~ $signed(((reg141 ?
                      wire77 : reg205) && (reg296 ?
                      reg136 : reg699)))) : ($signed($unsigned($unsigned(wire74))) ?
                      reg117 : (!reg90)));
              reg743 <= ((wire78[(4'h9):(1'h0)] ?
                      reg268[(1'h1):(1'h1)] : {($signed(reg169) | reg711[(4'h8):(1'h1)]),
                          {(reg708 ? reg295 : reg723)},
                          reg228}) ?
                  (^~($signed({wire241,
                      reg158,
                      reg296}) | reg732)) : (~$unsigned((~|((8'haf) ?
                      reg719 : (8'h9c))))));
              reg744 = reg257[(5'h1e):(5'h1b)];
            end
          else
            begin
              reg744 = {($unsigned(((8'ha2) != $signed(reg182))) >= $unsigned(({(8'ha8),
                      reg314} != $unsigned(reg171))))};
              reg745 = (~&reg304[(4'hf):(3'h6)]);
              reg746 <= (~&$unsigned($unsigned({reg217})));
              reg747 = ({(reg177 ?
                          (&$unsigned(reg195)) : reg206[(2'h3):(2'h2)]),
                      $unsigned((^~wire683[(2'h2):(1'h0)]))} ?
                  (+$unsigned((~$unsigned(reg195)))) : ($signed((reg262[(2'h2):(1'h0)] ?
                          (reg254 ? reg741 : wire241) : reg254)) ?
                      $signed(({reg715, reg234, reg291} ?
                          $signed(reg719) : (reg740 ?
                              wire77 : reg121))) : reg304));
              reg748 = $signed(((({wire164} ?
                          $signed(reg257) : (reg142 * reg743)) ?
                      $unsigned(reg151) : $signed((~^reg302))) ?
                  {(^(~^reg687))} : reg747));
              reg749 = $unsigned((($unsigned($unsigned(reg283)) * reg191[(3'h5):(2'h2)]) ?
                  (7'h46) : (^~(|{reg125, reg175, reg182}))));
              reg750 = (~(7'h50));
            end
          reg751 = reg699[(4'hc):(3'h6)];
          for (forvar752 = (1'h0); (forvar752 < (3'h5)); forvar752 = (forvar752 + (1'h1)))
            begin
              reg753 = (((~wire77) ?
                  $unsigned(($signed(reg205) ?
                      reg714[(3'h6):(2'h3)] : (reg718 ?
                          wire164 : reg145))) : (reg209[(4'hd):(4'h9)] ?
                      reg324 : (((8'h9e) ? reg256 : reg738) ?
                          reg182[(5'h16):(5'h15)] : (+reg718)))) << (-(reg283 ?
                  (-$signed(reg737)) : reg117)));
              reg754 = reg266[(5'h12):(1'h0)];
              reg755 = $signed($signed({reg191[(2'h2):(1'h0)],
                  ((reg168 ? reg747 : reg746) ?
                      ((8'h9f) ? reg83 : (7'h50)) : {reg234})}));
              reg756 <= $unsigned($unsigned((&(~|{(7'h46), reg204, reg304}))));
              reg757 <= reg218;
              reg758 = {$signed(reg213[(3'h5):(2'h2)]),
                  (reg756 << $signed($signed({reg171, (7'h4b), reg232})))};
              reg759 = $signed(reg228);
            end
        end
      if ((~|((((reg206 * reg696) < (&reg194)) ?
          wire730[(5'h16):(2'h3)] : $unsigned($signed(reg248))) <= $unsigned(((reg90 >>> reg274) >= $unsigned((8'hb6)))))))
        begin
          for (forvar760 = (1'h0); (forvar760 < (1'h0)); forvar760 = (forvar760 + (1'h1)))
            begin
              reg761 = $unsigned(reg130);
              reg762 = $unsigned($signed(((~|{wire241,
                  reg711,
                  reg264}) << $unsigned(reg186))));
              reg763 <= (~^reg175);
              reg764 <= (({$signed($unsigned(reg279))} ?
                      (!$unsigned((^reg734))) : reg701[(4'h8):(3'h5)]) ?
                  ((~reg738) || (7'h53)) : (^~({$unsigned(reg755),
                      (^reg761),
                      $unsigned(reg90)} - ($signed(reg260) ?
                      $signed(reg746) : $signed(reg276)))));
            end
          reg765 = {(+(~^$signed($unsigned(reg736)))),
              reg256[(4'hc):(4'ha)],
              (~{(-reg262[(2'h3):(1'h1)])})};
          if ((&($unsigned($signed((reg205 ? reg239 : reg201))) ?
              $signed($signed((reg191 <= reg108))) : ($signed((-reg746)) & $unsigned((&reg269))))))
            begin
              reg766 = reg313;
              reg767 = {reg733};
              reg768 <= reg741[(4'hb):(4'h9)];
              reg769 = (8'ha1);
              reg770 <= ((&{$signed($signed((7'h48))),
                      reg233,
                      $signed((|reg182))}) ?
                  ($unsigned(wire163) >>> reg732[(5'h14):(4'hf)]) : $unsigned($signed($unsigned((^(8'had))))));
              reg771 <= $signed($signed(reg134));
            end
          else
            begin
              reg766 = $unsigned((7'h49));
              reg768 <= ((~|wire76) ?
                  (~|(reg724[(3'h5):(1'h1)] > ($unsigned(reg262) ?
                      reg275[(5'h10):(2'h2)] : ((7'h44) ?
                          reg213 : reg145)))) : reg275);
              reg769 = (!((^(~|$unsigned(wire74))) ?
                  (!reg291[(4'h9):(3'h6)]) : (-(((8'h9d) - reg763) ?
                      reg320 : (|reg133)))));
              reg770 <= $unsigned(reg276);
              reg771 <= {$signed(wire77)};
              reg772 <= $unsigned((~^$unsigned((((7'h54) ? reg711 : reg135) ?
                  reg736 : (8'hbb)))));
              reg773 <= $unsigned(($signed($signed(reg125)) ?
                  reg228 : ($signed($unsigned(reg228)) ?
                      reg734 : $signed((wire76 ^ reg177)))));
            end
        end
      else
        begin
          for (forvar760 = (1'h0); (forvar760 < (2'h2)); forvar760 = (forvar760 + (1'h1)))
            begin
              reg763 <= (~&((~|reg743[(1'h0):(1'h0)]) >>> $unsigned(((reg83 ?
                      reg772 : reg773) ?
                  reg761 : (!reg767)))));
              reg764 <= (+{(($unsigned((8'had)) ?
                      (8'hac) : (reg264 ?
                          reg175 : (7'h48))) < ($signed(wire241) ?
                      {reg266} : (reg686 << reg120)))});
              reg768 <= $unsigned(((reg227 ?
                  $signed($unsigned(reg275)) : reg256[(4'he):(3'h5)]) == $signed(reg257[(5'h14):(4'he)])));
              reg770 <= (+(+$signed(($signed(wire78) ?
                  {reg175, wire163, reg136} : reg742[(5'h10):(4'hd)]))));
              reg771 <= $unsigned((|((reg263 ?
                  $unsigned(reg763) : $unsigned(reg710)) > (7'h52))));
              reg774 = reg162;
            end
        end
      reg775 <= (reg756 ? $signed((~|(!(reg305 >>> reg256)))) : {reg194});
      reg776 <= (($unsigned($signed($signed(reg104))) ?
          reg295 : (($unsigned((7'h46)) + (reg248 ?
              wire72 : wire240)) | (reg761 ?
              reg158 : (8'hb1)))) ^~ ({(reg740 && ((8'hb0) || wire74))} ?
          reg253 : (reg743 > ((reg133 ? reg733 : reg111) ?
              $signed(forvar760) : wire241[(4'hb):(3'h7)]))));
      reg777 = reg746[(2'h3):(2'h2)];
      reg778 = $signed($unsigned($unsigned(reg304[(5'h14):(4'h8)])));
      if (((^~(({reg743, reg291, (7'h46)} >>> $signed(reg167)) ~^ reg177)) ?
          $unsigned($signed($unsigned((reg777 && reg774)))) : $unsigned((~(reg711 ?
              $unsigned(wire163) : reg759[(1'h0):(1'h0)])))))
        begin
          for (forvar779 = (1'h0); (forvar779 < (3'h4)); forvar779 = (forvar779 + (1'h1)))
            begin
              reg780 = $signed($unsigned($signed(((8'hb0) ?
                  (reg291 ? reg305 : reg747) : $unsigned(wire79)))));
              reg781 <= reg228;
            end
          reg782 <= {(|(reg256 != reg745[(2'h3):(2'h3)])), reg315};
          reg783 <= ($unsigned($unsigned($unsigned((reg742 | (8'hb6))))) != reg766[(2'h3):(2'h2)]);
          reg784 <= reg218[(3'h7):(3'h7)];
        end
      else
        begin
          reg779 = (~^((+(^(^(8'hac)))) ?
              wire77 : ($signed(reg261) ?
                  ((wire730 - reg781) != $signed(reg135)) : ((reg716 + reg302) ?
                      reg748 : (~&reg719)))));
          if ({reg222[(4'h8):(2'h3)], $unsigned(reg753), reg769})
            begin
              reg780 = $unsigned(reg766);
              reg785 = (reg217[(4'h8):(4'h8)] | (|$unsigned(($unsigned(reg775) ?
                  (reg130 & (8'h9d)) : $unsigned(reg322)))));
              reg786 = reg687;
              reg787 = {reg89,
                  $signed(((~|(reg233 ?
                      reg749 : reg167)) <= $unsigned(((7'h42) ?
                      reg213 : reg758))))};
              reg788 = (!(~^({$unsigned(wire72)} >= $unsigned((&forvar731)))));
            end
          else
            begin
              reg780 = {$unsigned((|$signed((reg218 ? reg90 : reg248)))),
                  reg763};
              reg785 = reg744[(2'h3):(2'h3)];
              reg786 = (!(~^reg777[(5'h10):(3'h4)]));
              reg787 = $unsigned($unsigned(reg756));
            end
          reg789 = (|$unsigned($signed((|$unsigned(reg142)))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar790 = (1'h0); (forvar790 < (1'h0)); forvar790 = (forvar790 + (1'h1)))
        begin
          reg791 <= reg205[(3'h7):(2'h2)];
          if ((~&reg255))
            begin
              reg792 = ($signed(reg263) ?
                  $signed((~|{(reg768 ? reg169 : reg274),
                      (reg263 ? (8'hb0) : reg701),
                      reg260[(5'h1d):(5'h1a)]})) : $unsigned(((&(7'h4f)) - $unsigned(reg178[(5'h1c):(4'hc)]))));
              reg793 <= ($unsigned($unsigned(reg260)) ?
                  $unsigned($signed((~|reg262))) : (forvar790[(3'h4):(2'h3)] ^~ (8'h9e)));
              reg794 = $signed(reg90[(4'hf):(1'h0)]);
              reg795 = reg145;
              reg796 = $unsigned(($unsigned($signed(reg325)) ?
                  ((reg264 ? (!reg743) : (wire683 ? reg274 : reg270)) ?
                      (reg281[(4'h8):(3'h6)] ~^ (reg218 ?
                          (8'hb5) : reg253)) : reg701[(4'hd):(4'ha)]) : $signed(((reg206 <= reg260) ?
                      wire74 : (reg263 ? reg248 : reg98)))));
              reg797 = (({((+(8'ha7)) >> (~reg200)),
                      (reg165[(3'h5):(3'h5)] << reg775[(1'h0):(1'h0)]),
                      (8'had)} > (!($unsigned(reg746) >= ((8'hb7) ^~ reg254)))) ?
                  $signed(reg256) : (^~(((reg315 << (8'hae)) >>> $signed(reg98)) <<< (reg232[(5'h1d):(5'h1d)] ?
                      $signed(reg194) : $signed(reg723)))));
              reg798 = (~&wire75[(4'he):(3'h6)]);
            end
          else
            begin
              reg792 = reg256;
              reg793 <= reg186;
              reg799 <= reg756[(1'h0):(1'h0)];
              reg800 <= reg276;
            end
          for (forvar801 = (1'h0); (forvar801 < (3'h6)); forvar801 = (forvar801 + (1'h1)))
            begin
              reg802 <= $unsigned(reg699);
              reg803 <= (((^reg716[(4'hd):(1'h1)]) ?
                  ((~&reg715[(3'h4):(2'h3)]) ?
                      reg158 : {reg263[(3'h4):(2'h3)],
                          reg113[(5'h1b):(5'h10)]}) : reg210) && $signed($signed({$signed((7'h43)),
                  $unsigned((7'h54))})));
              reg804 = ((-($signed((reg200 || reg312)) << reg737)) ?
                  (reg737 ^~ (-$signed(((8'hb9) || reg262)))) : ((((~reg209) ?
                      reg186 : $signed(reg90)) || reg295[(5'h10):(1'h1)]) ~^ $signed(reg687[(1'h0):(1'h0)])));
              reg805 <= reg262;
              reg806 <= ((reg262 ^ (reg794 - {$signed(reg723),
                      $signed(reg195),
                      (reg735 ? reg305 : reg310)})) ?
                  $signed(($unsigned($signed((7'h56))) ?
                      $signed(reg800[(1'h1):(1'h1)]) : ({reg130,
                          reg167,
                          reg227} | (reg268 ? reg716 : wire241)))) : reg232);
              reg807 <= (~reg168[(2'h3):(1'h1)]);
              reg808 <= (+(+wire241));
            end
        end
      reg809 <= $signed($unsigned(reg293[(2'h2):(1'h1)]));
      for (forvar810 = (1'h0); (forvar810 < (3'h4)); forvar810 = (forvar810 + (1'h1)))
        begin
          if ($unsigned(((!$unsigned({reg195})) ^~ (reg324[(2'h2):(1'h0)] ^ $signed((reg256 ~^ reg260))))))
            begin
              reg811 <= reg191;
              reg812 = ($unsigned({($unsigned(reg743) != $unsigned(reg218)),
                  (reg136[(2'h3):(1'h1)] * (reg228 ?
                      reg797 : reg186))}) ~^ (|$unsigned({reg708[(4'he):(1'h1)],
                  $signed(reg278),
                  (reg756 && reg227)})));
              reg813 <= (!(reg716 ?
                  $signed($unsigned((reg268 ?
                      reg152 : reg757))) : ((^~(reg313 <<< reg701)) ?
                      ((reg781 & reg304) ?
                          (reg102 ?
                              reg205 : reg741) : $unsigned((8'hae))) : ({reg268} ?
                          ((8'hbb) ?
                              reg756 : (8'ha7)) : reg181[(4'he):(1'h0)]))));
              reg814 <= reg710[(1'h1):(1'h0)];
            end
          else
            begin
              reg811 <= reg802[(4'hc):(4'hb)];
              reg813 <= {((+{(reg152 ? wire79 : reg814),
                      reg715[(1'h0):(1'h0)],
                      {reg264, reg718}}) <<< reg718[(4'hf):(3'h7)]),
                  reg181};
              reg814 <= $unsigned((!$unsigned($signed((reg723 & reg194)))));
              reg815 = ($unsigned(reg321) ~^ reg256[(3'h5):(2'h2)]);
              reg816 = (^$signed((reg727 ?
                  reg803 : ($unsigned(reg715) ?
                      $unsigned(reg130) : (reg171 ? reg293 : reg83)))));
            end
          for (forvar817 = (1'h0); (forvar817 < (1'h1)); forvar817 = (forvar817 + (1'h1)))
            begin
              reg818 <= (8'ha8);
              reg819 <= (+((reg807 * $unsigned({reg737,
                  reg310,
                  (8'hab)})) << {(~$signed(reg83)),
                  ((8'ha6) ? reg312 : $unsigned(reg111)),
                  ($signed(reg217) ?
                      ((8'ha1) ? reg115 : reg262) : {reg791, reg111})}));
            end
        end
      reg820 = reg258[(3'h4):(2'h2)];
      reg821 = (|(^(~^wire72[(2'h2):(1'h1)])));
      reg822 <= (~(reg816 * $unsigned((7'h50))));
      for (forvar823 = (1'h0); (forvar823 < (3'h5)); forvar823 = (forvar823 + (1'h1)))
        begin
          reg824 <= reg296;
          reg825 <= {reg152[(1'h1):(1'h1)], $signed(reg256)};
          for (forvar826 = (1'h0); (forvar826 < (3'h6)); forvar826 = (forvar826 + (1'h1)))
            begin
              reg827 <= ($signed($unsigned(reg312)) ?
                  ($unsigned($signed(reg142[(2'h2):(1'h1)])) >>> reg692[(2'h2):(1'h0)]) : (forvar823 ?
                      reg162 : (~|($unsigned(reg803) ?
                          $unsigned(reg727) : ((7'h55) ? reg117 : (8'h9f))))));
              reg828 = forvar801[(5'h16):(2'h3)];
              reg829 = (~$signed((reg312[(4'hb):(4'h9)] >= (7'h41))));
            end
          if (($unsigned((-$unsigned((reg716 ?
              reg178 : (7'h4b))))) << (($signed(forvar801) ?
                  reg228[(2'h3):(2'h2)] : $signed((7'h40))) ?
              (8'h9c) : $signed((~&(^~reg796))))))
            begin
              reg830 = $signed(((-reg182) ?
                  (reg796 ?
                      (reg302 <= (+reg239)) : ((-reg773) <= reg175)) : reg275[(2'h2):(2'h2)]));
              reg831 = reg740[(2'h2):(2'h2)];
              reg832 = (reg687 > $signed(reg162[(2'h3):(2'h3)]));
              reg833 <= $signed(reg718[(4'hc):(1'h0)]);
              reg834 = reg281;
              reg835 <= $signed((^~(^~($unsigned(wire76) ?
                  (reg728 - reg182) : reg776[(2'h2):(2'h2)]))));
            end
          else
            begin
              reg830 = (&reg782);
              reg833 <= ($unsigned(reg772) ?
                  (($unsigned(reg120) ~^ reg295) ?
                      $signed(((forvar810 ? (8'hb8) : reg737) ?
                          $unsigned((8'ha4)) : wire241[(5'h14):(3'h6)])) : $signed($signed((-reg182)))) : reg764[(4'hb):(4'h9)]);
              reg835 <= $unsigned(($signed(wire163) ?
                  (~reg132[(4'ha):(3'h4)]) : $unsigned($unsigned((reg830 ^~ (7'h55))))));
              reg836 <= $signed($signed({(reg165[(5'h12):(5'h12)] ?
                      (reg699 ? reg743 : (8'ha8)) : {(8'ha2)}),
                  reg699}));
              reg837 <= (((!((|reg227) ? wire76 : (reg321 + reg763))) ?
                  {reg232,
                      $signed($unsigned(reg833)),
                      $unsigned((reg793 ?
                          reg315 : (8'ha3)))} : reg821) ^~ $unsigned({$unsigned((8'hb9))}));
              reg838 = (((^(wire76[(1'h1):(1'h0)] ?
                      (reg210 ?
                          reg804 : (8'hb8)) : reg218)) > $signed(((^~reg210) ?
                      reg314 : (~^reg763)))) ?
                  reg740 : {reg710, reg253});
            end
          reg839 = $signed(($unsigned((|forvar826[(5'h14):(5'h12)])) ~^ {$unsigned($unsigned((8'ha4))),
              reg135,
              {(wire683 - reg168), (+(7'h48)), reg791}}));
        end
    end
  assign wire840 = reg115[(4'h9):(1'h1)];
  always
    @(posedge clk) begin
      reg841 <= $signed(reg213[(4'hd):(4'hc)]);
    end
  assign wire842 = ($unsigned(((wire241 ^~ wire77[(2'h3):(2'h2)]) ?
                           reg783 : {(reg233 ? reg141 : (7'h49)), (&reg108)})) ?
                       {{((8'hb9) ?
                                   reg194[(3'h6):(2'h2)] : (reg322 >>> (7'h4f))),
                               (reg228 ?
                                   (reg268 ? (8'ha6) : reg158) : {reg206,
                                       reg737,
                                       reg822}),
                               $signed(reg278[(1'h0):(1'h0)])}} : $unsigned(($signed($signed(reg701)) ?
                           reg741[(4'he):(2'h3)] : $unsigned(reg191[(1'h1):(1'h1)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module326
#(parameter param680 = ((((((7'h42) ? (8'ha4) : (7'h57)) ? (~&(7'h41)) : ((8'hb4) >>> (7'h4a))) && {{(8'hbe)}, ((8'hb1) > (7'h4e)), ((8'h9d) ? (7'h42) : (8'hb5))}) - ((&(~&(8'hb7))) >= (7'h4e))) ? (7'h40) : {(!((~(8'haa)) != (7'h47)))}), 
parameter param681 = param680, 
parameter param682 = (param681 & param680))
(y, clk, wire331, wire330, wire329, wire328, wire327);
  output wire [(32'h1673):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire331;
  input wire signed [(5'h1b):(1'h0)] wire330;
  input wire signed [(5'h1f):(1'h0)] wire329;
  input wire [(4'hc):(1'h0)] wire328;
  input wire [(5'h14):(1'h0)] wire327;
  wire [(5'h1d):(1'h0)] wire577;
  wire signed [(2'h2):(1'h0)] wire525;
  wire [(4'ha):(1'h0)] wire469;
  wire signed [(2'h2):(1'h0)] wire447;
  wire [(2'h2):(1'h0)] wire446;
  wire signed [(5'h13):(1'h0)] wire445;
  wire [(5'h1b):(1'h0)] wire420;
  wire [(4'hc):(1'h0)] wire419;
  wire [(4'h9):(1'h0)] wire363;
  wire [(2'h2):(1'h0)] wire335;
  wire signed [(5'h17):(1'h0)] wire334;
  wire [(4'hc):(1'h0)] wire333;
  wire [(2'h3):(1'h0)] wire332;
  reg [(5'h1d):(1'h0)] reg679 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg678 = (1'h0);
  reg [(4'h9):(1'h0)] reg676 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg672 = (1'h0);
  reg [(5'h14):(1'h0)] reg668 = (1'h0);
  reg [(5'h1c):(1'h0)] reg667 = (1'h0);
  reg [(5'h18):(1'h0)] reg665 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg662 = (1'h0);
  reg [(3'h7):(1'h0)] reg658 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg656 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg654 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg653 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg652 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg644 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg643 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg639 = (1'h0);
  reg [(5'h1b):(1'h0)] reg637 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg636 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg635 = (1'h0);
  reg [(5'h17):(1'h0)] reg634 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg633 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg631 = (1'h0);
  reg [(2'h2):(1'h0)] reg629 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg627 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg626 = (1'h0);
  reg [(3'h5):(1'h0)] reg624 = (1'h0);
  reg [(5'h18):(1'h0)] reg622 = (1'h0);
  reg [(5'h10):(1'h0)] reg619 = (1'h0);
  reg [(4'h9):(1'h0)] reg618 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg616 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg614 = (1'h0);
  reg [(5'h16):(1'h0)] reg613 = (1'h0);
  reg [(5'h13):(1'h0)] reg611 = (1'h0);
  reg [(4'hf):(1'h0)] reg610 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg609 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg608 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg607 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg603 = (1'h0);
  reg [(5'h18):(1'h0)] reg602 = (1'h0);
  reg [(4'h8):(1'h0)] reg601 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg598 = (1'h0);
  reg [(4'he):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg590 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg587 = (1'h0);
  reg [(3'h4):(1'h0)] reg586 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg583 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg582 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg575 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg574 = (1'h0);
  reg [(5'h15):(1'h0)] reg573 = (1'h0);
  reg [(3'h7):(1'h0)] reg572 = (1'h0);
  reg [(5'h18):(1'h0)] reg571 = (1'h0);
  reg [(4'hc):(1'h0)] reg568 = (1'h0);
  reg [(4'h8):(1'h0)] reg564 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg563 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg560 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg557 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg554 = (1'h0);
  reg [(5'h12):(1'h0)] reg553 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg549 = (1'h0);
  reg [(5'h17):(1'h0)] reg545 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg543 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg542 = (1'h0);
  reg [(5'h14):(1'h0)] reg539 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg538 = (1'h0);
  reg [(5'h1f):(1'h0)] reg537 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg536 = (1'h0);
  reg [(5'h13):(1'h0)] reg534 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg531 = (1'h0);
  reg [(4'hb):(1'h0)] reg530 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg528 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg524 = (1'h0);
  reg [(4'ha):(1'h0)] reg523 = (1'h0);
  reg [(2'h2):(1'h0)] reg520 = (1'h0);
  reg signed [(4'he):(1'h0)] reg519 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg518 = (1'h0);
  reg [(4'hd):(1'h0)] reg507 = (1'h0);
  reg [(2'h2):(1'h0)] reg505 = (1'h0);
  reg [(4'h9):(1'h0)] reg503 = (1'h0);
  reg [(3'h5):(1'h0)] reg501 = (1'h0);
  reg [(4'hc):(1'h0)] reg494 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg492 = (1'h0);
  reg [(5'h13):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg481 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg477 = (1'h0);
  reg [(5'h15):(1'h0)] reg474 = (1'h0);
  reg [(5'h18):(1'h0)] reg471 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg465 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg462 = (1'h0);
  reg [(4'ha):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg452 = (1'h0);
  reg [(5'h12):(1'h0)] reg448 = (1'h0);
  reg [(5'h1f):(1'h0)] reg441 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg438 = (1'h0);
  reg [(5'h1d):(1'h0)] reg437 = (1'h0);
  reg [(5'h13):(1'h0)] reg436 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg435 = (1'h0);
  reg [(3'h4):(1'h0)] reg434 = (1'h0);
  reg [(5'h17):(1'h0)] reg430 = (1'h0);
  reg [(5'h14):(1'h0)] reg425 = (1'h0);
  reg [(5'h18):(1'h0)] reg421 = (1'h0);
  reg [(5'h1e):(1'h0)] reg418 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg417 = (1'h0);
  reg [(2'h3):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg412 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg411 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg399 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg396 = (1'h0);
  reg [(5'h13):(1'h0)] reg393 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg390 = (1'h0);
  reg [(3'h5):(1'h0)] reg389 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg388 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg386 = (1'h0);
  reg [(5'h1a):(1'h0)] reg383 = (1'h0);
  reg [(5'h16):(1'h0)] reg377 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg376 = (1'h0);
  reg [(3'h5):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg371 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg369 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg361 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg358 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg354 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg351 = (1'h0);
  reg [(5'h1c):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg348 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg343 = (1'h0);
  reg [(3'h4):(1'h0)] reg341 = (1'h0);
  reg [(4'ha):(1'h0)] reg340 = (1'h0);
  reg [(5'h1a):(1'h0)] reg677 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg675 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg674 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg673 = (1'h0);
  reg [(5'h14):(1'h0)] reg671 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar670 = (1'h0);
  reg [(4'h9):(1'h0)] forvar669 = (1'h0);
  reg [(5'h1e):(1'h0)] reg666 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg663 = (1'h0);
  reg [(5'h16):(1'h0)] reg661 = (1'h0);
  reg [(5'h1f):(1'h0)] reg660 = (1'h0);
  reg [(5'h12):(1'h0)] reg659 = (1'h0);
  reg [(4'hc):(1'h0)] reg657 = (1'h0);
  reg [(3'h6):(1'h0)] reg655 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg650 = (1'h0);
  reg [(3'h6):(1'h0)] forvar649 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg648 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg647 = (1'h0);
  reg [(4'hf):(1'h0)] reg646 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg645 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar642 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg641 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar640 = (1'h0);
  reg [(5'h11):(1'h0)] reg638 = (1'h0);
  reg [(5'h10):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg630 = (1'h0);
  reg [(4'hc):(1'h0)] reg628 = (1'h0);
  reg [(3'h4):(1'h0)] reg625 = (1'h0);
  reg [(2'h3):(1'h0)] forvar623 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar621 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg620 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg617 = (1'h0);
  reg [(5'h17):(1'h0)] reg615 = (1'h0);
  reg [(5'h12):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg606 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg605 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg604 = (1'h0);
  reg [(5'h13):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg599 = (1'h0);
  reg [(5'h14):(1'h0)] reg597 = (1'h0);
  reg [(3'h4):(1'h0)] reg596 = (1'h0);
  reg signed [(4'he):(1'h0)] reg594 = (1'h0);
  reg [(4'hb):(1'h0)] reg593 = (1'h0);
  reg [(4'ha):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg591 = (1'h0);
  reg [(5'h19):(1'h0)] reg589 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg588 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg585 = (1'h0);
  reg [(3'h6):(1'h0)] forvar584 = (1'h0);
  reg [(5'h16):(1'h0)] reg581 = (1'h0);
  reg [(5'h14):(1'h0)] reg580 = (1'h0);
  reg [(5'h10):(1'h0)] forvar579 = (1'h0);
  reg [(4'h9):(1'h0)] forvar578 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg576 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar565 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg569 = (1'h0);
  reg [(2'h3):(1'h0)] reg567 = (1'h0);
  reg [(4'h8):(1'h0)] reg566 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg565 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg561 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg555 = (1'h0);
  reg [(5'h13):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg550 = (1'h0);
  reg [(4'hc):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg547 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar546 = (1'h0);
  reg [(5'h15):(1'h0)] reg544 = (1'h0);
  reg [(4'ha):(1'h0)] reg541 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg540 = (1'h0);
  reg [(4'hc):(1'h0)] forvar535 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg533 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg532 = (1'h0);
  reg [(4'ha):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg527 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar526 = (1'h0);
  reg [(5'h1b):(1'h0)] reg522 = (1'h0);
  reg [(5'h10):(1'h0)] reg521 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg513 = (1'h0);
  reg [(4'h8):(1'h0)] forvar512 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg517 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg516 = (1'h0);
  reg [(3'h4):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg514 = (1'h0);
  reg [(3'h4):(1'h0)] forvar513 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg512 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg511 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg510 = (1'h0);
  reg [(3'h5):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg508 = (1'h0);
  reg [(4'hf):(1'h0)] reg506 = (1'h0);
  reg [(2'h2):(1'h0)] reg504 = (1'h0);
  reg [(3'h5):(1'h0)] reg502 = (1'h0);
  reg [(5'h16):(1'h0)] reg500 = (1'h0);
  reg [(5'h1b):(1'h0)] reg499 = (1'h0);
  reg [(4'h9):(1'h0)] reg498 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg497 = (1'h0);
  reg [(4'he):(1'h0)] reg496 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar495 = (1'h0);
  reg [(4'h9):(1'h0)] reg493 = (1'h0);
  reg [(5'h12):(1'h0)] forvar491 = (1'h0);
  reg [(4'hb):(1'h0)] reg490 = (1'h0);
  reg [(4'ha):(1'h0)] reg489 = (1'h0);
  reg [(5'h1d):(1'h0)] reg488 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg487 = (1'h0);
  reg [(3'h4):(1'h0)] reg486 = (1'h0);
  reg [(5'h15):(1'h0)] reg485 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg484 = (1'h0);
  reg [(2'h3):(1'h0)] reg483 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg479 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg476 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg475 = (1'h0);
  reg [(5'h11):(1'h0)] forvar473 = (1'h0);
  reg [(4'hb):(1'h0)] forvar472 = (1'h0);
  reg [(5'h1d):(1'h0)] reg470 = (1'h0);
  reg [(5'h12):(1'h0)] reg468 = (1'h0);
  reg [(4'he):(1'h0)] reg467 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg466 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg464 = (1'h0);
  reg [(5'h1c):(1'h0)] reg454 = (1'h0);
  reg [(5'h1f):(1'h0)] reg450 = (1'h0);
  reg [(5'h12):(1'h0)] forvar449 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg463 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar461 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg460 = (1'h0);
  reg [(3'h6):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg457 = (1'h0);
  reg [(5'h1b):(1'h0)] reg456 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar454 = (1'h0);
  reg [(4'ha):(1'h0)] reg451 = (1'h0);
  reg [(5'h15):(1'h0)] forvar450 = (1'h0);
  reg [(2'h2):(1'h0)] reg449 = (1'h0);
  reg signed [(4'he):(1'h0)] reg444 = (1'h0);
  reg [(3'h5):(1'h0)] reg443 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg440 = (1'h0);
  reg [(5'h16):(1'h0)] reg439 = (1'h0);
  reg [(3'h4):(1'h0)] reg433 = (1'h0);
  reg signed [(4'he):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg431 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg429 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg427 = (1'h0);
  reg [(3'h7):(1'h0)] forvar426 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar424 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg423 = (1'h0);
  reg [(5'h1a):(1'h0)] reg422 = (1'h0);
  reg [(2'h2):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar415 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg414 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg410 = (1'h0);
  reg [(5'h12):(1'h0)] reg409 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg408 = (1'h0);
  reg [(5'h13):(1'h0)] reg407 = (1'h0);
  reg [(4'ha):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg404 = (1'h0);
  reg [(4'hb):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg391 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar385 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg401 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar399 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg397 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg394 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg392 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar391 = (1'h0);
  reg [(5'h17):(1'h0)] reg387 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg385 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg384 = (1'h0);
  reg [(4'hf):(1'h0)] reg382 = (1'h0);
  reg [(4'hd):(1'h0)] reg381 = (1'h0);
  reg [(4'hc):(1'h0)] reg380 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg379 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg378 = (1'h0);
  reg [(4'he):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg373 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg372 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg367 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg366 = (1'h0);
  reg [(3'h7):(1'h0)] forvar365 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar364 = (1'h0);
  reg [(5'h19):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg360 = (1'h0);
  reg [(4'h9):(1'h0)] reg357 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar356 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg355 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg353 = (1'h0);
  reg [(4'hd):(1'h0)] reg352 = (1'h0);
  reg [(5'h1c):(1'h0)] reg350 = (1'h0);
  reg [(5'h1a):(1'h0)] reg347 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg345 = (1'h0);
  reg [(5'h1f):(1'h0)] reg342 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar339 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg338 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar337 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar336 = (1'h0);
  assign y = {wire577,
                 wire525,
                 wire469,
                 wire447,
                 wire446,
                 wire445,
                 wire420,
                 wire419,
                 wire363,
                 wire335,
                 wire334,
                 wire333,
                 wire332,
                 reg679,
                 reg678,
                 reg676,
                 reg672,
                 reg668,
                 reg667,
                 reg665,
                 reg662,
                 reg658,
                 reg656,
                 reg654,
                 reg653,
                 reg652,
                 reg644,
                 reg643,
                 reg639,
                 reg637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 reg631,
                 reg629,
                 reg627,
                 reg626,
                 reg624,
                 reg622,
                 reg619,
                 reg618,
                 reg616,
                 reg614,
                 reg613,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg603,
                 reg602,
                 reg601,
                 reg598,
                 reg595,
                 reg590,
                 reg587,
                 reg586,
                 reg583,
                 reg582,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 reg571,
                 reg568,
                 reg564,
                 reg563,
                 reg560,
                 reg557,
                 reg556,
                 reg554,
                 reg553,
                 reg552,
                 reg549,
                 reg545,
                 reg543,
                 reg542,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 reg534,
                 reg531,
                 reg530,
                 reg528,
                 reg524,
                 reg523,
                 reg520,
                 reg519,
                 reg518,
                 reg507,
                 reg505,
                 reg503,
                 reg501,
                 reg494,
                 reg492,
                 reg482,
                 reg481,
                 reg478,
                 reg477,
                 reg474,
                 reg471,
                 reg465,
                 reg461,
                 reg462,
                 reg458,
                 reg455,
                 reg453,
                 reg452,
                 reg448,
                 reg441,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg430,
                 reg425,
                 reg421,
                 reg418,
                 reg417,
                 reg413,
                 reg412,
                 reg411,
                 reg406,
                 reg403,
                 reg399,
                 reg400,
                 reg398,
                 reg396,
                 reg393,
                 reg390,
                 reg389,
                 reg388,
                 reg386,
                 reg383,
                 reg377,
                 reg376,
                 reg375,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg361,
                 reg359,
                 reg358,
                 reg354,
                 reg351,
                 reg349,
                 reg348,
                 reg344,
                 reg343,
                 reg341,
                 reg340,
                 reg677,
                 reg675,
                 reg674,
                 reg673,
                 reg671,
                 forvar670,
                 forvar669,
                 reg666,
                 reg664,
                 reg663,
                 reg661,
                 reg660,
                 reg659,
                 reg657,
                 reg655,
                 reg651,
                 reg650,
                 forvar649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 forvar642,
                 reg641,
                 forvar640,
                 reg638,
                 reg632,
                 reg630,
                 reg628,
                 reg625,
                 forvar623,
                 forvar621,
                 reg620,
                 reg617,
                 reg615,
                 reg612,
                 reg606,
                 reg605,
                 reg604,
                 reg600,
                 reg599,
                 reg597,
                 reg596,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg589,
                 reg588,
                 reg585,
                 forvar584,
                 reg581,
                 reg580,
                 forvar579,
                 forvar578,
                 reg576,
                 forvar565,
                 reg570,
                 reg569,
                 reg567,
                 reg566,
                 reg565,
                 reg562,
                 reg561,
                 reg559,
                 reg558,
                 reg555,
                 reg551,
                 reg550,
                 reg548,
                 reg547,
                 forvar546,
                 reg544,
                 reg541,
                 reg540,
                 forvar535,
                 reg533,
                 reg532,
                 reg529,
                 reg527,
                 forvar526,
                 reg522,
                 reg521,
                 reg513,
                 forvar512,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 forvar513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg506,
                 reg504,
                 reg502,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 forvar495,
                 reg493,
                 forvar491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg480,
                 reg479,
                 reg476,
                 reg475,
                 forvar473,
                 forvar472,
                 reg470,
                 reg468,
                 reg467,
                 reg466,
                 reg464,
                 reg454,
                 reg450,
                 forvar449,
                 reg463,
                 forvar461,
                 reg460,
                 reg459,
                 reg457,
                 reg456,
                 forvar454,
                 reg451,
                 forvar450,
                 reg449,
                 reg444,
                 reg443,
                 reg442,
                 reg440,
                 reg439,
                 reg433,
                 reg432,
                 reg431,
                 reg429,
                 reg428,
                 reg427,
                 forvar426,
                 forvar424,
                 reg423,
                 reg422,
                 reg416,
                 forvar415,
                 reg414,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg405,
                 reg404,
                 reg402,
                 reg391,
                 forvar385,
                 reg401,
                 forvar399,
                 reg397,
                 reg395,
                 reg394,
                 reg392,
                 forvar391,
                 reg387,
                 reg385,
                 reg384,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg374,
                 reg373,
                 reg372,
                 reg367,
                 reg366,
                 forvar365,
                 forvar364,
                 reg362,
                 reg360,
                 reg357,
                 forvar356,
                 reg355,
                 reg353,
                 reg352,
                 reg350,
                 reg347,
                 reg346,
                 reg345,
                 reg342,
                 forvar339,
                 reg338,
                 forvar337,
                 forvar336,
                 (1'h0)};
  assign wire332 = $unsigned($signed((($unsigned(wire328) ?
                           $signed(wire327) : wire331) ?
                       (^~(8'ha9)) : wire327[(4'h9):(1'h0)])));
  assign wire333 = {((~|wire331[(1'h0):(1'h0)]) ?
                           $signed($unsigned($signed(wire331))) : (8'hb6)),
                       (wire332 << wire328),
                       {(wire327 ? $unsigned($signed(wire331)) : wire331),
                           wire329,
                           ((~((7'h4d) < wire332)) * (wire327 >= (7'h53)))}};
  assign wire334 = $signed($unsigned($unsigned((wire332[(1'h1):(1'h0)] ?
                       wire332 : (wire329 << wire327)))));
  assign wire335 = ($unsigned((~|wire330)) ~^ ($unsigned(wire330[(5'h13):(4'hc)]) >> (~wire327)));
  always
    @(posedge clk) begin
      for (forvar336 = (1'h0); (forvar336 < (2'h2)); forvar336 = (forvar336 + (1'h1)))
        begin
          for (forvar337 = (1'h0); (forvar337 < (2'h3)); forvar337 = (forvar337 + (1'h1)))
            begin
              reg338 = wire327[(1'h0):(1'h0)];
            end
        end
      for (forvar339 = (1'h0); (forvar339 < (1'h1)); forvar339 = (forvar339 + (1'h1)))
        begin
          if ((7'h44))
            begin
              reg340 <= ((~^(wire329 ?
                      ($unsigned((7'h45)) ?
                          $signed(wire331) : (reg338 > (8'h9f))) : (-wire332[(1'h1):(1'h0)]))) ?
                  forvar336[(2'h2):(1'h0)] : (^$unsigned(((&(7'h57)) - {forvar336,
                      wire333}))));
              reg341 <= {(+$signed(($signed(wire334) | reg340[(3'h6):(3'h5)]))),
                  (&$signed((|wire328)))};
              reg342 = wire328;
              reg343 <= wire327[(3'h4):(2'h3)];
              reg344 <= (wire331 * wire334);
              reg345 = $signed(reg342);
            end
          else
            begin
              reg342 = (!reg345);
              reg345 = $signed($unsigned($signed(wire333[(4'hc):(1'h0)])));
            end
          if (forvar339)
            begin
              reg346 = ($signed($signed(reg340[(1'h1):(1'h0)])) ?
                  forvar339[(3'h4):(2'h3)] : wire327[(4'hd):(1'h0)]);
              reg347 = $signed((wire329 ^~ forvar336[(4'hb):(4'ha)]));
              reg348 <= $signed(reg346);
              reg349 <= (!wire332);
              reg350 = wire330[(4'hf):(4'h8)];
            end
          else
            begin
              reg348 <= (~^wire335[(2'h2):(1'h0)]);
              reg350 = $unsigned((~(-(reg343 && (reg346 <= wire332)))));
              reg351 <= reg344;
            end
          if ($signed(reg342))
            begin
              reg352 = wire329[(5'h13):(4'hf)];
              reg353 = $signed(reg346);
              reg354 <= (+reg346[(2'h2):(1'h0)]);
            end
          else
            begin
              reg354 <= $unsigned(forvar339);
              reg355 = (~|reg348);
            end
          for (forvar356 = (1'h0); (forvar356 < (3'h6)); forvar356 = (forvar356 + (1'h1)))
            begin
              reg357 = {$unsigned((reg343[(3'h6):(3'h5)] || (reg345[(5'h16):(5'h12)] >> (reg344 == reg355))))};
              reg358 <= reg355;
              reg359 <= wire333[(1'h0):(1'h0)];
              reg360 = (((~^$signed((wire332 ~^ reg352))) + (~|$signed(((8'hbb) << reg348)))) * ((~|((wire332 | reg342) ?
                  (~wire335) : $signed(forvar339))) == $signed($unsigned(forvar336))));
              reg361 <= reg344;
              reg362 = {({((~reg355) ?
                          (forvar339 << reg355) : $unsigned(wire330)),
                      $unsigned(reg358[(4'hb):(3'h5)])} > forvar356[(1'h0):(1'h0)]),
                  {reg358[(4'h8):(2'h3)]}};
            end
        end
    end
  assign wire363 = $unsigned((({(reg361 <<< wire329),
                           {wire334, reg358},
                           wire331} ?
                       $signed(((7'h53) ?
                           reg348 : reg358)) : ($unsigned(reg358) >> $signed(wire327))) >> reg354));
  always
    @(posedge clk) begin
      for (forvar364 = (1'h0); (forvar364 < (1'h0)); forvar364 = (forvar364 + (1'h1)))
        begin
          for (forvar365 = (1'h0); (forvar365 < (3'h6)); forvar365 = (forvar365 + (1'h1)))
            begin
              reg366 = (8'ha5);
              reg367 = $unsigned($signed({reg351[(5'h1a):(4'hd)]}));
              reg368 <= ({$signed((|$unsigned(wire334)))} && wire328[(1'h1):(1'h0)]);
              reg369 <= (~{($unsigned(reg348) << ($signed(reg358) ?
                      {wire335, reg366} : wire330))});
            end
          if ((~^$unsigned((|((8'h9f) | (wire335 < reg354))))))
            begin
              reg370 <= $unsigned($unsigned(reg340[(1'h0):(1'h0)]));
              reg371 <= $signed($unsigned(((8'ha3) ?
                  (wire363 < $signed(reg359)) : wire330[(4'hf):(3'h5)])));
            end
          else
            begin
              reg372 = (({$signed((7'h57)),
                          (wire333 ? (&reg361) : wire335[(1'h1):(1'h1)])} ?
                      reg354[(3'h5):(1'h1)] : reg344) ?
                  $signed((+$signed(reg371))) : ($unsigned({(^reg343)}) ?
                      ({$unsigned(reg369)} + (~&(wire335 != wire332))) : (~^(~^((7'h4d) && wire333)))));
              reg373 = $unsigned((!(($unsigned(reg351) ?
                  wire334 : reg372[(5'h10):(1'h0)]) * (wire363[(3'h4):(1'h1)] < (wire329 ?
                  reg367 : (7'h43))))));
              reg374 = $signed({$signed($unsigned(wire335)),
                  (wire334[(5'h12):(2'h3)] ?
                      reg368 : ((wire334 & forvar365) ?
                          (^~reg359) : forvar365[(3'h6):(2'h2)])),
                  reg343[(4'ha):(3'h7)]});
              reg375 <= (reg366 ?
                  reg348 : (wire331[(1'h1):(1'h0)] ?
                      $unsigned(((reg368 ? wire333 : wire327) ?
                          (+(7'h40)) : reg341)) : $unsigned($unsigned({wire332,
                          reg366,
                          reg340}))));
              reg376 <= wire333[(1'h1):(1'h1)];
              reg377 <= ((((reg366 ? (~reg376) : reg368) ?
                      reg367 : ({reg373, wire331, reg366} ?
                          {reg359, wire327, wire328} : $unsigned(reg354))) ?
                  ($signed((wire330 ?
                      wire327 : wire328)) ~^ (reg351 >= (reg372 & reg372))) : reg349) >= reg354[(3'h5):(2'h3)]);
            end
          reg378 = reg349[(3'h5):(3'h5)];
          reg379 = $unsigned((8'ha9));
          reg380 = reg367;
          reg381 = (|((^~(wire331[(4'hc):(1'h0)] ?
                  $signed(wire333) : (8'hb6))) ?
              $signed(reg358[(5'h10):(4'h8)]) : (wire335[(1'h1):(1'h0)] ^~ wire332[(2'h3):(2'h3)])));
          reg382 = $signed($unsigned($unsigned($signed(wire329))));
        end
      reg383 <= $unsigned($signed({(^~(-reg373))}));
      reg384 = ((!((!(|reg381)) ?
          $signed({reg372, wire334}) : reg340)) ~^ $signed($signed((reg344 ?
          {reg378, reg358} : $signed(reg366)))));
      if (wire330[(1'h0):(1'h0)])
        begin
          reg385 = (&((|(^reg374)) ?
              $signed(wire333[(1'h1):(1'h1)]) : (~&forvar364[(3'h5):(2'h3)])));
          if ((8'ha1))
            begin
              reg386 <= reg381[(2'h2):(2'h2)];
              reg387 = (!(reg366[(2'h3):(1'h0)] ~^ $signed(reg377[(4'hb):(1'h1)])));
              reg388 <= $unsigned($signed($unsigned((reg376 * $signed(wire363)))));
              reg389 <= ($signed($signed(wire329[(4'he):(1'h0)])) | (!(+$unsigned(reg343[(5'h14):(4'hf)]))));
              reg390 <= (^reg389);
            end
          else
            begin
              reg387 = (~|$unsigned($unsigned(($signed(wire331) ?
                  $signed(reg385) : (&wire333)))));
              reg388 <= (|reg358[(2'h2):(2'h2)]);
            end
          for (forvar391 = (1'h0); (forvar391 < (2'h2)); forvar391 = (forvar391 + (1'h1)))
            begin
              reg392 = $unsigned((reg373[(5'h16):(4'hf)] ?
                  $signed((reg348 <= (~&wire331))) : (|$signed(reg382))));
              reg393 <= ($unsigned($unsigned(reg340)) ?
                  ((7'h49) ?
                      $unsigned((wire330[(5'h1a):(4'hb)] <= reg344)) : $unsigned($signed((!wire329)))) : $signed((-$unsigned($unsigned(reg343)))));
              reg394 = reg343[(4'h8):(4'h8)];
              reg395 = (reg351 ?
                  $signed((({reg386} ?
                      reg373 : (reg387 < reg349)) * $signed((!reg379)))) : (($unsigned(((7'h46) ?
                      reg372 : forvar391)) < ((reg379 >>> reg392) ~^ ((8'haf) ?
                      reg393 : reg377))) > reg351[(3'h4):(2'h2)]));
              reg396 <= ($unsigned(wire363[(3'h6):(3'h4)]) ^ $unsigned(wire333[(4'h9):(3'h5)]));
              reg397 = ((reg393 ?
                  (~$unsigned($signed(reg361))) : $unsigned($unsigned(((7'h49) ?
                      reg369 : wire328)))) << reg396);
            end
          reg398 <= $signed({reg349,
              $unsigned($unsigned((reg361 || reg379))),
              wire329[(4'he):(3'h7)]});
          for (forvar399 = (1'h0); (forvar399 < (1'h0)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg400 <= (reg370 | $signed(wire327[(3'h4):(3'h4)]));
            end
          reg401 = reg389[(1'h0):(1'h0)];
        end
      else
        begin
          for (forvar385 = (1'h0); (forvar385 < (2'h2)); forvar385 = (forvar385 + (1'h1)))
            begin
              reg387 = reg397[(2'h2):(2'h2)];
              reg388 <= (~&(~^$unsigned((~&(wire328 ? (8'hab) : (8'hb2))))));
              reg391 = (&(((+{wire335, reg351, reg371}) ?
                  $unsigned(reg348) : (wire333 ?
                      $signed((8'ha2)) : (&reg361))) == $signed(((^~(8'hbc)) ?
                  reg377 : $signed(reg392)))));
              reg393 <= (~&$unsigned({((wire331 ? (7'h4f) : reg361) ?
                      $unsigned(reg386) : {reg367, reg380, reg390})}));
              reg394 = ($unsigned((~^(reg386 ?
                      reg398[(4'ha):(1'h1)] : forvar364[(2'h2):(1'h1)]))) ?
                  reg361 : ({wire333} ?
                      $signed(reg359[(5'h10):(3'h4)]) : $signed(reg387)));
              reg396 <= (reg391 ?
                  ($unsigned($signed((forvar391 > (8'hb4)))) ?
                      ((&{reg380, reg340}) ?
                          $signed(((8'hb2) ?
                              wire331 : forvar399)) : reg349[(2'h2):(2'h2)]) : (!(|reg374))) : wire331);
              reg398 <= reg382[(4'he):(3'h7)];
            end
          if (((reg401[(4'hc):(4'h8)] ?
              (((wire363 ^ (8'hbd)) ?
                  (7'h50) : $signed((7'h54))) + wire331[(3'h4):(3'h4)]) : ($unsigned((forvar385 ?
                      (8'hbc) : reg400)) ?
                  (forvar391 ? $unsigned(wire329) : reg370) : ((!reg398) ?
                      $signed(reg354) : reg371))) <= $unsigned(((~&(-reg387)) ?
              reg349[(5'h1a):(3'h4)] : $unsigned((reg349 ? reg396 : reg390))))))
            begin
              reg399 <= (((($unsigned(reg351) ?
                      ((8'hab) & (8'ha0)) : $unsigned((8'hb5))) ?
                  $unsigned($signed(reg398)) : (((7'h56) && reg343) ?
                      $unsigned(wire331) : $unsigned(reg340))) < reg385[(5'h18):(2'h2)]) ^ (+{reg400,
                  $unsigned(reg401[(4'hd):(2'h3)])}));
              reg401 = reg385;
              reg402 = (~(^(-{(reg396 <<< reg377)})));
              reg403 <= (((+reg393[(4'hf):(1'h0)]) ?
                  (($unsigned(reg369) ?
                      wire335[(1'h1):(1'h0)] : reg381[(1'h0):(1'h0)]) ~^ wire363[(3'h6):(3'h6)]) : (^~$unsigned($unsigned((7'h52))))) != ((($unsigned(wire331) || (reg376 ?
                          reg376 : (8'hb5))) ?
                      (-{(7'h57), (7'h4f)}) : {((7'h4b) ? (8'hb1) : wire335),
                          reg380}) ?
                  $signed((~|reg341)) : ($signed($signed(reg367)) ^ ((reg396 ?
                          wire329 : reg393) ?
                      {reg368, reg372} : wire327))));
            end
          else
            begin
              reg399 <= {reg394};
              reg401 = $unsigned((-(!reg378)));
            end
          reg404 = $signed(reg403);
          if ((!$signed(({{forvar364, wire331}, (reg398 ? reg372 : reg388)} ?
              (8'hac) : $signed(reg378)))))
            begin
              reg405 = (reg344 ? $unsigned((8'ha2)) : reg398[(5'h10):(3'h7)]);
              reg406 <= (^~reg378);
              reg407 = ((reg383 >= ((^wire331[(3'h6):(2'h3)]) ?
                      $signed(reg378) : (~|$unsigned(reg370)))) ?
                  reg340[(1'h0):(1'h0)] : ((|($unsigned((8'hb3)) ~^ reg343[(5'h15):(4'h8)])) ?
                      reg385 : reg400[(3'h4):(1'h1)]));
              reg408 = ($signed($unsigned({reg382,
                  (^~reg394)})) || $unsigned(((~|(^~reg391)) ?
                  reg366 : $unsigned(wire332[(2'h3):(2'h2)]))));
              reg409 = wire333;
              reg410 = $unsigned((forvar365 ?
                  $unsigned(reg390[(3'h5):(2'h2)]) : (-(reg403[(1'h1):(1'h0)] ?
                      {reg405} : (reg387 ? wire330 : (8'hac))))));
            end
          else
            begin
              reg405 = ((reg375[(3'h4):(3'h4)] ~^ reg395) ?
                  wire333[(4'h8):(3'h5)] : $unsigned((!{(!reg366)})));
              reg406 <= ((|($unsigned((reg389 ? reg371 : (8'had))) ?
                      reg404 : (~^$signed(reg404)))) ?
                  (({(reg370 != (8'ha0)),
                          wire335[(1'h0):(1'h0)]} > $unsigned($signed(reg401))) ?
                      forvar385[(2'h2):(1'h0)] : ((forvar399[(4'h8):(1'h0)] ?
                          reg359 : ((8'hbc) >>> reg381)) <<< (&$signed(reg366)))) : $unsigned(wire363));
              reg407 = ((wire363 | reg370) ?
                  (reg375[(3'h4):(1'h0)] != (reg393 & reg391)) : ({$signed($signed(reg386)),
                          (^~(reg392 ? reg393 : reg351))} ?
                      reg399[(4'hf):(3'h4)] : ($signed($unsigned(reg385)) ?
                          (+(~|reg389)) : ((reg368 || reg387) ~^ (^reg361)))));
              reg408 = (reg387 ?
                  $unsigned(forvar385[(1'h1):(1'h1)]) : ($signed($signed($unsigned(reg401))) >= (((reg401 ?
                          reg402 : reg395) ?
                      reg397 : $unsigned((8'hac))) & $signed((reg375 ?
                      wire335 : reg373)))));
              reg409 = (-(($signed((~^reg344)) ?
                      {(reg408 ? reg351 : reg384),
                          $unsigned(reg361)} : reg391) ?
                  ((~|reg383) ~^ reg376[(2'h2):(1'h1)]) : reg410));
              reg411 <= $unsigned(((7'h51) ?
                  (8'ha5) : ($signed((reg391 ? reg368 : reg396)) ?
                      (^reg379) : $unsigned(((8'hae) ? reg408 : wire363)))));
              reg412 <= wire334[(3'h6):(3'h4)];
            end
          reg413 <= (+reg341);
          reg414 = reg408;
          for (forvar415 = (1'h0); (forvar415 < (1'h0)); forvar415 = (forvar415 + (1'h1)))
            begin
              reg416 = $unsigned({$unsigned(reg374),
                  $unsigned($unsigned((reg374 & reg397))),
                  wire331[(4'h9):(3'h4)]});
              reg417 <= $unsigned($signed((|$unsigned((wire329 < wire363)))));
            end
        end
      reg418 <= {((|reg401[(3'h7):(3'h5)]) ?
              (~&$unsigned({reg344})) : (~&(((8'h9e) >= wire327) * reg388))),
          {$unsigned({reg378, $signed(reg408), ((8'ha2) ? (7'h53) : reg375)}),
              $unsigned(reg394[(4'he):(4'hb)])},
          (^~$signed(((~reg340) ? (~|(7'h44)) : $signed(wire331))))};
    end
  assign wire419 = ((~&$unsigned((&{wire328}))) > ($unsigned((~&$unsigned(reg403))) ?
                       reg358[(5'h1c):(5'h10)] : reg349[(5'h15):(2'h2)]));
  assign wire420 = (8'hb0);
  always
    @(posedge clk) begin
      reg421 <= (reg341 ? reg400 : reg358);
      reg422 = (wire331[(3'h4):(3'h4)] ?
          $unsigned(({$unsigned(reg361)} ?
              $signed($unsigned(reg376)) : $unsigned((reg341 < reg341)))) : $signed($unsigned($signed((reg390 | reg393)))));
      reg423 = (-(reg421 || (((^wire334) ?
          ((8'hb3) ?
              reg403 : wire332) : {reg413}) < $signed($signed((8'hab))))));
    end
  always
    @(posedge clk) begin
      for (forvar424 = (1'h0); (forvar424 < (3'h5)); forvar424 = (forvar424 + (1'h1)))
        begin
          reg425 <= $unsigned((($signed((reg377 ^ (8'hbd))) >> forvar424) << reg389));
          for (forvar426 = (1'h0); (forvar426 < (2'h3)); forvar426 = (forvar426 + (1'h1)))
            begin
              reg427 = reg396;
              reg428 = reg361[(4'he):(4'he)];
              reg429 = $signed(forvar426);
              reg430 <= reg398;
              reg431 = $unsigned($signed({wire419, reg383}));
              reg432 = (|(^$unsigned(reg396[(5'h11):(2'h3)])));
              reg433 = reg432;
            end
          if ({(^~$signed((8'hab)))})
            begin
              reg434 <= {{$signed(((reg348 ? wire332 : reg389) != (-reg340)))},
                  ({wire328[(4'hb):(2'h2)],
                          ((reg411 ?
                              wire363 : reg344) | reg432[(3'h6):(1'h1)])} ?
                      $signed($signed($unsigned(reg354))) : $unsigned(reg396[(3'h6):(3'h6)])),
                  (((reg403[(5'h10):(3'h4)] & reg343[(3'h6):(2'h3)]) ^ $unsigned({reg399})) <<< reg376)};
              reg435 <= (((reg421 ?
                  ({(7'h54), wire332} ?
                      $unsigned(reg399) : (!reg403)) : (~|(reg368 ?
                      reg388 : reg434))) - ((+reg358) >> $signed(reg430[(4'hd):(4'hd)]))) - (7'h54));
              reg436 <= (-reg354[(3'h5):(1'h0)]);
              reg437 <= $signed(reg370);
              reg438 <= reg361;
            end
          else
            begin
              reg439 = (~&(($unsigned(wire329[(5'h19):(4'hc)]) << $unsigned($signed(reg403))) ?
                  ({reg425[(3'h7):(1'h0)], reg398, (reg358 < reg371)} ?
                      reg425 : reg348[(3'h4):(2'h3)]) : $signed((((8'hb7) ?
                      reg386 : reg398) && reg371))));
            end
          reg440 = $signed(wire333[(4'hc):(4'ha)]);
          reg441 <= ((^~reg435[(1'h1):(1'h0)]) << (reg358 ?
              wire363 : wire332[(2'h3):(1'h1)]));
        end
      reg442 = (((^(wire363[(1'h1):(1'h1)] - wire419)) && (~($signed(wire334) ?
              reg377 : $signed(reg375)))) ?
          ((($unsigned(reg431) ?
                  (wire334 ? reg369 : reg351) : $unsigned((7'h58))) ?
              reg358[(4'hf):(4'h9)] : $unsigned((reg430 ?
                  reg369 : wire330))) > ($signed((7'h57)) ?
              (reg377 <= reg340) : reg437)) : $unsigned($unsigned($unsigned((+reg434)))));
      reg443 = (reg390 >>> reg389);
      reg444 = ($unsigned({(&(reg348 ?
              (8'hbe) : forvar426))}) != $signed((^~(~|(|reg375)))));
    end
  assign wire445 = $signed((wire419 ~^ reg437[(5'h16):(5'h14)]));
  assign wire446 = $unsigned(reg343);
  assign wire447 = {wire446[(1'h1):(1'h1)],
                       (^wire327[(5'h11):(2'h3)]),
                       $signed((~$signed((reg438 ^~ wire363))))};
  always
    @(posedge clk) begin
      reg448 <= $signed($signed($unsigned((&wire334[(4'h8):(3'h7)]))));
    end
  always
    @(posedge clk) begin
      if (({$unsigned($unsigned((~|reg441)))} ?
          (&(($signed(reg398) | $signed(reg358)) ?
              ($signed((7'h52)) | (reg448 ?
                  reg343 : wire447)) : (|$signed(reg417)))) : reg437[(5'h16):(3'h6)]))
        begin
          reg449 = (7'h48);
          for (forvar450 = (1'h0); (forvar450 < (1'h0)); forvar450 = (forvar450 + (1'h1)))
            begin
              reg451 = $signed($unsigned($unsigned({(reg425 != wire334)})));
            end
          reg452 <= $unsigned(($signed(reg425[(1'h0):(1'h0)]) ?
              ($unsigned(reg344[(5'h15):(2'h3)]) || {$unsigned(reg343),
                  $unsigned((7'h41))}) : $signed($unsigned($unsigned(reg418)))));
          reg453 <= reg398;
          for (forvar454 = (1'h0); (forvar454 < (1'h1)); forvar454 = (forvar454 + (1'h1)))
            begin
              reg455 <= reg358[(5'h10):(3'h7)];
              reg456 = (+($unsigned(((~reg436) || $unsigned(reg441))) ^ (reg430 != ((7'h52) > $signed(reg389)))));
              reg457 = $signed({reg389[(2'h3):(2'h2)],
                  ((+$unsigned(reg354)) ?
                      ((~^reg386) ?
                          (reg425 ?
                              wire445 : reg453) : wire363[(2'h3):(2'h3)]) : (reg449 ?
                          $unsigned(reg400) : $signed(reg344)))});
              reg458 <= wire446;
              reg459 = $signed(($unsigned((((8'hb4) - reg400) <<< reg348[(3'h4):(1'h1)])) ?
                  (+(8'ha1)) : wire419));
            end
          if ((($unsigned((reg448[(2'h3):(2'h3)] && reg455[(2'h2):(1'h1)])) ?
              (^(reg343[(3'h7):(2'h3)] ?
                  $unsigned((8'hbc)) : wire327)) : ($signed((wire330 ?
                      reg406 : reg437)) ?
                  {(wire332 > wire420)} : $signed($unsigned(wire333)))) * $signed({(reg388[(2'h2):(1'h1)] ?
                  (-reg456) : $unsigned(reg400)),
              $signed((reg441 ? reg403 : reg458)),
              $signed(reg393[(3'h7):(3'h6)])})))
            begin
              reg460 = reg388[(1'h0):(1'h0)];
            end
          else
            begin
              reg460 = $signed($unsigned(reg412));
            end
          for (forvar461 = (1'h0); (forvar461 < (3'h5)); forvar461 = (forvar461 + (1'h1)))
            begin
              reg462 <= ($signed((-({reg458, reg396} ?
                      wire329[(4'h8):(1'h0)] : $unsigned(reg435)))) ?
                  wire334 : ($unsigned(reg458) ?
                      reg386[(2'h2):(2'h2)] : (({reg399} ?
                          $signed((8'hb1)) : (~&reg403)) * ((reg398 ?
                              reg389 : reg434) ?
                          wire447 : (~reg437)))));
              reg463 = reg383[(5'h14):(4'he)];
            end
        end
      else
        begin
          for (forvar449 = (1'h0); (forvar449 < (3'h4)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg450 = {(wire329 ?
                      $signed($unsigned($unsigned(reg354))) : reg383[(4'ha):(1'h1)]),
                  (8'hb5)};
              reg451 = reg358;
              reg452 <= reg411;
              reg453 <= (|$unsigned($signed((+{reg396, reg393, reg354}))));
              reg454 = ((^(^((reg388 ^~ forvar449) < $unsigned((8'hb0))))) ?
                  $unsigned(reg359) : forvar449[(2'h3):(1'h1)]);
              reg456 = (7'h51);
            end
          if (wire446[(1'h1):(1'h0)])
            begin
              reg458 <= ($unsigned({wire327[(4'hd):(2'h2)],
                  reg390}) & $unsigned((~|$signed((reg369 ?
                  reg458 : reg411)))));
              reg459 = reg359[(4'he):(3'h5)];
            end
          else
            begin
              reg458 <= (((((reg449 ? reg396 : reg430) >>> (reg430 ?
                          wire445 : wire419)) ?
                      ((^reg361) > (-(7'h46))) : reg459) << ((~reg398[(4'h8):(4'h8)]) ?
                      $unsigned(reg361[(3'h6):(2'h3)]) : (wire420[(5'h17):(5'h16)] ?
                          reg457 : (reg458 != (8'h9c))))) ?
                  (reg441[(4'h9):(1'h0)] ?
                      $unsigned($unsigned($unsigned(reg383))) : (~&reg376[(3'h6):(2'h3)])) : $unsigned(reg375[(3'h5):(1'h0)]));
              reg461 <= {$signed(($unsigned(((8'had) ? reg437 : (8'hba))) ?
                      (reg412 ?
                          (+reg343) : (reg354 >> (7'h53))) : {$signed(reg359)}))};
              reg463 = (({(reg399[(4'he):(3'h4)] == (reg349 ?
                      reg375 : (7'h56)))} ^ ((~|$unsigned((8'hab))) + $signed($unsigned(reg376)))) <<< ((reg456 ?
                      reg406 : (~^reg452)) ?
                  (8'haa) : $signed(reg358)));
              reg464 = (8'h9e);
              reg465 <= (reg399[(5'h14):(3'h6)] >= (^~{$unsigned(((8'hab) == reg453)),
                  $signed($unsigned(reg441)),
                  reg389}));
              reg466 = ($unsigned($unsigned((forvar449 ?
                  (reg455 ?
                      reg463 : (7'h49)) : (~|reg456)))) | (reg438[(4'h9):(4'h8)] > $unsigned((^~(reg406 ?
                  (8'haf) : reg437)))));
            end
        end
      reg467 = $signed(($unsigned((8'ha7)) ?
          (reg466 ?
              ((~|reg457) <= (~reg411)) : {reg435,
                  (wire446 ? reg435 : reg462)}) : (reg400[(1'h1):(1'h1)] ?
              (reg403[(5'h12):(4'he)] > wire419[(4'h9):(1'h1)]) : (reg435 ~^ $unsigned(reg371)))));
      reg468 = {(($signed((forvar461 != reg421)) | {reg396[(4'hb):(3'h6)],
                  forvar449}) ?
              $unsigned(wire333[(3'h4):(2'h3)]) : wire419[(4'h8):(3'h4)]),
          (reg466[(5'h13):(4'h8)] | (((^~(8'ha3)) ?
                  reg375[(3'h4):(3'h4)] : $unsigned(reg359)) ?
              (((8'hb9) << (8'ha0)) || $unsigned(wire446)) : {(wire327 ?
                      reg437 : wire419)})),
          $unsigned($signed(reg435))};
    end
  assign wire469 = (7'h4b);
  always
    @(posedge clk) begin
      reg470 = ((($unsigned($unsigned(reg340)) ?
          reg349 : (~$unsigned(reg458))) - reg465) >> $unsigned(reg418[(1'h1):(1'h1)]));
      reg471 <= (&$signed(wire445[(5'h12):(5'h12)]));
      for (forvar472 = (1'h0); (forvar472 < (1'h0)); forvar472 = (forvar472 + (1'h1)))
        begin
          for (forvar473 = (1'h0); (forvar473 < (1'h1)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 <= reg448[(4'ha):(3'h7)];
              reg475 = reg441;
              reg476 = (reg430[(5'h17):(2'h2)] || {($unsigned(reg448[(3'h7):(2'h2)]) - ($signed((8'hae)) + wire419[(1'h0):(1'h0)]))});
              reg477 <= $unsigned(reg368[(5'h16):(4'he)]);
              reg478 <= (($unsigned(((reg403 ^~ reg368) ?
                  (~reg371) : $unsigned(reg465))) | {(reg354[(2'h3):(1'h0)] ?
                      forvar472[(3'h5):(3'h4)] : $signed(reg475))}) << (($signed(reg411) ?
                      $signed(reg406[(4'hb):(4'ha)]) : {(reg438 ~^ reg343)}) ?
                  {reg471, $signed($unsigned(reg438))} : reg458));
            end
          reg479 = (((7'h52) << ($signed((wire331 <= reg453)) > reg461[(4'h8):(3'h5)])) ?
              {$unsigned({$signed(reg458),
                      (~^reg438)})} : $unsigned({(^$unsigned(forvar473)),
                  (((8'ha9) ? reg377 : (8'ha7)) << (~&reg476))}));
          reg480 = (-(~(~&$unsigned(reg376))));
          if ((wire331[(4'hb):(1'h1)] ?
              reg413 : $signed($signed({$signed(reg343)}))))
            begin
              reg481 <= {(|$unsigned((reg389 ?
                      ((8'hbf) - (8'haa)) : {reg369, reg349, wire334}))),
                  ({reg461} << (reg386 >>> $signed((reg477 ?
                      reg376 : reg386))))};
              reg482 <= ($signed($signed(($unsigned(reg412) == (+reg453)))) ?
                  $unsigned((^$signed($signed(reg393)))) : $signed((reg413 ?
                      {(^~reg359), (reg361 > reg471)} : wire335)));
              reg483 = $signed((&$signed(reg344)));
            end
          else
            begin
              reg483 = wire420;
              reg484 = (({$signed((reg470 ? reg375 : (8'ha4))),
                          reg348[(1'h0):(1'h0)]} ?
                      ($unsigned({wire332, wire419, reg448}) ?
                          $unsigned((reg349 ?
                              reg399 : reg383)) : wire329) : wire447[(2'h2):(1'h1)]) ?
                  $signed((|reg343[(4'ha):(3'h4)])) : ($signed((reg370 ?
                          wire469[(4'h8):(3'h5)] : (reg340 ?
                              reg393 : reg480))) ?
                      (reg438 | ((~&wire332) ?
                          (^wire363) : reg377[(5'h10):(4'hf)])) : (reg403 ?
                          (^(reg413 ? wire446 : (7'h4a))) : reg483)));
              reg485 = {$signed((8'hac)),
                  (reg361 ? reg418[(5'h13):(3'h4)] : reg483[(2'h2):(2'h2)])};
              reg486 = reg389[(3'h4):(2'h2)];
              reg487 = $signed(($unsigned(wire363[(1'h0):(1'h0)]) ?
                  $unsigned($unsigned((reg413 != wire420))) : reg361));
              reg488 = reg471;
            end
          reg489 = (~&(reg349 ? reg351 : $signed((~&$signed(reg396)))));
          reg490 = wire329;
          for (forvar491 = (1'h0); (forvar491 < (1'h0)); forvar491 = (forvar491 + (1'h1)))
            begin
              reg492 <= (8'hb2);
              reg493 = $signed(($signed((~|{reg430,
                  reg375})) + ($unsigned(reg490[(3'h7):(2'h2)]) ?
                  ($signed(reg351) <<< $signed(reg482)) : $signed((+reg349)))));
            end
        end
      reg494 <= $signed({wire327[(3'h5):(1'h1)]});
      for (forvar495 = (1'h0); (forvar495 < (2'h2)); forvar495 = (forvar495 + (1'h1)))
        begin
          if ((reg418[(5'h12):(5'h11)] + {{($unsigned(reg351) * $signed(wire446)),
                  (^~reg488[(3'h6):(3'h6)]),
                  (|$signed(reg417))}}))
            begin
              reg496 = $unsigned((~|$unsigned($unsigned($signed(wire332)))));
            end
          else
            begin
              reg496 = (+(reg489 > $unsigned((reg396[(5'h15):(3'h4)] ?
                  $unsigned(reg421) : $unsigned(reg436)))));
              reg497 = ({$unsigned($signed(reg375)),
                  ($signed(reg359[(5'h16):(3'h5)]) ?
                      ($signed(reg477) ^ reg492) : reg461)} * {reg383[(1'h0):(1'h0)],
                  (reg483[(1'h0):(1'h0)] ?
                      (~|reg477) : $signed($signed((8'hb3))))});
              reg498 = $signed(reg421[(2'h3):(2'h2)]);
              reg499 = $unsigned((7'h42));
              reg500 = (7'h53);
              reg501 <= $signed($unsigned(reg375[(3'h4):(3'h4)]));
            end
          if ($unsigned($signed($signed(({(7'h53)} ? reg417 : reg452)))))
            begin
              reg502 = $unsigned(((~(reg475 < $unsigned((8'ha1)))) & $unsigned($unsigned(reg477[(3'h6):(2'h3)]))));
              reg503 <= $signed({(7'h42)});
              reg504 = $unsigned((wire332 ?
                  reg453[(3'h6):(3'h6)] : ($unsigned($unsigned(reg340)) >> (wire332[(1'h1):(1'h0)] <= $signed(reg403)))));
              reg505 <= ((7'h42) - (^(^~forvar472[(4'h9):(4'h9)])));
              reg506 = (-((~|$signed((8'h9f))) ?
                  reg493 : $signed($signed(((7'h4e) ? reg376 : reg462)))));
              reg507 <= (reg441 << $unsigned((!((reg455 <= (8'ha0)) ^ {reg421}))));
              reg508 = {(~|((reg489[(3'h4):(1'h0)] == reg489[(3'h4):(2'h2)]) <= (reg489[(3'h4):(2'h2)] >>> (reg358 >>> reg497)))),
                  reg344[(5'h19):(5'h19)],
                  (reg421 >= reg502)};
            end
          else
            begin
              reg503 <= $signed(((reg485[(3'h4):(2'h3)] ?
                      $signed(reg475) : ((reg488 ? reg488 : reg485) ?
                          {(8'hb2), reg430, reg470} : (!wire330))) ?
                  {$signed(((7'h55) - reg388)),
                      (((8'ha9) && reg351) ? reg341 : (^reg413)),
                      $signed($unsigned(reg369))} : $unsigned($signed((reg369 - reg359)))));
            end
          reg509 = reg403[(5'h11):(4'h9)];
          reg510 = ({$unsigned(reg501),
              reg488[(4'ha):(2'h2)],
              reg494[(4'hc):(1'h1)]} ^ (8'hbb));
        end
      if ({reg369,
          reg476,
          (reg351 * (|($unsigned(reg358) ?
              (reg490 ? reg458 : reg461) : $signed(reg498))))})
        begin
          reg511 = (|reg341);
          reg512 = $signed(({(!{reg480, reg437}),
              (reg411[(3'h4):(1'h1)] - (reg358 ? reg412 : reg471))} * reg500));
          for (forvar513 = (1'h0); (forvar513 < (1'h0)); forvar513 = (forvar513 + (1'h1)))
            begin
              reg514 = (^forvar513);
            end
          reg515 = (!{$signed(((reg399 != reg503) ?
                  $unsigned(reg396) : wire469))});
          if (($signed({(^reg412[(5'h17):(4'he)])}) ?
              ($signed({(reg508 ? reg497 : reg480),
                  (reg436 ? (8'ha8) : reg370),
                  reg354}) < (~|reg341)) : ((reg348 ?
                      (~|$unsigned(reg354)) : $unsigned(reg448)) ?
                  $unsigned($signed(reg398)) : $unsigned(reg500))))
            begin
              reg516 = (reg344[(5'h15):(5'h13)] ?
                  {reg361[(4'h8):(1'h1)],
                      wire333[(3'h4):(3'h4)]} : $signed(($unsigned(reg400) * (reg425[(1'h0):(1'h0)] ?
                      {wire446} : {reg486, reg389}))));
              reg517 = (!reg359);
              reg518 <= ((!$signed((+(!reg502)))) ?
                  $signed(reg500[(4'hf):(3'h5)]) : {forvar491,
                      reg515[(2'h3):(2'h2)],
                      $unsigned((|$unsigned(reg461)))});
            end
          else
            begin
              reg516 = reg371;
            end
        end
      else
        begin
          reg511 = ($unsigned((reg487[(2'h2):(1'h1)] > (!$signed(reg388)))) ?
              ((^$unsigned((~^(8'hb8)))) ?
                  (~^((reg458 + reg507) == reg441[(5'h1e):(1'h0)])) : (-(reg341[(1'h0):(1'h0)] && (forvar472 ?
                      reg461 : reg448)))) : $unsigned($unsigned(reg484)));
          for (forvar512 = (1'h0); (forvar512 < (3'h5)); forvar512 = (forvar512 + (1'h1)))
            begin
              reg513 = wire445[(5'h11):(4'he)];
              reg514 = $signed(($signed(reg512) == reg358[(5'h16):(1'h1)]));
            end
          reg518 <= ($unsigned(reg349[(5'h11):(4'ha)]) ?
              reg418 : (-reg511[(2'h2):(1'h1)]));
          reg519 <= reg461;
          reg520 <= (($signed($unsigned((reg487 ^ reg437))) | $signed((7'h45))) ?
              reg506[(4'hc):(3'h4)] : reg488[(4'he):(1'h0)]);
        end
      reg521 = forvar513[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg522 = (((reg406[(5'h1b):(4'h8)] ~^ (~&$unsigned(wire332))) && (wire445 && reg441[(5'h11):(5'h10)])) * reg383);
      reg523 <= $unsigned(({({wire328, reg368} ?
              $signed((7'h56)) : $signed(wire334)),
          $signed($unsigned(reg417)),
          {{reg507, (8'haf)}}} ^~ {(~$unsigned(reg417)),
          ((8'hb4) == ((8'ha4) ? wire335 : reg461))}));
      reg524 <= $unsigned((($signed(reg503) ^ ((reg376 ?
              (8'hbd) : reg377) | wire447)) ?
          ((~|reg399) && wire328) : reg421[(2'h3):(2'h2)]));
    end
  assign wire525 = (^~{$unsigned((wire447[(1'h0):(1'h0)] + (reg412 ?
                           reg377 : (7'h44)))),
                       {reg400[(4'h9):(1'h0)], {reg519}}});
  always
    @(posedge clk) begin
      for (forvar526 = (1'h0); (forvar526 < (3'h4)); forvar526 = (forvar526 + (1'h1)))
        begin
          reg527 = reg377;
          if ({($signed(reg341[(1'h1):(1'h0)]) & reg465[(1'h1):(1'h1)])})
            begin
              reg528 <= ({reg393[(3'h7):(3'h5)]} && (({(-reg413)} ?
                      $unsigned(reg435[(2'h2):(2'h2)]) : wire328[(3'h7):(3'h5)]) ?
                  $unsigned(wire419) : (($unsigned(reg361) || {reg425,
                      reg471,
                      reg351}) - reg383[(5'h17):(2'h3)])));
              reg529 = $signed((({reg430, $unsigned(wire419), (-(7'h44))} ?
                  (((7'h47) >> (8'hab)) >>> (reg361 << reg520)) : (~(reg351 >>> reg471))) ~^ (((reg343 ?
                  wire335 : reg400) ~^ $unsigned(reg471)) < (7'h4e))));
              reg530 <= $signed(reg393);
              reg531 <= $signed(reg441[(5'h18):(3'h6)]);
              reg532 = $signed((($unsigned((~&reg436)) + $unsigned(forvar526[(3'h7):(1'h0)])) >>> (($signed(forvar526) >= (wire469 <<< reg412)) ?
                  (((8'hb1) ?
                      reg399 : (7'h57)) | ((7'h44) ^~ reg399)) : reg465)));
              reg533 = $unsigned({(reg494 ?
                      ((reg400 == reg340) ?
                          $signed(wire329) : reg455) : reg354[(2'h3):(1'h1)]),
                  (reg474[(4'ha):(4'h9)] ?
                      ((~^reg524) + $unsigned(reg376)) : {$unsigned(reg494)}),
                  $unsigned((+(reg390 ? wire334 : reg340)))});
            end
          else
            begin
              reg528 <= wire335;
              reg530 <= ((^($signed($signed(reg390)) >> reg393[(2'h2):(1'h0)])) ?
                  (~|$signed({(reg388 ?
                          reg340 : reg529)})) : $unsigned($unsigned(forvar526[(4'ha):(3'h7)])));
              reg532 = reg354;
              reg534 <= reg399[(2'h3):(1'h0)];
            end
          for (forvar535 = (1'h0); (forvar535 < (1'h0)); forvar535 = (forvar535 + (1'h1)))
            begin
              reg536 <= reg377;
            end
          reg537 <= reg435[(2'h2):(2'h2)];
          if ({wire363,
              ((!(((8'hbf) ? wire328 : reg533) >>> $unsigned((7'h41)))) ?
                  reg376 : wire330[(4'h9):(3'h5)]),
              reg403})
            begin
              reg538 <= (reg398 ? $unsigned(wire333[(3'h4):(1'h0)]) : reg406);
              reg539 <= {(~^($unsigned(reg532) ?
                      {$signed((7'h55)),
                          $unsigned(wire331),
                          $signed(reg453)} : $signed($unsigned(reg536)))),
                  $signed(($signed($signed(reg453)) ?
                      reg421[(5'h14):(5'h12)] : (reg393 >>> ((7'h44) >>> reg361)))),
                  $signed({(-(-reg343)), reg481})};
              reg540 = reg430[(4'hd):(2'h2)];
            end
          else
            begin
              reg538 <= {($signed((-(reg471 - reg411))) ?
                      (((reg348 ? wire419 : (7'h41)) ?
                          reg531[(5'h14):(4'hf)] : {reg371,
                              reg400,
                              reg361}) < (+(8'ha6))) : ($signed((+reg533)) > reg376[(3'h7):(3'h5)]))};
              reg540 = reg462;
              reg541 = (~(^((reg441 ? reg530 : $unsigned(wire332)) ?
                  reg406[(5'h1a):(5'h12)] : ((7'h44) ?
                      $signed(reg529) : (reg376 ? reg340 : reg348)))));
              reg542 <= ((8'hb7) ?
                  $signed($signed($unsigned((reg461 << reg520)))) : (^(reg412[(5'h10):(3'h5)] << {wire445[(4'ha):(4'h8)],
                      (reg478 >>> reg530)})));
              reg543 <= reg421;
              reg544 = reg438;
            end
          reg545 <= $signed($signed((!$unsigned((reg430 ?
              (7'h54) : (8'ha5))))));
          for (forvar546 = (1'h0); (forvar546 < (2'h3)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 = reg349[(4'hb):(1'h1)];
            end
        end
      if ((+reg547))
        begin
          if ($signed((reg537 || $signed(reg393))))
            begin
              reg548 = $unsigned(wire328[(4'hc):(2'h3)]);
              reg549 <= $unsigned($unsigned($signed({(reg341 ?
                      reg537 : wire331),
                  ((7'h48) - (7'h51)),
                  reg540})));
            end
          else
            begin
              reg549 <= {$signed($unsigned($unsigned((reg418 ?
                      reg452 : (8'h9c)))))};
              reg550 = wire446[(1'h1):(1'h1)];
              reg551 = reg531[(3'h6):(3'h5)];
              reg552 <= (reg547[(5'h17):(4'h8)] ?
                  reg340[(3'h4):(2'h3)] : wire447[(1'h1):(1'h1)]);
              reg553 <= $unsigned(((~reg538) + reg455));
              reg554 <= reg529[(4'h8):(3'h7)];
              reg555 = ((((~|(reg376 ? (8'ha3) : reg551)) ?
                      {$unsigned(reg396), $unsigned(reg524)} : (~{wire363,
                          reg465})) ?
                  (7'h40) : reg494) ^ ((~reg461) ?
                  {(~&(reg505 ? reg418 : reg530)),
                      reg400[(3'h5):(3'h4)],
                      $signed((forvar546 >= reg371))} : (reg393 ?
                      (8'hbc) : ($unsigned(wire327) & $signed(reg494)))));
            end
          if ((reg344[(5'h13):(1'h0)] ? reg453 : reg396[(4'h8):(2'h3)]))
            begin
              reg556 <= ($unsigned(reg438[(4'hc):(3'h6)]) ?
                  reg554[(4'hd):(4'hc)] : $unsigned((reg406[(5'h15):(3'h6)] >>> $signed((~reg477)))));
              reg557 <= wire363;
              reg558 = $signed((^$signed((reg430[(5'h11):(4'hb)] ?
                  $signed(wire329) : reg455))));
            end
          else
            begin
              reg556 <= $unsigned($unsigned((7'h4b)));
              reg558 = $signed(reg552[(2'h3):(2'h3)]);
              reg559 = reg361;
              reg560 <= {(7'h48), (-$unsigned($signed((reg434 == reg458))))};
              reg561 = {(!$signed((reg549 <= (reg351 ? reg411 : (7'h41))))),
                  (~|reg503[(4'h8):(3'h4)]),
                  reg448};
              reg562 = wire420[(5'h17):(3'h4)];
              reg563 <= (($signed($unsigned(reg553)) ?
                      $signed((!reg548)) : $signed((~^{(7'h4c), (7'h43)}))) ?
                  $signed($signed((7'h57))) : $signed(((wire335 ?
                          (reg452 ? reg478 : reg537) : $signed(reg396)) ?
                      {$unsigned(reg531),
                          {reg471, reg461, (8'hbe)}} : $unsigned((^~reg561)))));
            end
          reg564 <= (((^~(&(-reg403))) ~^ $signed((-$signed(wire332)))) ?
              (^~$signed((&$unsigned(reg540)))) : $unsigned(wire447[(1'h1):(1'h0)]));
        end
      else
        begin
          reg549 <= $signed(((reg393 ~^ $signed((~|reg529))) ~^ (((reg369 ?
                  reg341 : (8'hba)) > (reg542 & reg532)) ?
              reg393 : ((+reg369) < (reg524 ? (8'haa) : reg344)))));
          if ($unsigned((reg544[(3'h5):(3'h5)] >> reg383)))
            begin
              reg552 <= $signed((($unsigned(reg458[(2'h2):(2'h2)]) ^ (!$unsigned(reg562))) ?
                  reg343[(5'h12):(4'hb)] : (($unsigned(reg436) ?
                      $unsigned(reg393) : wire328[(4'hc):(1'h0)]) ^ reg351)));
              reg553 <= ($unsigned(reg544) ?
                  $signed($signed((((7'h52) ? (8'hbb) : reg386) ?
                      $unsigned((7'h4b)) : reg561[(5'h19):(2'h3)]))) : $unsigned(reg390[(2'h2):(1'h0)]));
              reg554 <= ((($signed(reg413[(2'h2):(1'h0)]) ~^ ($unsigned(reg554) ?
                      {reg501, reg545, (7'h44)} : (wire446 >> wire327))) ?
                  wire332 : {(~^{(8'ha2)}),
                      (((8'ha7) ? reg411 : reg557) ?
                          $signed(reg368) : $unsigned(reg477)),
                      $signed(((8'ha8) ?
                          reg448 : (8'hb4)))}) <<< reg386[(1'h0):(1'h0)]);
              reg555 = (7'h54);
              reg558 = (7'h42);
            end
          else
            begin
              reg552 <= reg563;
              reg553 <= reg503;
              reg555 = $unsigned((reg474[(2'h2):(1'h0)] ?
                  {($signed(reg482) < (reg390 ? reg412 : wire332)),
                      {$unsigned(reg540), (!reg436), wire329}} : reg417));
              reg556 <= $signed($signed($unsigned(reg518[(1'h1):(1'h1)])));
              reg558 = (!reg507);
            end
        end
      if ((|$signed({wire331[(4'ha):(3'h5)],
          (reg438[(3'h5):(3'h4)] <= wire420),
          (wire447 ? (reg458 ? (8'haf) : reg551) : (reg458 ^~ (8'ha4)))})))
        begin
          if ((^$signed(reg343)))
            begin
              reg565 = (|($signed($unsigned((wire447 >= reg559))) ?
                  (^wire334) : reg441[(5'h1b):(5'h15)]));
              reg566 = $unsigned(reg558);
              reg567 = $unsigned({reg551[(5'h10):(5'h10)]});
              reg568 <= wire420;
            end
          else
            begin
              reg565 = reg494[(2'h3):(2'h3)];
              reg566 = reg532;
              reg567 = (-($unsigned($signed($signed(reg540))) ?
                  {reg538,
                      reg453,
                      {$signed(reg406),
                          $signed(reg494)}} : (reg452[(3'h5):(3'h4)] ?
                      reg556[(1'h1):(1'h1)] : $unsigned($signed(reg390)))));
              reg569 = $unsigned(reg351);
              reg570 = (&($unsigned($unsigned(wire447[(1'h1):(1'h0)])) ?
                  (reg494[(3'h6):(2'h3)] ?
                      reg396 : reg531[(5'h12):(4'hb)]) : ($signed(reg435[(1'h0):(1'h0)]) >>> (-reg531))));
            end
        end
      else
        begin
          for (forvar565 = (1'h0); (forvar565 < (3'h5)); forvar565 = (forvar565 + (1'h1)))
            begin
              reg568 <= (^~$signed($unsigned(reg527)));
              reg571 <= reg529[(1'h0):(1'h0)];
            end
          reg572 <= $signed((($unsigned($signed(reg568)) < ($signed(reg564) ?
              reg458[(4'h8):(2'h3)] : (reg544 < (7'h4e)))) - (|reg527[(5'h11):(1'h1)])));
          reg573 <= $signed(reg477[(5'h10):(3'h4)]);
          reg574 <= reg418[(1'h0):(1'h0)];
          reg575 <= (((~|($unsigned(wire334) ?
                      ((7'h49) ? reg399 : reg411) : $signed(reg528))) ?
                  ((((7'h4b) >> wire330) ?
                      (reg571 - reg377) : $unsigned(reg531)) ^~ reg507) : reg537[(3'h6):(2'h3)]) ?
              $signed({(reg430 <= reg471),
                  $signed((^~wire447)),
                  (|(~|reg388))}) : (!{reg370,
                  $unsigned((~reg557)),
                  reg421[(5'h11):(3'h7)]}));
        end
      reg576 = $unsigned({$signed(wire363)});
    end
  assign wire577 = (7'h4e);
  always
    @(posedge clk) begin
      for (forvar578 = (1'h0); (forvar578 < (2'h2)); forvar578 = (forvar578 + (1'h1)))
        begin
          for (forvar579 = (1'h0); (forvar579 < (3'h6)); forvar579 = (forvar579 + (1'h1)))
            begin
              reg580 = $unsigned(reg455[(3'h4):(1'h0)]);
              reg581 = (|(+$unsigned(($unsigned((8'ha1)) ?
                  ((8'hba) != (8'hb8)) : reg478[(4'h9):(2'h3)]))));
              reg582 <= $unsigned(reg530[(3'h7):(2'h2)]);
              reg583 <= (reg452 >>> (reg538[(2'h2):(1'h1)] != (~wire334)));
            end
          for (forvar584 = (1'h0); (forvar584 < (1'h1)); forvar584 = (forvar584 + (1'h1)))
            begin
              reg585 = reg545;
              reg586 <= (-(!$unsigned((((8'ha3) ?
                  reg574 : reg545) >= (^~(7'h43))))));
              reg587 <= $unsigned(wire331[(4'hd):(2'h3)]);
              reg588 = (|reg452);
              reg589 = ($unsigned((!$unsigned(reg537[(3'h4):(2'h2)]))) == reg585);
            end
          if ((~^{$unsigned(((8'ha3) >>> (reg536 ? (8'ha6) : reg575)))}))
            begin
              reg590 <= ((~($signed(((8'hbb) & reg351)) ?
                      reg563[(1'h0):(1'h0)] : (((8'hb6) & reg453) > $unsigned(reg572)))) ?
                  ((~|((reg418 ?
                      reg582 : (8'ha6)) + reg359)) < (~|reg505)) : $unsigned(forvar584));
            end
          else
            begin
              reg591 = (^$unsigned((reg563[(2'h2):(1'h0)] ?
                  (|(wire577 ? (8'hb7) : reg538)) : reg481[(4'hf):(1'h1)])));
              reg592 = ($unsigned(wire332[(2'h3):(2'h2)]) ?
                  (~^(((7'h47) < $unsigned(reg389)) ?
                      (+reg536) : $signed((reg539 <= (8'ha2))))) : (($unsigned((~(8'hb0))) <<< (~&$unsigned(reg474))) >= reg574));
              reg593 = (!$unsigned(($signed((reg560 ? reg376 : reg590)) ?
                  reg481[(5'h14):(5'h13)] : reg536[(3'h7):(2'h3)])));
              reg594 = ({reg582} <<< ((~$signed(reg437)) >>> reg412));
            end
        end
      if ((reg348 ?
          ((wire329[(5'h1c):(1'h0)] - ((reg368 || reg351) ?
                  reg351[(5'h13):(5'h10)] : (+reg481))) ?
              wire446[(1'h0):(1'h0)] : $unsigned((((8'ha8) >> (8'hb2)) ?
                  $unsigned(wire328) : (reg542 ? reg370 : reg471)))) : reg386))
        begin
          reg595 <= $unsigned({reg403,
              {({(8'hbe), reg448, reg375} ?
                      $signed(reg518) : $unsigned(reg554)),
                  $signed(reg436[(3'h6):(2'h3)])},
              $unsigned({$signed((7'h4b)), $unsigned(reg538)})});
          reg596 = (7'h45);
        end
      else
        begin
          if ((&wire333))
            begin
              reg596 = $signed($unsigned(reg503));
            end
          else
            begin
              reg596 = reg507[(2'h2):(1'h1)];
              reg597 = (~&(~&(~&$unsigned(reg371))));
              reg598 <= (~&{reg534[(5'h12):(4'hb)],
                  (reg477 ?
                      $unsigned($unsigned(reg341)) : $signed($signed(reg563))),
                  $unsigned(reg543[(4'h8):(3'h5)])});
              reg599 = $unsigned((^(7'h51)));
            end
          if ({(8'h9f)})
            begin
              reg600 = $unsigned(({wire577} ? (8'hb6) : reg492));
              reg601 <= {$signed({((+reg452) > reg581[(2'h3):(1'h0)]),
                      (((8'hbe) >> reg421) >>> {(8'ha8), reg542})})};
              reg602 <= {$unsigned(({{reg412, reg600}, ((7'h47) + wire419)} ?
                      reg448 : $unsigned(reg582[(3'h5):(2'h3)])))};
              reg603 <= wire327[(3'h6):(1'h0)];
              reg604 = reg482;
              reg605 = ((8'hb4) ?
                  ($unsigned(($unsigned(wire327) == (~&(8'hb6)))) || reg531) : {$signed((reg588 << (reg542 & (8'ha5)))),
                      reg598,
                      reg520});
              reg606 = reg583;
            end
          else
            begin
              reg600 = (~|({wire446,
                      (reg452[(4'h9):(3'h6)] >>> (reg425 ^ forvar578)),
                      reg417[(1'h0):(1'h0)]} ?
                  (($signed(reg601) ?
                          reg520[(1'h1):(1'h1)] : wire332[(1'h1):(1'h1)]) ?
                      (reg370 ?
                          reg520 : reg505) : reg587[(1'h1):(1'h0)]) : $unsigned({reg598[(5'h13):(3'h7)],
                      reg400[(1'h1):(1'h1)]})));
              reg604 = (~&$signed($signed(wire445[(5'h13):(1'h1)])));
              reg607 <= reg377;
            end
          if ((reg430[(2'h3):(1'h1)] ?
              ($signed(forvar578[(4'h9):(1'h1)]) ?
                  $signed($unsigned($unsigned(reg505))) : {$signed(reg605),
                      ((|reg595) ?
                          (|(7'h40)) : reg518)}) : ($signed(reg518[(1'h1):(1'h0)]) ?
                  $signed(($unsigned(reg553) ~^ (-(8'hba)))) : ($signed($signed((8'hae))) ?
                      (|reg590) : $unsigned((reg568 ^~ reg412))))))
            begin
              reg608 <= ({{reg564[(3'h7):(3'h7)],
                      (!(reg437 | reg390)),
                      $unsigned(reg343)},
                  (((reg388 ? reg563 : reg386) ?
                      (reg524 ? reg369 : wire328) : (reg461 ?
                          (7'h51) : reg341)) <<< reg474),
                  {wire334,
                      $signed(reg545),
                      ($unsigned(reg477) ?
                          reg600 : (reg386 | reg503))}} + (~&$unsigned(((reg591 >> reg572) ?
                  (!(7'h41)) : ((8'hb8) >= reg545)))));
              reg609 <= $unsigned(({(!(+(8'h9d))),
                      (+(reg600 ? reg477 : reg572))} ?
                  (+$signed((&reg602))) : (reg602 >= $unsigned((~|wire445)))));
              reg610 <= reg600;
              reg611 <= $signed(({(^(8'hb8)), reg406} ?
                  (reg383 >= reg518[(4'h9):(2'h3)]) : reg590[(5'h1a):(4'hd)]));
              reg612 = $unsigned($unsigned({(&reg494[(2'h2):(2'h2)]),
                  wire327}));
              reg613 <= reg393[(4'hd):(4'hc)];
              reg614 <= (^~(reg534 ? wire577 : reg441));
            end
          else
            begin
              reg608 <= ((!(((wire363 ? (8'ha8) : reg368) ?
                      $unsigned(reg383) : (wire446 ? reg393 : (8'ha3))) ?
                  ((!reg593) ? (+reg588) : (reg413 | reg592)) : ((wire327 ?
                          reg538 : reg572) ?
                      (~|(7'h4e)) : (&reg588)))) ^ (8'h9e));
              reg612 = $signed(({((reg375 <= reg390) & $signed(wire447)),
                      $unsigned($signed(reg536)),
                      reg543[(5'h11):(3'h7)]} ?
                  forvar579[(3'h5):(3'h5)] : reg549));
              reg615 = reg377[(4'h9):(1'h0)];
            end
          if ((8'hb6))
            begin
              reg616 <= wire328;
            end
          else
            begin
              reg617 = $signed($unsigned((-$unsigned($signed(reg434)))));
              reg618 <= $signed(wire525);
              reg619 <= (|((~|reg371[(5'h11):(5'h11)]) >= reg534[(3'h6):(2'h3)]));
              reg620 = {$unsigned(({(!reg568), $unsigned(reg538)} ?
                      reg601[(1'h1):(1'h1)] : (^~reg591[(4'ha):(4'h8)]))),
                  reg375[(3'h4):(3'h4)],
                  $unsigned($signed(reg507[(4'hd):(3'h6)]))};
            end
        end
      for (forvar621 = (1'h0); (forvar621 < (1'h0)); forvar621 = (forvar621 + (1'h1)))
        begin
          reg622 <= (8'h9c);
          for (forvar623 = (1'h0); (forvar623 < (2'h2)); forvar623 = (forvar623 + (1'h1)))
            begin
              reg624 <= $unsigned(reg501[(2'h2):(2'h2)]);
              reg625 = $unsigned((reg518[(1'h0):(1'h0)] ?
                  ($unsigned(reg624) ^ $signed((reg519 ?
                      reg571 : reg441))) : reg607));
            end
          if ((reg543 > {$unsigned(((wire332 ? reg349 : reg474) >>> {reg572,
                  reg619})),
              $unsigned($signed((wire328 - reg613)))}))
            begin
              reg626 <= $signed(reg519[(2'h2):(2'h2)]);
              reg627 <= $unsigned($signed((^~$unsigned((^~reg351)))));
              reg628 = $unsigned(({reg615[(5'h12):(3'h4)]} ?
                  (&$unsigned((forvar584 < reg481))) : $unsigned({reg396,
                      reg611[(4'h9):(2'h2)]})));
              reg629 <= reg441[(4'h9):(3'h4)];
              reg630 = {reg413};
              reg631 <= (~^forvar578[(4'h8):(2'h3)]);
            end
          else
            begin
              reg628 = (~reg518);
              reg629 <= (reg629[(1'h0):(1'h0)] ?
                  (^~$unsigned(reg585[(5'h14):(1'h1)])) : $unsigned($unsigned({(~|reg612),
                      forvar621,
                      wire328})));
              reg631 <= ((((reg560[(3'h4):(1'h0)] ~^ reg344[(5'h13):(3'h4)]) != reg629) <<< (8'hba)) ?
                  {$unsigned($signed((+reg393))), wire329} : {(reg478 ?
                          wire332 : (wire330 ? (^reg471) : reg534)),
                      reg530});
            end
          if ($unsigned(reg430[(4'hb):(2'h3)]))
            begin
              reg632 = $unsigned(reg537[(3'h7):(2'h2)]);
              reg633 <= $unsigned((^~reg582[(2'h2):(2'h2)]));
              reg634 <= reg571;
              reg635 <= reg523;
              reg636 <= $unsigned($unsigned((reg343 & (~^(-reg552)))));
              reg637 <= {reg602[(4'ha):(3'h6)], reg354[(3'h4):(3'h4)]};
              reg638 = reg386[(2'h2):(1'h0)];
            end
          else
            begin
              reg633 <= $signed((~&$signed(reg361[(4'hc):(3'h6)])));
              reg638 = (+(reg351[(5'h12):(4'hc)] ?
                  (reg478 >= ((8'haf) ?
                      $unsigned(reg626) : (~(8'hb2)))) : $unsigned($signed((reg581 * reg616)))));
            end
          reg639 <= $signed(($unsigned($unsigned({reg361, reg585})) ?
              (reg636 ?
                  ((|wire419) ?
                      reg593 : $signed((8'hbf))) : (~|(reg481 <<< reg592))) : (((reg361 ?
                      (8'hb5) : reg597) ?
                  (+reg627) : $unsigned(reg583)) | reg616[(1'h1):(1'h0)])));
        end
      for (forvar640 = (1'h0); (forvar640 < (1'h1)); forvar640 = (forvar640 + (1'h1)))
        begin
          reg641 = ((^(&$unsigned(((8'haa) ? forvar621 : reg602)))) ?
              {(~&((|reg605) ? reg344[(2'h2):(1'h1)] : reg609)),
                  reg608} : reg368);
          for (forvar642 = (1'h0); (forvar642 < (3'h6)); forvar642 = (forvar642 + (1'h1)))
            begin
              reg643 <= reg358[(5'h17):(5'h12)];
              reg644 <= (reg582[(4'h9):(4'h9)] << {(((reg545 ?
                          (7'h4d) : (8'ha1)) ?
                      $unsigned(reg611) : reg631[(4'hf):(2'h2)]) <<< (^(reg390 ?
                      reg620 : reg629))),
                  reg597[(3'h4):(2'h3)],
                  $signed(reg354)});
              reg645 = (((((reg595 ?
                      reg531 : reg574) > reg418) << reg624) ^ $unsigned(reg403[(3'h6):(3'h5)])) ?
                  reg574[(5'h12):(4'h8)] : $unsigned($unsigned((|wire445[(4'hb):(4'hb)]))));
              reg646 = reg605;
              reg647 = forvar621;
              reg648 = reg430[(4'hc):(3'h7)];
            end
          for (forvar649 = (1'h0); (forvar649 < (1'h0)); forvar649 = (forvar649 + (1'h1)))
            begin
              reg650 = (&{forvar621[(4'h9):(2'h3)],
                  (($signed(wire332) ? {(8'ha6)} : (~|(8'hb2))) ?
                      reg474[(1'h0):(1'h0)] : $unsigned(reg389[(1'h0):(1'h0)]))});
              reg651 = (&reg596);
              reg652 <= $signed($unsigned($unsigned($unsigned((forvar579 - reg389)))));
              reg653 <= $signed($signed((7'h44)));
              reg654 <= $unsigned((reg492 ?
                  $signed((^$signed(wire577))) : (!reg647)));
              reg655 = ($signed($unsigned(($unsigned((8'hbf)) < $signed(reg452)))) ?
                  (reg608 == reg341) : reg437);
              reg656 <= $signed(((~$unsigned($signed(reg631))) ?
                  (((reg344 << reg494) == $signed(reg610)) ?
                      ($unsigned(reg399) ?
                          (reg603 ?
                              reg461 : wire525) : (~^reg648)) : $signed($signed(reg376))) : reg412[(4'h9):(1'h0)]));
            end
          if (($signed($unsigned($unsigned($signed((8'ha9))))) >>> $unsigned(((~|reg393[(1'h1):(1'h0)]) ^ $unsigned((reg634 == reg406))))))
            begin
              reg657 = {{$signed(reg631), reg564, reg652},
                  ((reg539 ? reg537 : $unsigned((reg610 >> reg452))) ?
                      (7'h55) : ($signed({forvar621, reg543, (7'h4f)}) ?
                          reg361 : $signed($signed((8'ha3))))),
                  ($unsigned(reg607[(3'h7):(3'h6)]) * {{$signed(wire469),
                          (~reg644)}})};
              reg658 <= $signed($signed((^(|(|reg572)))));
              reg659 = reg477[(1'h0):(1'h0)];
              reg660 = $signed(reg351);
              reg661 = reg643[(4'h8):(1'h1)];
              reg662 <= (reg452 << reg505[(2'h2):(2'h2)]);
              reg663 = ((|((reg614 ? {reg657, reg654, reg651} : (~&reg534)) ?
                  $unsigned((reg589 ?
                      (7'h40) : reg564)) : reg581)) >= (((reg629[(1'h1):(1'h1)] && (reg660 >>> reg492)) || $signed($signed((7'h50)))) ?
                  ($unsigned((wire363 <= wire469)) ?
                      $signed((~^wire525)) : $unsigned((~wire447))) : ((~|reg608) & $unsigned(forvar640[(4'hb):(1'h0)]))));
            end
          else
            begin
              reg658 <= {$signed($signed($unsigned((reg607 <<< reg341)))),
                  reg389,
                  (wire420 ? ($signed($signed(wire419)) >> (8'ha7)) : reg523)};
              reg662 <= reg455;
              reg663 = reg616;
              reg664 = (~&$unsigned(reg436));
              reg665 <= wire331[(4'hb):(4'h9)];
              reg666 = reg665[(3'h6):(3'h6)];
            end
          reg667 <= wire446[(2'h2):(1'h0)];
          reg668 <= ((reg341[(1'h0):(1'h0)] * (($signed(reg646) >> reg639[(4'hc):(3'h7)]) ~^ $signed($unsigned(reg549)))) <= ($signed(((~|reg411) ?
                  reg524 : reg371[(4'ha):(4'ha)])) ?
              reg556[(4'h8):(4'h8)] : {(~(reg658 < (8'h9c))),
                  reg343[(4'hb):(4'h9)]}));
        end
      for (forvar669 = (1'h0); (forvar669 < (1'h1)); forvar669 = (forvar669 + (1'h1)))
        begin
          for (forvar670 = (1'h0); (forvar670 < (1'h1)); forvar670 = (forvar670 + (1'h1)))
            begin
              reg671 = ((~&(~&reg591[(3'h5):(3'h4)])) ?
                  {$unsigned($unsigned({reg478, reg406, reg633})),
                      $signed($unsigned((reg637 ? reg604 : reg421))),
                      (((~^reg400) | $signed(reg645)) >= ($signed((7'h50)) ?
                          wire577 : $signed(wire525)))} : {reg358});
              reg672 <= wire419;
              reg673 = reg661;
              reg674 = (8'hac);
              reg675 = (reg629[(1'h0):(1'h0)] ?
                  $unsigned((((7'h47) || {reg627, reg644}) ?
                      reg610 : reg574)) : (^{reg655,
                      $unsigned($signed(reg370))}));
              reg676 <= reg528;
            end
          reg677 = (reg598 ?
              $signed($signed($unsigned($unsigned(reg668)))) : reg481[(2'h3):(2'h3)]);
          reg678 <= $unsigned($signed(reg675));
        end
      reg679 <= reg358[(5'h12):(2'h2)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2467
#(parameter param2802 = (((&((+(8'hb8)) ? (~^(7'h46)) : ((8'hb9) <= (7'h53)))) ? (((-(8'ha3)) ? (-(8'hae)) : (-(8'hb6))) ? (|((8'h9f) * (8'h9c))) : {(7'h47)}) : ((((8'hb2) >= (7'h40)) || ((8'ha2) <= (7'h4c))) ? {((8'hb7) ? (7'h56) : (7'h54)), ((7'h44) << (7'h4d)), ((8'hac) ? (8'hb3) : (8'h9d))} : ((~&(8'hbb)) != ((8'haa) - (7'h46))))) != ((^~((7'h47) << ((7'h49) ? (7'h41) : (7'h41)))) && (((~|(8'hbb)) ? ((7'h52) <= (8'h9c)) : (^~(7'h48))) ? (|((8'haa) | (8'ha8))) : ((^~(8'hb0)) ? ((8'hba) ? (7'h4d) : (7'h52)) : {(8'hae)})))), 
parameter param2803 = param2802)
(y, clk, wire2472, wire2471, wire2470, wire2469, wire2468);
  output wire [(32'h1667):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire2472;
  input wire signed [(3'h7):(1'h0)] wire2471;
  input wire [(5'h12):(1'h0)] wire2470;
  input wire [(4'hb):(1'h0)] wire2469;
  input wire [(5'h13):(1'h0)] wire2468;
  wire [(5'h11):(1'h0)] wire2696;
  wire [(5'h1e):(1'h0)] wire2695;
  wire [(5'h15):(1'h0)] wire2694;
  wire [(5'h1f):(1'h0)] wire2664;
  wire [(4'hf):(1'h0)] wire2663;
  wire signed [(4'hb):(1'h0)] wire2662;
  wire [(5'h1c):(1'h0)] wire2640;
  wire [(5'h1f):(1'h0)] wire2475;
  wire signed [(5'h11):(1'h0)] wire2474;
  wire signed [(4'ha):(1'h0)] wire2473;
  reg signed [(2'h3):(1'h0)] reg2801 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2799 = (1'h0);
  reg [(5'h11):(1'h0)] reg2797 = (1'h0);
  reg [(5'h11):(1'h0)] reg2796 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2795 = (1'h0);
  reg [(3'h4):(1'h0)] reg2792 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2790 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2789 = (1'h0);
  reg [(3'h6):(1'h0)] reg2787 = (1'h0);
  reg [(3'h7):(1'h0)] reg2786 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2783 = (1'h0);
  reg [(3'h5):(1'h0)] reg2781 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2779 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2778 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2776 = (1'h0);
  reg [(5'h11):(1'h0)] reg2775 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2772 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2770 = (1'h0);
  reg [(5'h12):(1'h0)] reg2768 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2765 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2764 = (1'h0);
  reg [(5'h15):(1'h0)] reg2763 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2762 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2761 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2757 = (1'h0);
  reg [(5'h16):(1'h0)] reg2751 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2750 = (1'h0);
  reg [(4'hd):(1'h0)] reg2748 = (1'h0);
  reg [(3'h7):(1'h0)] reg2747 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2746 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2744 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2743 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2742 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2738 = (1'h0);
  reg [(4'hc):(1'h0)] reg2737 = (1'h0);
  reg [(5'h12):(1'h0)] reg2735 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2733 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2731 = (1'h0);
  reg [(5'h14):(1'h0)] reg2730 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2729 = (1'h0);
  reg [(4'hb):(1'h0)] reg2727 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2726 = (1'h0);
  reg [(4'hd):(1'h0)] reg2724 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2723 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2722 = (1'h0);
  reg [(5'h19):(1'h0)] reg2721 = (1'h0);
  reg [(3'h6):(1'h0)] reg2718 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2717 = (1'h0);
  reg [(5'h18):(1'h0)] reg2716 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2714 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2710 = (1'h0);
  reg [(5'h11):(1'h0)] reg2709 = (1'h0);
  reg [(4'h8):(1'h0)] reg2707 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2706 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2704 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2702 = (1'h0);
  reg [(4'hd):(1'h0)] reg2701 = (1'h0);
  reg [(4'hc):(1'h0)] reg2700 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2693 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2690 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2688 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2685 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2684 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2679 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2676 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2675 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2674 = (1'h0);
  reg [(5'h19):(1'h0)] reg2671 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2670 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2668 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2660 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2659 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2656 = (1'h0);
  reg [(4'hd):(1'h0)] reg2655 = (1'h0);
  reg [(5'h16):(1'h0)] reg2654 = (1'h0);
  reg [(3'h5):(1'h0)] reg2651 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2649 = (1'h0);
  reg [(4'hb):(1'h0)] reg2646 = (1'h0);
  reg [(3'h6):(1'h0)] reg2641 = (1'h0);
  reg [(5'h15):(1'h0)] reg2638 = (1'h0);
  reg [(3'h4):(1'h0)] reg2635 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2634 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2630 = (1'h0);
  reg [(2'h3):(1'h0)] reg2627 = (1'h0);
  reg [(5'h14):(1'h0)] reg2625 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2617 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2615 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2614 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2613 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2611 = (1'h0);
  reg [(4'hf):(1'h0)] reg2608 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2605 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2604 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2602 = (1'h0);
  reg [(3'h6):(1'h0)] reg2599 = (1'h0);
  reg [(5'h19):(1'h0)] reg2597 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2596 = (1'h0);
  reg [(5'h16):(1'h0)] reg2594 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2593 = (1'h0);
  reg [(5'h15):(1'h0)] reg2591 = (1'h0);
  reg [(4'hd):(1'h0)] reg2590 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2589 = (1'h0);
  reg [(3'h6):(1'h0)] reg2588 = (1'h0);
  reg [(5'h14):(1'h0)] reg2586 = (1'h0);
  reg [(5'h14):(1'h0)] reg2583 = (1'h0);
  reg [(2'h3):(1'h0)] reg2582 = (1'h0);
  reg [(4'hc):(1'h0)] reg2580 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2579 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2578 = (1'h0);
  reg [(2'h3):(1'h0)] reg2577 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2556 = (1'h0);
  reg [(5'h14):(1'h0)] reg2574 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2573 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2571 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2569 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2567 = (1'h0);
  reg [(4'hc):(1'h0)] reg2565 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2564 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2562 = (1'h0);
  reg [(4'he):(1'h0)] reg2561 = (1'h0);
  reg [(2'h3):(1'h0)] reg2559 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2558 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2557 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2555 = (1'h0);
  reg [(4'ha):(1'h0)] reg2553 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2551 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2547 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2545 = (1'h0);
  reg [(4'h8):(1'h0)] reg2544 = (1'h0);
  reg [(4'h9):(1'h0)] reg2543 = (1'h0);
  reg [(5'h16):(1'h0)] reg2542 = (1'h0);
  reg [(5'h14):(1'h0)] reg2541 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2539 = (1'h0);
  reg [(4'hf):(1'h0)] reg2538 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2537 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2536 = (1'h0);
  reg [(2'h2):(1'h0)] reg2531 = (1'h0);
  reg [(5'h10):(1'h0)] reg2528 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2526 = (1'h0);
  reg [(4'he):(1'h0)] reg2525 = (1'h0);
  reg [(3'h4):(1'h0)] reg2523 = (1'h0);
  reg [(4'hc):(1'h0)] reg2521 = (1'h0);
  reg [(5'h19):(1'h0)] reg2520 = (1'h0);
  reg [(4'ha):(1'h0)] reg2517 = (1'h0);
  reg [(5'h15):(1'h0)] reg2515 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2510 = (1'h0);
  reg [(5'h17):(1'h0)] reg2504 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2513 = (1'h0);
  reg [(4'h8):(1'h0)] reg2507 = (1'h0);
  reg [(3'h4):(1'h0)] reg2501 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2497 = (1'h0);
  reg [(3'h5):(1'h0)] reg2495 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2493 = (1'h0);
  reg [(3'h4):(1'h0)] reg2488 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2487 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2486 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2484 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2480 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2478 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2800 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2798 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar2794 = (1'h0);
  reg [(4'hf):(1'h0)] reg2793 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2791 = (1'h0);
  reg [(5'h19):(1'h0)] reg2784 = (1'h0);
  reg [(5'h16):(1'h0)] forvar2782 = (1'h0);
  reg [(3'h6):(1'h0)] reg2788 = (1'h0);
  reg [(5'h16):(1'h0)] reg2785 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2784 = (1'h0);
  reg [(4'hc):(1'h0)] reg2782 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2780 = (1'h0);
  reg [(5'h14):(1'h0)] reg2777 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2774 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2773 = (1'h0);
  reg [(5'h16):(1'h0)] reg2771 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2769 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2767 = (1'h0);
  reg [(5'h12):(1'h0)] reg2766 = (1'h0);
  reg [(3'h4):(1'h0)] reg2760 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2759 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2758 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2756 = (1'h0);
  reg [(5'h14):(1'h0)] reg2755 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2754 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2753 = (1'h0);
  reg [(4'hc):(1'h0)] reg2752 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2748 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2749 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2745 = (1'h0);
  reg [(5'h15):(1'h0)] reg2741 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2740 = (1'h0);
  reg [(5'h14):(1'h0)] reg2739 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2737 = (1'h0);
  reg [(4'h8):(1'h0)] reg2725 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2736 = (1'h0);
  reg [(5'h18):(1'h0)] reg2734 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2732 = (1'h0);
  reg [(4'h9):(1'h0)] reg2728 = (1'h0);
  reg [(5'h12):(1'h0)] forvar2725 = (1'h0);
  reg [(3'h6):(1'h0)] reg2720 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2719 = (1'h0);
  reg [(2'h2):(1'h0)] reg2715 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2713 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2712 = (1'h0);
  reg [(3'h6):(1'h0)] reg2711 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2708 = (1'h0);
  reg [(5'h17):(1'h0)] reg2705 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2703 = (1'h0);
  reg [(4'hf):(1'h0)] reg2699 = (1'h0);
  reg [(3'h7):(1'h0)] reg2698 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2697 = (1'h0);
  reg [(5'h15):(1'h0)] reg2692 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2691 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2689 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2687 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2686 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2683 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2682 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2681 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2680 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2677 = (1'h0);
  reg [(5'h12):(1'h0)] reg2673 = (1'h0);
  reg [(5'h13):(1'h0)] reg2672 = (1'h0);
  reg [(5'h14):(1'h0)] reg2669 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2667 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2666 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2665 = (1'h0);
  reg [(5'h12):(1'h0)] reg2661 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2658 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2657 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2653 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2652 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar2650 = (1'h0);
  reg [(3'h5):(1'h0)] reg2648 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2647 = (1'h0);
  reg [(5'h12):(1'h0)] reg2645 = (1'h0);
  reg [(5'h12):(1'h0)] reg2644 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2643 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2642 = (1'h0);
  reg [(4'h9):(1'h0)] reg2639 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2637 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2636 = (1'h0);
  reg [(5'h15):(1'h0)] reg2633 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2632 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2631 = (1'h0);
  reg [(5'h18):(1'h0)] reg2629 = (1'h0);
  reg [(4'ha):(1'h0)] reg2628 = (1'h0);
  reg [(5'h12):(1'h0)] reg2626 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2624 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2623 = (1'h0);
  reg [(5'h11):(1'h0)] reg2622 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2621 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2620 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2619 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2618 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2616 = (1'h0);
  reg [(2'h2):(1'h0)] reg2612 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar2610 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2609 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2607 = (1'h0);
  reg [(5'h18):(1'h0)] reg2606 = (1'h0);
  reg [(5'h15):(1'h0)] reg2603 = (1'h0);
  reg [(2'h3):(1'h0)] reg2601 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2600 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2598 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2595 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2592 = (1'h0);
  reg [(3'h4):(1'h0)] reg2587 = (1'h0);
  reg [(4'hc):(1'h0)] reg2585 = (1'h0);
  reg [(4'h9):(1'h0)] reg2584 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2581 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2576 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2575 = (1'h0);
  reg [(3'h7):(1'h0)] reg2572 = (1'h0);
  reg [(4'hb):(1'h0)] reg2570 = (1'h0);
  reg [(5'h10):(1'h0)] reg2568 = (1'h0);
  reg [(4'ha):(1'h0)] reg2566 = (1'h0);
  reg [(2'h3):(1'h0)] reg2563 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2560 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2556 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2554 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2552 = (1'h0);
  reg [(4'he):(1'h0)] reg2550 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2549 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2548 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2546 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2540 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2535 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2534 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2533 = (1'h0);
  reg [(2'h3):(1'h0)] reg2532 = (1'h0);
  reg [(3'h4):(1'h0)] reg2530 = (1'h0);
  reg [(5'h19):(1'h0)] reg2529 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2527 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2524 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2522 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2519 = (1'h0);
  reg [(5'h18):(1'h0)] reg2518 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2516 = (1'h0);
  reg [(5'h14):(1'h0)] reg2514 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2512 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2511 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2510 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2509 = (1'h0);
  reg [(3'h4):(1'h0)] reg2508 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2506 = (1'h0);
  reg [(5'h13):(1'h0)] reg2505 = (1'h0);
  reg [(5'h16):(1'h0)] forvar2504 = (1'h0);
  reg [(4'h8):(1'h0)] reg2503 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2502 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2500 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar2499 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2498 = (1'h0);
  reg [(5'h15):(1'h0)] reg2496 = (1'h0);
  reg [(5'h12):(1'h0)] reg2494 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2492 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2491 = (1'h0);
  reg [(4'h8):(1'h0)] reg2490 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2489 = (1'h0);
  reg [(3'h7):(1'h0)] reg2485 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2483 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2482 = (1'h0);
  reg [(3'h7):(1'h0)] reg2481 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2479 = (1'h0);
  reg [(4'hd):(1'h0)] reg2477 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2476 = (1'h0);
  assign y = {wire2696,
                 wire2695,
                 wire2694,
                 wire2664,
                 wire2663,
                 wire2662,
                 wire2640,
                 wire2475,
                 wire2474,
                 wire2473,
                 reg2801,
                 reg2799,
                 reg2797,
                 reg2796,
                 reg2795,
                 reg2792,
                 reg2790,
                 reg2789,
                 reg2787,
                 reg2786,
                 reg2783,
                 reg2781,
                 reg2779,
                 reg2778,
                 reg2776,
                 reg2775,
                 reg2772,
                 reg2770,
                 reg2768,
                 reg2765,
                 reg2764,
                 reg2763,
                 reg2762,
                 reg2761,
                 reg2757,
                 reg2751,
                 reg2750,
                 reg2748,
                 reg2747,
                 reg2746,
                 reg2744,
                 reg2743,
                 reg2742,
                 reg2738,
                 reg2737,
                 reg2735,
                 reg2733,
                 reg2731,
                 reg2730,
                 reg2729,
                 reg2727,
                 reg2726,
                 reg2724,
                 reg2723,
                 reg2722,
                 reg2721,
                 reg2718,
                 reg2717,
                 reg2716,
                 reg2714,
                 reg2710,
                 reg2709,
                 reg2707,
                 reg2706,
                 reg2704,
                 reg2702,
                 reg2701,
                 reg2700,
                 reg2693,
                 reg2690,
                 reg2688,
                 reg2685,
                 reg2684,
                 reg2679,
                 reg2678,
                 reg2676,
                 reg2675,
                 reg2674,
                 reg2671,
                 reg2670,
                 reg2668,
                 reg2660,
                 reg2659,
                 reg2656,
                 reg2655,
                 reg2654,
                 reg2651,
                 reg2649,
                 reg2646,
                 reg2641,
                 reg2638,
                 reg2635,
                 reg2634,
                 reg2630,
                 reg2627,
                 reg2625,
                 reg2617,
                 reg2615,
                 reg2614,
                 reg2613,
                 reg2611,
                 reg2608,
                 reg2605,
                 reg2604,
                 reg2602,
                 reg2599,
                 reg2597,
                 reg2596,
                 reg2594,
                 reg2593,
                 reg2591,
                 reg2590,
                 reg2589,
                 reg2588,
                 reg2586,
                 reg2583,
                 reg2582,
                 reg2580,
                 reg2579,
                 reg2578,
                 reg2577,
                 reg2556,
                 reg2574,
                 reg2573,
                 reg2571,
                 reg2569,
                 reg2567,
                 reg2565,
                 reg2564,
                 reg2562,
                 reg2561,
                 reg2559,
                 reg2558,
                 reg2557,
                 reg2555,
                 reg2553,
                 reg2551,
                 reg2547,
                 reg2545,
                 reg2544,
                 reg2543,
                 reg2542,
                 reg2541,
                 reg2539,
                 reg2538,
                 reg2537,
                 reg2536,
                 reg2531,
                 reg2528,
                 reg2526,
                 reg2525,
                 reg2523,
                 reg2521,
                 reg2520,
                 reg2517,
                 reg2515,
                 reg2510,
                 reg2504,
                 reg2513,
                 reg2507,
                 reg2501,
                 reg2497,
                 reg2495,
                 reg2493,
                 reg2488,
                 reg2487,
                 reg2486,
                 reg2484,
                 reg2480,
                 reg2478,
                 reg2800,
                 reg2798,
                 forvar2794,
                 reg2793,
                 reg2791,
                 reg2784,
                 forvar2782,
                 reg2788,
                 reg2785,
                 forvar2784,
                 reg2782,
                 reg2780,
                 reg2777,
                 reg2774,
                 reg2773,
                 reg2771,
                 reg2769,
                 reg2767,
                 reg2766,
                 reg2760,
                 reg2759,
                 reg2758,
                 reg2756,
                 reg2755,
                 forvar2754,
                 reg2753,
                 reg2752,
                 forvar2748,
                 reg2749,
                 reg2745,
                 reg2741,
                 forvar2740,
                 reg2739,
                 forvar2737,
                 reg2725,
                 reg2736,
                 reg2734,
                 reg2732,
                 reg2728,
                 forvar2725,
                 reg2720,
                 reg2719,
                 reg2715,
                 reg2713,
                 reg2712,
                 reg2711,
                 reg2708,
                 reg2705,
                 reg2703,
                 reg2699,
                 reg2698,
                 reg2697,
                 reg2692,
                 reg2691,
                 reg2689,
                 reg2687,
                 reg2686,
                 reg2683,
                 reg2682,
                 reg2681,
                 reg2680,
                 reg2677,
                 reg2673,
                 reg2672,
                 reg2669,
                 forvar2667,
                 reg2666,
                 forvar2665,
                 reg2661,
                 reg2658,
                 reg2657,
                 reg2653,
                 reg2652,
                 forvar2650,
                 reg2648,
                 forvar2647,
                 reg2645,
                 reg2644,
                 forvar2643,
                 reg2642,
                 reg2639,
                 reg2637,
                 forvar2636,
                 reg2633,
                 reg2632,
                 reg2631,
                 reg2629,
                 reg2628,
                 reg2626,
                 forvar2624,
                 reg2623,
                 reg2622,
                 reg2621,
                 reg2620,
                 reg2619,
                 reg2618,
                 reg2616,
                 reg2612,
                 forvar2610,
                 forvar2609,
                 reg2607,
                 reg2606,
                 reg2603,
                 reg2601,
                 reg2600,
                 forvar2598,
                 reg2595,
                 reg2592,
                 reg2587,
                 reg2585,
                 reg2584,
                 forvar2581,
                 forvar2576,
                 forvar2575,
                 reg2572,
                 reg2570,
                 reg2568,
                 reg2566,
                 reg2563,
                 reg2560,
                 forvar2556,
                 reg2554,
                 reg2552,
                 reg2550,
                 reg2549,
                 forvar2548,
                 reg2546,
                 reg2540,
                 reg2535,
                 reg2534,
                 reg2533,
                 reg2532,
                 reg2530,
                 reg2529,
                 reg2527,
                 reg2524,
                 reg2522,
                 reg2519,
                 reg2518,
                 reg2516,
                 reg2514,
                 reg2512,
                 reg2511,
                 forvar2510,
                 reg2509,
                 reg2508,
                 reg2506,
                 reg2505,
                 forvar2504,
                 reg2503,
                 reg2502,
                 reg2500,
                 forvar2499,
                 reg2498,
                 reg2496,
                 reg2494,
                 reg2492,
                 reg2491,
                 reg2490,
                 reg2489,
                 reg2485,
                 reg2483,
                 reg2482,
                 reg2481,
                 reg2479,
                 reg2477,
                 forvar2476,
                 (1'h0)};
  assign wire2473 = {wire2471,
                        $signed($signed((wire2471[(3'h4):(2'h3)] ?
                            (wire2469 | wire2472) : wire2471[(3'h4):(2'h2)])))};
  assign wire2474 = wire2468[(5'h13):(4'h8)];
  assign wire2475 = wire2470;
  always
    @(posedge clk) begin
      for (forvar2476 = (1'h0); (forvar2476 < (3'h4)); forvar2476 = (forvar2476 + (1'h1)))
        begin
          if ($unsigned((^(($signed((7'h53)) ?
              (wire2473 ~^ wire2471) : (wire2475 ?
                  wire2473 : forvar2476)) >> ((wire2471 ? wire2469 : wire2468) ?
              wire2475 : wire2472)))))
            begin
              reg2477 = wire2470;
              reg2478 <= ($signed((-{{wire2470, wire2471, wire2469},
                      (|(7'h4f))})) ?
                  (wire2473[(1'h1):(1'h1)] != wire2471[(3'h4):(2'h3)]) : wire2470);
              reg2479 = forvar2476[(3'h4):(2'h2)];
            end
          else
            begin
              reg2478 <= {wire2471[(3'h6):(3'h4)],
                  ({forvar2476[(4'hd):(1'h1)],
                      {(wire2469 ? (8'hbe) : wire2469),
                          wire2470[(4'h8):(3'h4)]},
                      wire2469[(4'h9):(1'h0)]} * (&({forvar2476, wire2472} ?
                      (reg2479 ? wire2470 : wire2475) : (wire2470 ?
                          wire2469 : wire2475))))};
              reg2480 <= reg2477[(3'h7):(3'h6)];
              reg2481 = (-(!((-reg2479[(3'h4):(1'h1)]) <= (~^{reg2478,
                  reg2479}))));
              reg2482 = $signed((~reg2479));
              reg2483 = wire2475;
              reg2484 <= $unsigned(reg2482[(4'hb):(2'h2)]);
              reg2485 = $unsigned(reg2480[(2'h2):(2'h2)]);
            end
          reg2486 <= (+(reg2483 ?
              $signed((+(&reg2485))) : reg2484[(5'h12):(3'h4)]));
          if (reg2480[(2'h2):(2'h2)])
            begin
              reg2487 <= (((~^{$unsigned(reg2486)}) - reg2483[(2'h2):(1'h0)]) >= reg2480);
              reg2488 <= ((~^$signed(reg2479)) ^ forvar2476);
              reg2489 = $unsigned({(|($unsigned(reg2486) & reg2478))});
              reg2490 = ((($unsigned(reg2486[(4'hb):(4'ha)]) == ((~wire2470) ?
                          $signed((7'h42)) : $signed(wire2469))) ?
                      wire2470 : wire2470) ?
                  reg2486 : {{wire2468[(4'he):(3'h5)],
                          ((^~wire2471) ?
                              $signed(wire2469) : $unsigned(wire2469)),
                          $unsigned({forvar2476, (8'hb4)})}});
              reg2491 = (~($unsigned((~|(reg2489 ?
                  reg2487 : (8'hb3)))) || (^((wire2472 || wire2470) ?
                  reg2485[(3'h5):(2'h3)] : (8'ha7)))));
              reg2492 = $unsigned({reg2485[(1'h1):(1'h1)]});
              reg2493 <= (|reg2490);
            end
          else
            begin
              reg2489 = ($unsigned(reg2493) <= (reg2478 - $unsigned(({(8'hb6),
                      reg2482} ?
                  reg2478[(4'hb):(2'h3)] : (^~reg2479)))));
              reg2490 = reg2477;
              reg2491 = (&{reg2486, reg2490[(3'h7):(1'h1)]});
              reg2492 = {((^(~|$unsigned(reg2480))) ?
                      ((~$signed(wire2475)) - reg2490) : $signed((8'hb4))),
                  $unsigned(reg2478[(2'h3):(2'h2)])};
              reg2493 <= (~reg2478);
              reg2494 = (~&$unsigned(({$signed(reg2481),
                  reg2481,
                  $signed(reg2480)} >>> $unsigned(wire2473))));
              reg2495 <= ($unsigned((^~wire2471[(1'h1):(1'h0)])) << $signed($signed((+reg2487))));
            end
          reg2496 = ($unsigned($unsigned(wire2468)) | $unsigned(((7'h53) ?
              reg2495 : {reg2480[(1'h1):(1'h0)]})));
          reg2497 <= $signed((&reg2488[(2'h3):(1'h0)]));
          reg2498 = $signed($signed((^~reg2481[(1'h0):(1'h0)])));
          for (forvar2499 = (1'h0); (forvar2499 < (1'h0)); forvar2499 = (forvar2499 + (1'h1)))
            begin
              reg2500 = ($unsigned(($unsigned((reg2487 ?
                      wire2470 : wire2468)) ^~ wire2475)) ?
                  wire2471[(3'h5):(1'h0)] : $signed((reg2496 <= reg2486)));
              reg2501 <= reg2482;
              reg2502 = ((|$signed(((~|reg2501) ? reg2488 : forvar2499))) ?
                  forvar2499[(3'h4):(3'h4)] : ({(~&reg2491),
                      wire2472[(1'h0):(1'h0)],
                      $unsigned((wire2470 ?
                          (8'h9c) : (8'ha8)))} == reg2495[(2'h2):(1'h0)]));
              reg2503 = reg2494;
            end
        end
      if (reg2480)
        begin
          for (forvar2504 = (1'h0); (forvar2504 < (3'h5)); forvar2504 = (forvar2504 + (1'h1)))
            begin
              reg2505 = $unsigned(reg2485);
              reg2506 = $unsigned(reg2485);
              reg2507 <= ({(((reg2503 ?
                          reg2482 : wire2473) != $unsigned((8'ha4))) ~^ {(~reg2479),
                          $signed(wire2474),
                          reg2480})} ?
                  (reg2486[(3'h6):(2'h2)] > (-((8'hb0) ?
                      (~&reg2479) : $signed(wire2475)))) : {wire2475[(4'hb):(3'h4)],
                      reg2505});
              reg2508 = ({$signed((~&$unsigned(reg2501))),
                  (|(-reg2500))} || (~&forvar2504));
              reg2509 = (~|(+$signed((~(reg2486 << forvar2499)))));
            end
          for (forvar2510 = (1'h0); (forvar2510 < (3'h4)); forvar2510 = (forvar2510 + (1'h1)))
            begin
              reg2511 = ((reg2485[(3'h7):(3'h4)] && ((((7'h40) > (8'hb4)) ^ (forvar2499 ?
                  reg2496 : wire2473)) <= $unsigned($signed(reg2502)))) * $unsigned((~{((8'haf) ^ reg2494),
                  $signed(reg2481)})));
              reg2512 = (reg2498[(1'h0):(1'h0)] ?
                  forvar2499[(5'h18):(3'h6)] : reg2489[(5'h16):(4'he)]);
              reg2513 <= ((({(wire2475 & wire2469)} ?
                      ((reg2485 == reg2483) | $unsigned((8'hbb))) : $unsigned((reg2503 ?
                          reg2483 : (7'h57)))) < (reg2487[(2'h2):(1'h1)] ^ (~$unsigned(reg2479)))) ?
                  ($signed(reg2495[(2'h2):(1'h0)]) || reg2488[(2'h2):(1'h0)]) : $signed($unsigned($unsigned(reg2491))));
            end
          reg2514 = reg2485;
        end
      else
        begin
          if ({((((~|reg2481) & $signed(reg2486)) << reg2491[(1'h1):(1'h0)]) << $unsigned(($unsigned((8'had)) ?
                  reg2502[(3'h6):(3'h5)] : (~^reg2507))))})
            begin
              reg2504 <= (reg2489 ?
                  reg2501 : ($unsigned(((^reg2482) ?
                      reg2488[(3'h4):(2'h3)] : ((8'ha5) ?
                          wire2474 : reg2480))) && $signed(reg2509)));
              reg2507 <= reg2478[(4'hb):(3'h5)];
            end
          else
            begin
              reg2504 <= reg2509;
              reg2505 = reg2489;
              reg2507 <= (wire2472[(4'h8):(3'h4)] || (~((reg2487[(1'h1):(1'h1)] || reg2485[(2'h3):(1'h0)]) > $unsigned(reg2494[(4'hd):(4'hb)]))));
              reg2510 <= $unsigned(reg2477[(4'h9):(4'h9)]);
              reg2511 = ({$signed($unsigned($signed((7'h43))))} ?
                  $unsigned(((^~(reg2494 || reg2490)) <<< $unsigned((!reg2487)))) : reg2507);
              reg2512 = {{(reg2512 && reg2489[(2'h2):(2'h2)]),
                      $signed((~$signed(reg2479)))},
                  wire2471};
              reg2513 <= $signed((reg2497[(5'h17):(5'h10)] ?
                  reg2479 : ($signed(reg2481) ?
                      (~^reg2510[(5'h11):(2'h3)]) : (((8'hb8) < reg2482) ^ forvar2499))));
            end
          if (($signed(($unsigned(reg2511) ?
                  (^{reg2478,
                      reg2498}) : ($unsigned(reg2505) * $signed(forvar2504)))) ?
              $unsigned(forvar2504) : (+($signed($unsigned(wire2471)) || $unsigned($unsigned(reg2502))))))
            begin
              reg2514 = (wire2475 ?
                  (reg2506[(5'h14):(2'h3)] ?
                      ((reg2484[(3'h4):(2'h3)] <<< (reg2482 ^~ wire2468)) ?
                          ((reg2482 ? reg2493 : (8'h9c)) ?
                              {reg2477,
                                  (8'hbd)} : reg2484[(5'h13):(4'h8)]) : ((~&reg2484) ?
                              $signed(wire2468) : (reg2491 ?
                                  reg2489 : reg2509))) : forvar2510[(4'hc):(4'h8)]) : reg2512[(5'h14):(4'he)]);
            end
          else
            begin
              reg2515 <= $unsigned({$signed((((8'ha4) ?
                      forvar2510 : reg2484) & (8'had))),
                  wire2471,
                  ($signed((wire2474 & reg2485)) || reg2513[(5'h16):(5'h10)])});
              reg2516 = (+reg2505);
              reg2517 <= reg2479;
              reg2518 = (((^~{(wire2474 ? reg2491 : reg2514),
                  reg2477[(4'h9):(4'h8)]}) || ((|{wire2473,
                  (8'hba)}) == wire2473[(3'h5):(3'h5)])) < (reg2485 ?
                  $signed((^~$signed(reg2509))) : (reg2492 * (reg2484[(4'h8):(1'h0)] && $signed(reg2517)))));
              reg2519 = reg2516;
              reg2520 <= reg2482;
              reg2521 <= $unsigned($signed((reg2516[(5'h13):(3'h5)] ^ reg2520)));
            end
          reg2522 = $signed($signed(((!(reg2506 << forvar2510)) < wire2468)));
          reg2523 <= $signed(reg2492);
          if ((~^($signed($signed((!(8'hb2)))) ?
              $unsigned(((wire2473 ? (8'hbe) : reg2488) ?
                  $unsigned(wire2470) : reg2481)) : $signed(({reg2492} ?
                  (8'ha6) : (+reg2498))))))
            begin
              reg2524 = reg2492[(5'h15):(4'hf)];
              reg2525 <= {reg2486[(4'hb):(3'h7)],
                  {$unsigned(wire2468),
                      $unsigned(($signed(reg2485) - (reg2487 ?
                          reg2497 : reg2498)))}};
              reg2526 <= (~|$unsigned($unsigned((&reg2495[(1'h1):(1'h0)]))));
              reg2527 = reg2493[(4'h9):(3'h7)];
            end
          else
            begin
              reg2525 <= reg2486[(4'he):(4'hd)];
              reg2526 <= $signed($unsigned($signed($unsigned(reg2501))));
              reg2528 <= (~^(~^reg2498[(5'h1c):(2'h3)]));
              reg2529 = (+(forvar2476 ?
                  wire2468[(3'h7):(3'h6)] : (((^(7'h54)) ?
                      (reg2479 ?
                          wire2473 : reg2512) : reg2491) >> $unsigned(forvar2510[(5'h1c):(5'h1b)]))));
            end
          if ($signed(($signed(wire2475[(2'h3):(1'h0)]) <= reg2497)))
            begin
              reg2530 = $unsigned($unsigned((reg2504[(4'h9):(3'h4)] ?
                  ((reg2486 << reg2510) ?
                      {reg2517,
                          wire2475,
                          reg2489} : reg2500[(3'h6):(1'h0)]) : (-$signed(reg2489)))));
            end
          else
            begin
              reg2530 = ((($signed($signed(reg2488)) ?
                      $unsigned((+reg2513)) : (-(&(7'h56)))) >= {((7'h48) ?
                          {reg2528, reg2495} : reg2530),
                      reg2529}) ?
                  $unsigned(reg2527[(5'h1a):(5'h15)]) : ($unsigned(((~^reg2483) ?
                      $signed(reg2527) : $unsigned(reg2492))) | forvar2476));
              reg2531 <= wire2475[(3'h6):(2'h3)];
            end
        end
      if ($unsigned({$signed(((8'hae) ?
              ((7'h45) ~^ (8'hae)) : $signed(reg2479))),
          $unsigned(((reg2478 ? (8'hbd) : reg2496) ?
              reg2495[(1'h0):(1'h0)] : $signed((7'h4b))))}))
        begin
          reg2532 = reg2503;
          reg2533 = reg2520[(5'h16):(5'h16)];
          reg2534 = reg2495;
          reg2535 = $signed(reg2494);
        end
      else
        begin
          reg2532 = ($signed(reg2477[(1'h0):(1'h0)]) ?
              forvar2510[(5'h1a):(5'h11)] : ($unsigned(reg2522[(3'h4):(1'h1)]) == (forvar2499[(5'h10):(4'h9)] ?
                  reg2514 : (!reg2534[(4'hc):(4'hc)]))));
          if ($unsigned(wire2469))
            begin
              reg2536 <= reg2488[(2'h3):(1'h1)];
            end
          else
            begin
              reg2533 = $unsigned(((((reg2517 ? reg2491 : reg2492) ?
                  (reg2478 ? (8'hb3) : (7'h51)) : (reg2531 ?
                      reg2482 : wire2471)) ~^ $signed(reg2503[(3'h6):(1'h0)])) <<< {$unsigned({reg2511})}));
              reg2536 <= (forvar2510[(5'h11):(5'h11)] - $signed((-$signed((reg2528 ?
                  (7'h40) : reg2508)))));
              reg2537 <= $signed($unsigned(({reg2509[(3'h7):(1'h1)],
                      (-reg2498)} ?
                  (reg2502[(5'h10):(2'h3)] ?
                      (reg2496 ?
                          reg2510 : reg2486) : reg2535[(4'h9):(3'h4)]) : $signed($unsigned(reg2478)))));
              reg2538 <= $signed(reg2485[(1'h1):(1'h1)]);
              reg2539 <= (~|($signed((~$signed(reg2537))) ?
                  $unsigned(($unsigned(reg2495) << $signed(reg2524))) : {({reg2525} ?
                          (~&reg2522) : $signed(reg2502))}));
              reg2540 = (reg2525 << (+(|$signed(reg2478[(4'hc):(2'h2)]))));
              reg2541 <= $signed((^(~^(-reg2536[(2'h2):(2'h2)]))));
            end
          reg2542 <= reg2486;
          reg2543 <= $signed(reg2484);
          if (reg2519[(4'he):(3'h7)])
            begin
              reg2544 <= ((-(reg2494[(4'h8):(3'h4)] == reg2482[(4'ha):(3'h4)])) >>> (^~(((reg2492 ?
                          (7'h42) : reg2496) ?
                      reg2534 : $unsigned(reg2478)) ?
                  (!$unsigned(reg2511)) : (~&(reg2536 <= reg2497)))));
              reg2545 <= reg2527;
            end
          else
            begin
              reg2546 = reg2525[(4'hb):(4'hb)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg2547 <= $unsigned((7'h52));
      if ({$signed(((8'ha7) ? reg2488 : $signed({reg2515, reg2531, (8'hbe)})))})
        begin
          for (forvar2548 = (1'h0); (forvar2548 < (3'h6)); forvar2548 = (forvar2548 + (1'h1)))
            begin
              reg2549 = reg2513;
              reg2550 = (reg2521 * $unsigned((&{reg2486[(2'h2):(1'h0)],
                  {(7'h4d), reg2528},
                  $unsigned((8'h9f))})));
              reg2551 <= (((reg2539[(4'h8):(2'h3)] ?
                      ({reg2528} & $unsigned(reg2484)) : wire2475[(1'h1):(1'h0)]) >>> (&$signed((reg2526 ?
                      (8'hbc) : (7'h53))))) ?
                  (^~$unsigned($unsigned(reg2497[(4'hd):(2'h2)]))) : $signed(((^reg2504) ~^ (-(reg2539 >>> reg2531)))));
              reg2552 = $signed(($unsigned($unsigned((~|reg2542))) ?
                  {((8'hb7) == (-reg2523)),
                      ($unsigned(reg2544) && reg2497[(4'h9):(3'h5)]),
                      (reg2504[(3'h5):(2'h3)] ^~ reg2523[(1'h1):(1'h0)])} : (|reg2537[(2'h3):(2'h2)])));
              reg2553 <= reg2484;
              reg2554 = $unsigned($unsigned($signed(((reg2543 ?
                  reg2549 : reg2488) <<< (^reg2552)))));
              reg2555 <= reg2504[(4'hf):(4'hb)];
            end
          for (forvar2556 = (1'h0); (forvar2556 < (1'h1)); forvar2556 = (forvar2556 + (1'h1)))
            begin
              reg2557 <= ($unsigned($signed($unsigned($unsigned(reg2553)))) <= (($unsigned((reg2541 ?
                      (8'ha6) : reg2486)) ?
                  ((-wire2472) ?
                      $unsigned(wire2470) : {reg2536,
                          reg2539}) : $unsigned(reg2487)) & forvar2548));
              reg2558 <= (reg2555[(2'h2):(1'h1)] == $unsigned(((reg2520 ?
                      ((8'hb2) + (8'hbc)) : reg2510[(4'hf):(4'ha)]) ?
                  ((&(8'haf)) ? $signed(forvar2548) : (~&(8'haa))) : ((reg2528 ?
                      reg2521 : reg2526) | (~^reg2550)))));
              reg2559 <= $signed(((~^({wire2470,
                      (8'hb8),
                      forvar2556} > $unsigned(reg2487))) ?
                  {reg2526} : $signed(((!wire2471) ?
                      ((7'h4c) >>> reg2497) : $signed(reg2478)))));
              reg2560 = (!($signed(reg2510) ?
                  $unsigned(reg2486[(4'ha):(4'h9)]) : (reg2487[(1'h0):(1'h0)] ?
                      $signed((reg2507 ?
                          reg2558 : reg2507)) : $unsigned({(7'h48),
                          reg2536,
                          reg2551}))));
              reg2561 <= $signed(($unsigned($signed(reg2539)) ?
                  (~reg2552[(3'h4):(1'h1)]) : $signed($signed((|(8'ha7))))));
            end
          if (((~($signed((reg2486 ? (7'h4c) : reg2495)) ?
                  ($signed(reg2507) ?
                      $signed(wire2473) : (reg2558 & reg2558)) : ((reg2531 ?
                          reg2510 : wire2471) ?
                      (-(8'hb8)) : reg2543[(1'h1):(1'h1)]))) ?
              (reg2541[(5'h12):(2'h3)] > (+reg2531)) : $signed($unsigned({(reg2542 | reg2497)}))))
            begin
              reg2562 <= (reg2486 >>> $unsigned({$signed((reg2554 * reg2550)),
                  (|(7'h44)),
                  $signed((reg2484 >= reg2557))}));
              reg2563 = (^(8'hb3));
              reg2564 <= ($signed(($unsigned($signed(reg2557)) ?
                      (8'hbc) : {reg2543[(2'h3):(1'h1)],
                          $signed(reg2513),
                          (~&wire2470)})) ?
                  ((reg2560[(2'h2):(1'h0)] ?
                      ((&wire2469) ^ $unsigned((8'haa))) : ($signed((8'ha7)) ?
                          (~^(7'h48)) : reg2547)) || $unsigned({(reg2538 ?
                          reg2501 : reg2501),
                      $signed(reg2484),
                      ((7'h4c) + reg2559)})) : (-((~^$unsigned(reg2517)) + reg2513)));
              reg2565 <= reg2563[(2'h2):(1'h1)];
              reg2566 = {{((8'had) ^ $unsigned(wire2471)),
                      reg2493[(4'hb):(4'hb)],
                      (^~((reg2515 ?
                          reg2521 : reg2549) ^ (reg2523 <<< reg2549)))},
                  ($unsigned(reg2493[(5'h16):(5'h16)]) || (~&(((7'h4a) <= reg2501) <<< (wire2474 ?
                      (8'h9f) : reg2488)))),
                  {reg2487, {reg2549, reg2562}}};
            end
          else
            begin
              reg2562 <= $signed(reg2487);
              reg2563 = (reg2542[(3'h4):(1'h1)] ?
                  (~^$unsigned((reg2513[(2'h2):(2'h2)] == (!forvar2556)))) : reg2515);
              reg2564 <= $unsigned({($unsigned(reg2517[(4'h9):(4'h8)]) * reg2566)});
            end
          if ((($signed(reg2545) & $unsigned((-(!reg2547)))) - (~^reg2552)))
            begin
              reg2567 <= {reg2557[(5'h13):(3'h6)],
                  $unsigned((reg2549 >> reg2559)),
                  ((^~$unsigned({wire2468})) ?
                      ($signed($unsigned(reg2539)) ?
                          reg2542[(4'h8):(1'h0)] : $unsigned($unsigned(reg2497))) : (({reg2507,
                                  reg2528} ?
                              $signed(reg2555) : (7'h42)) ?
                          (~|{wire2470}) : ({(8'hbf),
                              wire2469} ~^ (reg2493 <<< reg2520))))};
              reg2568 = $signed(reg2555);
              reg2569 <= $signed(((~&reg2528[(4'he):(3'h7)]) && (8'hae)));
              reg2570 = $signed((7'h46));
            end
          else
            begin
              reg2567 <= $signed((-reg2567[(5'h19):(4'ha)]));
              reg2569 <= (!(8'ha6));
              reg2571 <= ($signed(((&$signed(reg2550)) ?
                  ($unsigned(reg2528) == (wire2472 ?
                      reg2517 : (8'haf))) : reg2552[(2'h3):(2'h3)])) <= reg2531);
              reg2572 = (reg2557 * wire2474);
              reg2573 <= wire2475[(5'h19):(3'h4)];
            end
          reg2574 <= reg2554;
        end
      else
        begin
          for (forvar2548 = (1'h0); (forvar2548 < (3'h4)); forvar2548 = (forvar2548 + (1'h1)))
            begin
              reg2551 <= ((~(((reg2547 ^ wire2475) - {reg2554,
                      reg2478}) || $signed(reg2501[(3'h4):(1'h0)]))) ?
                  reg2486[(2'h2):(1'h0)] : $signed(reg2557));
              reg2553 <= (~&$unsigned((7'h4d)));
              reg2555 <= forvar2556;
              reg2556 <= $signed({(reg2537[(2'h3):(2'h2)] ~^ ($signed(reg2555) * (!reg2547))),
                  (^~reg2570[(3'h5):(3'h4)])});
              reg2557 <= (~|(reg2560[(3'h6):(3'h4)] ?
                  (^((8'hac) ?
                      (reg2480 ~^ reg2559) : (reg2549 ?
                          reg2570 : (8'hba)))) : (~|(reg2558[(4'hc):(3'h4)] == {reg2574}))));
              reg2560 = (~|(reg2563[(1'h0):(1'h0)] ?
                  ((wire2469 == (~^(8'hb5))) ?
                      {$unsigned(reg2547),
                          $signed(reg2556),
                          (wire2473 & wire2468)} : ($signed(reg2561) <<< $unsigned(wire2471))) : {reg2545[(1'h1):(1'h1)],
                      {$unsigned(reg2565)}}));
            end
          reg2561 <= reg2484;
          reg2562 <= reg2510[(4'hf):(4'hb)];
          if (reg2478)
            begin
              reg2563 = reg2564[(5'h15):(4'hd)];
              reg2564 <= (($signed(((reg2557 + (8'hba)) | {reg2507,
                      wire2472,
                      reg2558})) ^~ reg2536) ?
                  (reg2526 ?
                      $unsigned(reg2563) : forvar2548) : (|((^~{wire2472}) * wire2468[(4'hc):(1'h1)])));
              reg2566 = reg2552[(1'h1):(1'h0)];
              reg2567 <= reg2488[(2'h3):(2'h2)];
              reg2569 <= (~(+(~reg2563)));
              reg2570 = reg2495;
              reg2571 <= reg2554[(3'h5):(3'h5)];
            end
          else
            begin
              reg2564 <= (|reg2553[(3'h4):(2'h3)]);
              reg2565 <= (reg2572[(1'h0):(1'h0)] ?
                  $signed((({reg2510, reg2564} >= (reg2557 ^ reg2531)) ?
                      (7'h45) : reg2564)) : reg2538[(3'h5):(1'h1)]);
              reg2566 = ((reg2507 ?
                      reg2515 : (($unsigned(reg2569) ?
                          $signed(wire2475) : reg2557[(5'h11):(2'h2)]) || ($unsigned(reg2562) ?
                          reg2556[(2'h2):(1'h0)] : reg2547[(4'ha):(1'h0)]))) ?
                  reg2484[(4'hd):(3'h4)] : (|$signed((reg2528[(4'h9):(2'h3)] ?
                      ((8'hbb) ? wire2473 : reg2521) : {(7'h4e)}))));
              reg2567 <= wire2471;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2575 = (1'h0); (forvar2575 < (3'h4)); forvar2575 = (forvar2575 + (1'h1)))
        begin
          for (forvar2576 = (1'h0); (forvar2576 < (3'h5)); forvar2576 = (forvar2576 + (1'h1)))
            begin
              reg2577 <= $unsigned($unsigned((8'ha2)));
              reg2578 <= $unsigned((reg2551 * ($signed($signed(reg2561)) ?
                  forvar2576[(1'h0):(1'h0)] : $signed((|reg2515)))));
            end
          reg2579 <= reg2547;
          reg2580 <= reg2523;
          for (forvar2581 = (1'h0); (forvar2581 < (1'h1)); forvar2581 = (forvar2581 + (1'h1)))
            begin
              reg2582 <= ($signed({$signed((reg2480 >> (7'h4b)))}) ?
                  (($signed($unsigned(reg2577)) ?
                      (8'hbb) : $signed($signed(forvar2575))) >= ((8'hb1) != reg2556)) : (~^(+($unsigned(reg2567) << reg2559))));
              reg2583 <= (reg2551[(1'h0):(1'h0)] ?
                  (reg2553[(3'h7):(1'h0)] ?
                      ({$signed(reg2565),
                          (reg2557 && reg2565)} >= ((reg2571 * reg2538) ?
                          $unsigned(reg2580) : (~|reg2501))) : (|reg2541[(5'h10):(4'h9)])) : reg2520[(3'h4):(3'h4)]);
              reg2584 = $signed(($signed((^~{(7'h4d), reg2547})) ?
                  $signed(reg2513[(4'hc):(4'h9)]) : reg2501));
              reg2585 = (~reg2556);
              reg2586 <= ($signed(reg2478) ?
                  ($unsigned((~&(~^reg2573))) >= reg2488[(1'h0):(1'h0)]) : (&$signed(((^forvar2581) & (8'ha4)))));
            end
          if (($unsigned(($unsigned((wire2468 <= reg2565)) ?
                  (!$unsigned(reg2513)) : ((^reg2578) == $signed(reg2545)))) ?
              (~&reg2513[(4'h9):(3'h7)]) : (reg2579[(4'h9):(4'h8)] == reg2567[(2'h3):(1'h1)])))
            begin
              reg2587 = $unsigned(reg2579);
              reg2588 <= forvar2575;
              reg2589 <= $unsigned((7'h4d));
              reg2590 <= ((~&reg2547) && (|(8'hb0)));
              reg2591 <= reg2488;
              reg2592 = ($unsigned({((reg2536 ^~ reg2583) < {wire2468}),
                  $unsigned((reg2565 ?
                      forvar2575 : wire2472))}) ~^ (~&$signed(reg2589[(2'h2):(1'h1)])));
            end
          else
            begin
              reg2588 <= ((((~|{reg2539, (8'ha4), reg2555}) ?
                  ((~^reg2488) ?
                      (reg2569 ?
                          (7'h4b) : reg2556) : (wire2470 <<< reg2567)) : $signed((-reg2493))) >>> {$signed((~&reg2558)),
                  $signed(reg2557),
                  ({reg2536,
                      (8'hab)} * (reg2562 >> reg2478))}) != ({$unsigned((reg2569 ?
                          reg2542 : reg2537))} ?
                  reg2501 : wire2474));
              reg2589 <= {$unsigned(($signed(reg2536[(1'h0):(1'h0)]) || ((reg2565 == reg2567) ?
                      wire2473 : (reg2531 ? reg2504 : reg2584)))),
                  ((wire2473 == (~|$unsigned(reg2571))) ? wire2475 : wire2471)};
              reg2592 = reg2557[(5'h18):(5'h13)];
              reg2593 <= reg2510;
              reg2594 <= (~^reg2567);
              reg2595 = {reg2510[(4'hf):(1'h1)]};
              reg2596 <= reg2521;
            end
          reg2597 <= wire2473[(3'h7):(2'h2)];
          for (forvar2598 = (1'h0); (forvar2598 < (2'h3)); forvar2598 = (forvar2598 + (1'h1)))
            begin
              reg2599 <= $unsigned(reg2553);
              reg2600 = forvar2581;
              reg2601 = wire2468[(4'h9):(3'h5)];
              reg2602 <= (~wire2472);
              reg2603 = (reg2517 == ((((forvar2576 >>> (8'ha9)) ?
                      reg2590[(4'h8):(1'h1)] : $signed(reg2579)) ?
                  ((~&reg2600) ?
                      $unsigned(reg2558) : $unsigned(reg2558)) : (((7'h4e) ?
                          reg2544 : (7'h41)) ?
                      (7'h42) : reg2578)) + $unsigned((8'ha3))));
              reg2604 <= reg2484[(5'h17):(4'h8)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg2605 <= ($signed((7'h4f)) ?
          ({($signed(reg2488) - (reg2545 >> reg2559))} > reg2555) : reg2501[(1'h1):(1'h0)]);
      reg2606 = $signed(reg2578[(5'h11):(5'h10)]);
      reg2607 = (wire2468[(4'h8):(4'h8)] ? reg2525 : (&reg2588[(3'h4):(2'h3)]));
      reg2608 <= reg2545[(5'h1d):(4'hb)];
    end
  always
    @(posedge clk) begin
      for (forvar2609 = (1'h0); (forvar2609 < (2'h2)); forvar2609 = (forvar2609 + (1'h1)))
        begin
          for (forvar2610 = (1'h0); (forvar2610 < (3'h5)); forvar2610 = (forvar2610 + (1'h1)))
            begin
              reg2611 <= reg2543;
              reg2612 = $signed((|reg2507));
              reg2613 <= ($unsigned(reg2580) ?
                  reg2557 : $unsigned((((&reg2580) ?
                      reg2556 : $signed(reg2590)) & $signed((^(7'h56))))));
              reg2614 <= $signed((reg2538[(4'h9):(2'h2)] <<< $unsigned((^~reg2561))));
              reg2615 <= (reg2612 ?
                  $signed(($signed({(7'h46)}) + (-(reg2547 <<< (8'ha4))))) : $unsigned(reg2583));
              reg2616 = reg2513;
              reg2617 <= $unsigned(reg2597[(5'h14):(4'h8)]);
            end
          reg2618 = reg2612;
          reg2619 = (+(reg2521 <= $signed((reg2613[(3'h7):(2'h2)] ?
              $signed((8'ha9)) : $unsigned(reg2521)))));
          reg2620 = (((reg2521[(2'h2):(1'h0)] <= (^~$unsigned(reg2604))) << {reg2619[(5'h15):(5'h11)],
              {$signed(reg2484), {reg2493, reg2564, reg2542}}}) & (^reg2501));
          reg2621 = $unsigned(({$unsigned((~&(7'h4c))),
              $signed(((7'h4c) ? reg2507 : reg2537))} | forvar2609));
          reg2622 = ($signed((|((7'h4a) ?
              reg2528 : reg2558[(5'h12):(4'he)]))) == ({(reg2569[(5'h12):(1'h1)] ?
                      $unsigned((7'h43)) : (|reg2536)),
                  reg2544[(3'h7):(3'h5)]} ?
              $signed((wire2468[(4'h9):(1'h0)] < {reg2617,
                  reg2569})) : $signed(reg2561[(4'hd):(4'hc)])));
        end
      reg2623 = $signed((~($signed($unsigned((7'h46))) - (+wire2468))));
      for (forvar2624 = (1'h0); (forvar2624 < (3'h4)); forvar2624 = (forvar2624 + (1'h1)))
        begin
          reg2625 <= (reg2558 ?
              ($signed($signed((reg2589 ? forvar2609 : reg2507))) ?
                  ($signed({reg2553,
                      reg2577}) >> reg2617) : (reg2484[(2'h3):(1'h1)] ?
                      (~(reg2478 <<< reg2480)) : (7'h4b))) : reg2515);
          reg2626 = $signed(((-$unsigned((reg2599 ?
              (8'h9c) : reg2618))) && forvar2624));
          if ($unsigned(reg2582[(2'h3):(2'h3)]))
            begin
              reg2627 <= ((^reg2515[(1'h1):(1'h1)]) ^~ $signed((|$signed((~^reg2542)))));
              reg2628 = (^reg2544);
              reg2629 = {reg2564,
                  (($signed({(8'hb3)}) ?
                      reg2608[(3'h4):(2'h3)] : (7'h56)) > (^~{{wire2469,
                          reg2623,
                          reg2579}})),
                  $signed((!((~reg2618) <<< (reg2556 ?
                      reg2562 : forvar2609))))};
              reg2630 <= $signed((reg2620[(4'ha):(3'h5)] ?
                  (~$unsigned($signed(reg2629))) : (reg2561[(2'h2):(2'h2)] <<< wire2473[(1'h0):(1'h0)])));
            end
          else
            begin
              reg2627 <= ($signed((-$unsigned($unsigned(reg2571)))) ?
                  {((~&reg2555[(3'h4):(1'h1)]) ?
                          ((reg2515 ? reg2544 : (7'h4f)) ?
                              {reg2586,
                                  reg2488,
                                  wire2469} : reg2577) : (^wire2470)),
                      reg2593[(4'ha):(4'h9)]} : (((reg2517[(1'h1):(1'h0)] != reg2591) ?
                      reg2564[(5'h17):(4'hf)] : reg2613[(3'h6):(1'h0)]) != reg2613));
              reg2628 = $signed((wire2469[(1'h0):(1'h0)] ?
                  $signed(((forvar2610 != reg2616) ?
                      reg2578[(4'hc):(4'h9)] : (reg2517 && reg2622))) : (+(~reg2593[(4'hc):(1'h1)]))));
              reg2630 <= $signed(($signed(reg2556) >>> reg2537[(3'h4):(2'h3)]));
              reg2631 = $unsigned($signed(($signed((|reg2521)) | {reg2504[(1'h1):(1'h0)],
                  (reg2605 ? (8'hbd) : reg2526),
                  (reg2531 ? (8'haa) : reg2517)})));
              reg2632 = $unsigned((8'hb9));
            end
          if ((~&$signed(reg2537)))
            begin
              reg2633 = ((!reg2486[(2'h3):(2'h3)]) ?
                  $signed((-(7'h4d))) : (&(^~reg2602)));
              reg2634 <= reg2591;
              reg2635 <= $signed(reg2630[(5'h17):(1'h0)]);
            end
          else
            begin
              reg2633 = reg2542;
            end
        end
      for (forvar2636 = (1'h0); (forvar2636 < (1'h1)); forvar2636 = (forvar2636 + (1'h1)))
        begin
          reg2637 = reg2542[(3'h4):(2'h2)];
          reg2638 <= $signed(({reg2488[(2'h3):(2'h2)]} - reg2567[(4'h9):(3'h6)]));
        end
      reg2639 = $signed((&wire2474[(4'hd):(3'h4)]));
    end
  assign wire2640 = {reg2588,
                        (reg2558 >>> reg2544[(3'h6):(2'h2)]),
                        (~|(reg2537[(3'h6):(3'h6)] ?
                            wire2468[(5'h11):(4'h9)] : (!((7'h57) ?
                                wire2472 : reg2583))))};
  always
    @(posedge clk) begin
      reg2641 <= reg2602[(3'h4):(2'h2)];
      reg2642 = reg2573;
      for (forvar2643 = (1'h0); (forvar2643 < (2'h3)); forvar2643 = (forvar2643 + (1'h1)))
        begin
          reg2644 = ((8'ha2) + reg2556);
          reg2645 = $signed(reg2597);
          reg2646 <= ($signed($unsigned($unsigned(reg2565[(3'h6):(2'h3)]))) ?
              reg2591[(4'h9):(1'h1)] : {reg2525[(4'h8):(3'h5)]});
          for (forvar2647 = (1'h0); (forvar2647 < (1'h0)); forvar2647 = (forvar2647 + (1'h1)))
            begin
              reg2648 = reg2515;
              reg2649 <= reg2605[(3'h6):(3'h5)];
            end
          for (forvar2650 = (1'h0); (forvar2650 < (3'h4)); forvar2650 = (forvar2650 + (1'h1)))
            begin
              reg2651 <= ((8'hbe) ?
                  ($unsigned({wire2469}) & (~^reg2613)) : reg2531[(1'h1):(1'h0)]);
              reg2652 = {reg2579};
              reg2653 = reg2539[(5'h14):(4'hb)];
              reg2654 <= reg2615[(2'h2):(1'h0)];
            end
          if ((^$unsigned(($signed(reg2608) == ($unsigned(reg2579) || (reg2488 ?
              reg2531 : reg2635))))))
            begin
              reg2655 <= (8'hb3);
              reg2656 <= {reg2567,
                  $signed($signed($signed($signed(reg2580)))),
                  reg2493[(5'h15):(4'h8)]};
              reg2657 = (^~$unsigned((^~{{reg2656}})));
              reg2658 = reg2577[(1'h0):(1'h0)];
            end
          else
            begin
              reg2655 <= (~^reg2513);
              reg2656 <= (((&reg2590[(2'h2):(1'h0)]) ?
                      reg2565[(4'h9):(1'h1)] : ($signed($signed(reg2648)) ?
                          reg2537[(1'h0):(1'h0)] : {reg2501,
                              (reg2642 ? reg2590 : reg2523)})) ?
                  (reg2582[(1'h1):(1'h0)] ?
                      ((reg2495[(1'h0):(1'h0)] >> (reg2656 >= reg2478)) ?
                          reg2590[(1'h1):(1'h0)] : {$signed(reg2617),
                              (reg2523 >= reg2515)}) : (^~$signed((reg2657 ?
                          reg2615 : reg2602)))) : {(reg2641[(1'h1):(1'h0)] > (~|(7'h45)))});
              reg2657 = {(reg2538 >> (-$signed((reg2593 ? reg2641 : (8'h9c))))),
                  $signed(($signed(reg2605) - reg2541[(4'h8):(1'h0)]))};
              reg2659 <= $unsigned((~^(|$signed((reg2648 ?
                  reg2638 : reg2613)))));
              reg2660 <= (~($unsigned(reg2641[(3'h4):(1'h0)]) >> (7'h42)));
            end
          reg2661 = ((wire2474[(4'he):(3'h6)] ?
                  $signed(reg2605[(1'h1):(1'h1)]) : (reg2635 + reg2590)) ?
              ($unsigned($unsigned(reg2487)) ?
                  ((|(reg2644 ~^ reg2523)) ?
                      ({reg2608,
                          reg2571} ^ $unsigned(reg2520)) : reg2602[(3'h5):(2'h2)]) : $signed((^(reg2579 ?
                      (8'hbb) : reg2590)))) : reg2517[(1'h0):(1'h0)]);
        end
    end
  assign wire2662 = (reg2656[(1'h1):(1'h0)] ~^ ((8'hbc) == $unsigned(($signed(reg2635) ?
                        {reg2586, reg2510} : $signed(reg2545)))));
  assign wire2663 = reg2504;
  assign wire2664 = (-$signed((((!wire2472) ^ ((7'h4e) ? reg2544 : wire2469)) ?
                        $signed(((7'h53) ? wire2473 : reg2578)) : reg2545)));
  always
    @(posedge clk) begin
      for (forvar2665 = (1'h0); (forvar2665 < (2'h2)); forvar2665 = (forvar2665 + (1'h1)))
        begin
          reg2666 = (reg2510[(4'ha):(1'h0)] < (7'h49));
          for (forvar2667 = (1'h0); (forvar2667 < (3'h5)); forvar2667 = (forvar2667 + (1'h1)))
            begin
              reg2668 <= reg2617[(3'h7):(3'h5)];
              reg2669 = reg2545[(5'h16):(1'h0)];
              reg2670 <= reg2590;
              reg2671 <= reg2646;
              reg2672 = (($unsigned({(reg2541 > reg2564), $signed(reg2608)}) ?
                      (((reg2555 ? wire2664 : reg2582) ?
                          $unsigned(reg2578) : ((7'h55) ~^ (7'h4a))) <<< reg2553) : reg2484[(4'hc):(4'hb)]) ?
                  ((~wire2474) * ((+reg2599[(3'h5):(1'h1)]) << reg2571[(5'h12):(1'h1)])) : wire2468[(4'hc):(4'hb)]);
              reg2673 = (&$signed(reg2597));
            end
          if (reg2495[(2'h3):(1'h1)])
            begin
              reg2674 <= (~|(&($unsigned(reg2589) ^ $signed($unsigned((7'h4b))))));
              reg2675 <= {reg2641, reg2625};
              reg2676 <= (reg2651[(2'h2):(2'h2)] ?
                  {{$signed((^~reg2669))}} : reg2589);
              reg2677 = ($signed(reg2553[(3'h6):(3'h4)]) + ($unsigned({(wire2663 != reg2536),
                      reg2520,
                      wire2640}) ?
                  (~|reg2599[(3'h6):(3'h4)]) : wire2471[(2'h3):(2'h2)]));
              reg2678 <= $unsigned($signed(($signed(reg2666[(3'h6):(1'h1)]) >> ($unsigned((8'hb7)) ?
                  (reg2525 ? wire2468 : reg2574) : (reg2571 + reg2520)))));
              reg2679 <= ({({$signed((7'h43))} ?
                      $unsigned((reg2627 ?
                          reg2651 : reg2617)) : reg2588[(2'h3):(2'h2)]),
                  ($signed($unsigned(reg2567)) ?
                      ($signed(reg2480) ?
                          $unsigned(reg2559) : (reg2526 - reg2513)) : $unsigned((reg2654 ?
                          reg2497 : (7'h45))))} >= reg2634[(4'hd):(3'h6)]);
              reg2680 = reg2611;
            end
          else
            begin
              reg2674 <= reg2677[(4'hc):(4'hb)];
            end
          reg2681 = wire2640[(1'h0):(1'h0)];
          if (reg2495[(1'h0):(1'h0)])
            begin
              reg2682 = (reg2676 ?
                  reg2582 : ($signed($signed({reg2673,
                      reg2675,
                      wire2664})) + reg2558));
              reg2683 = {(&$unsigned((~|reg2670))),
                  wire2663[(3'h6):(1'h1)],
                  ($unsigned({wire2469}) ? reg2526 : (8'hb5))};
              reg2684 <= reg2672;
              reg2685 <= $unsigned(reg2604);
            end
          else
            begin
              reg2682 = $signed($unsigned($unsigned((reg2630 ?
                  $unsigned(reg2531) : (reg2551 + reg2525)))));
              reg2684 <= $signed($signed(reg2651));
              reg2686 = ((!(&$signed((reg2567 ? reg2654 : (7'h55))))) ?
                  reg2677[(2'h3):(1'h0)] : reg2523[(2'h2):(1'h0)]);
              reg2687 = ($signed((reg2495 ?
                  (-(~^(8'hb8))) : reg2577)) <<< {wire2472[(2'h3):(2'h3)],
                  (reg2673 << {(reg2531 && reg2668)})});
              reg2688 <= reg2582[(2'h2):(1'h1)];
            end
        end
      reg2689 = reg2611;
      reg2690 <= $signed((~|((reg2493[(5'h1a):(4'hc)] ?
              wire2473 : reg2520[(5'h19):(5'h16)]) ?
          ((reg2504 ?
              reg2556 : reg2680) != reg2649) : $signed(((7'h44) <= reg2545)))));
      reg2691 = $signed((~^wire2470[(2'h3):(2'h2)]));
    end
  always
    @(posedge clk) begin
      reg2692 = wire2469;
      reg2693 <= $signed((reg2655[(3'h7):(3'h5)] < reg2495));
    end
  assign wire2694 = reg2635[(2'h2):(1'h1)];
  assign wire2695 = (($signed($signed((&(8'ha5)))) * $signed(({reg2531,
                                reg2486} ?
                            $signed(reg2605) : (reg2671 ?
                                (7'h47) : reg2488)))) ?
                        $signed(((7'h57) && reg2520)) : reg2523[(1'h0):(1'h0)]);
  assign wire2696 = (|reg2573[(5'h11):(4'hc)]);
  always
    @(posedge clk) begin
      reg2697 = (wire2694[(4'hf):(2'h3)] ?
          (~|reg2569[(2'h3):(1'h0)]) : (-reg2611));
      reg2698 = (reg2693 == reg2646[(4'ha):(2'h3)]);
      if (reg2536[(2'h3):(1'h1)])
        begin
          reg2699 = ((8'hb9) ?
              {(reg2495 ? (~|{reg2551}) : reg2593)} : (((^{reg2515,
                  reg2557,
                  reg2597}) || $signed(reg2536)) == $unsigned(({reg2526,
                      reg2659,
                      reg2693} ?
                  reg2544[(3'h6):(2'h2)] : {(8'ha8), reg2551, reg2605}))));
          reg2700 <= $signed((!$signed((reg2567[(5'h19):(4'hf)] - wire2662[(3'h7):(1'h1)]))));
          reg2701 <= wire2694;
          if ((reg2543[(4'h9):(4'h8)] - ((({reg2660} ?
                      (reg2604 ? reg2542 : wire2471) : {wire2695, reg2596}) ?
                  ({reg2562, reg2487, (7'h4d)} ?
                      (reg2573 ?
                          reg2668 : reg2544) : (wire2695 && reg2517)) : (-(~&reg2537))) ?
              reg2700 : $signed($signed((~|reg2569))))))
            begin
              reg2702 <= $signed($unsigned((+(~^(reg2556 - reg2520)))));
              reg2703 = (8'ha7);
              reg2704 <= reg2675;
              reg2705 = ($signed($unsigned(((|(8'ha4)) - {(8'hbc)}))) ?
                  reg2583[(5'h11):(4'h9)] : (7'h40));
              reg2706 <= (7'h4e);
            end
          else
            begin
              reg2702 <= reg2542[(5'h12):(1'h0)];
              reg2703 = reg2641[(2'h2):(2'h2)];
              reg2705 = reg2654;
              reg2706 <= (7'h50);
              reg2707 <= {(wire2475 && (~|($signed((8'h9f)) | (reg2510 == reg2608))))};
              reg2708 = (reg2613[(1'h1):(1'h0)] ?
                  (8'ha8) : ((((reg2478 >> reg2655) <= (~reg2671)) ?
                      ($signed(reg2615) >> {reg2561}) : reg2604[(4'ha):(2'h2)]) == (~^({reg2591} < $unsigned((7'h53))))));
            end
        end
      else
        begin
          reg2699 = ($signed((!reg2599)) || reg2547[(3'h5):(1'h0)]);
        end
      if (reg2704[(5'h18):(5'h11)])
        begin
          if (({($signed($signed((8'had))) ?
                      ((reg2487 >>> (8'hb3)) ?
                          wire2473[(1'h0):(1'h0)] : $unsigned(reg2541)) : (7'h40)),
                  $unsigned((^(|reg2693))),
                  reg2674[(4'he):(4'hb)]} ?
              reg2701[(3'h7):(3'h4)] : ((~^reg2513[(5'h15):(5'h10)]) >= (reg2517[(4'ha):(4'ha)] - $unsigned(reg2591)))))
            begin
              reg2709 <= reg2676;
              reg2710 <= wire2474;
              reg2711 = $unsigned(reg2678[(3'h7):(2'h3)]);
              reg2712 = {reg2615[(3'h4):(2'h3)],
                  $signed((reg2557[(4'hd):(4'hc)] <<< $unsigned((^~reg2670))))};
              reg2713 = (&$unsigned(reg2515[(3'h4):(3'h4)]));
            end
          else
            begin
              reg2709 <= reg2707;
              reg2711 = ((($unsigned({wire2695}) ?
                  (8'ha2) : (8'ha6)) ~^ {$signed($unsigned(reg2599)),
                  ((-reg2537) && (-wire2696)),
                  (~&$unsigned((8'ha9)))}) ^ (7'h4d));
              reg2714 <= (reg2513 ? (8'ha1) : $unsigned(reg2543));
              reg2715 = ({$signed(reg2685[(4'h9):(4'h9)]),
                      $unsigned($unsigned(reg2630))} ?
                  reg2707[(2'h2):(2'h2)] : reg2562);
              reg2716 <= {($unsigned($unsigned((reg2526 != reg2702))) ?
                      $unsigned(reg2547[(3'h7):(1'h0)]) : (&((~&reg2611) <<< reg2495[(2'h3):(2'h3)]))),
                  reg2709[(4'hd):(4'h8)],
                  reg2615[(1'h1):(1'h1)]};
            end
          reg2717 <= $signed($signed(($signed(reg2567[(1'h0):(1'h0)]) != reg2611[(4'hd):(4'hc)])));
          if (reg2713[(4'hb):(4'ha)])
            begin
              reg2718 <= (-$unsigned((|reg2671[(4'hd):(3'h4)])));
              reg2719 = (wire2663 ?
                  (8'ha5) : {wire2663,
                      ((~&$unsigned(reg2544)) ?
                          ($signed((7'h4f)) ?
                              reg2488 : (reg2525 ?
                                  reg2641 : wire2470)) : {((8'hab) & (8'hb5)),
                              {(8'hba), reg2555},
                              $signed((7'h55))}),
                      (^~($unsigned(reg2579) != {reg2597, (8'haf), reg2593}))});
              reg2720 = reg2487;
              reg2721 <= (~^(~((~(reg2709 == reg2704)) < ($signed((7'h4c)) && reg2707))));
            end
          else
            begin
              reg2719 = reg2564[(5'h12):(1'h1)];
              reg2721 <= $unsigned($unsigned(reg2501[(1'h1):(1'h0)]));
              reg2722 <= reg2604[(5'h10):(3'h5)];
              reg2723 <= reg2679[(4'hc):(3'h4)];
              reg2724 <= $unsigned((|reg2676[(3'h4):(1'h1)]));
            end
          for (forvar2725 = (1'h0); (forvar2725 < (1'h0)); forvar2725 = (forvar2725 + (1'h1)))
            begin
              reg2726 <= wire2474;
              reg2727 <= (^({($unsigned(reg2617) ?
                      $unsigned(reg2702) : (reg2571 + reg2649)),
                  $unsigned((reg2551 <<< reg2711))} >>> (reg2561[(1'h0):(1'h0)] ?
                  {reg2580[(4'hb):(4'hb)]} : reg2671)));
              reg2728 = (8'ha7);
              reg2729 <= ((~^($unsigned($unsigned(reg2634)) - reg2656[(1'h1):(1'h1)])) ?
                  ((reg2551 ?
                          ({wire2696,
                              reg2638} * reg2525) : ((~reg2513) >>> (+forvar2725))) ?
                      (reg2580 >> (-{reg2487})) : reg2656[(2'h2):(1'h0)]) : reg2574);
              reg2730 <= ({($unsigned((reg2510 <= (7'h48))) && $unsigned($signed((7'h52)))),
                      reg2565[(2'h3):(2'h2)],
                      (8'ha0)} ?
                  ($signed(wire2640) == $signed(reg2704[(5'h11):(4'ha)])) : wire2696[(4'ha):(3'h4)]);
            end
          if ((reg2709 - reg2630))
            begin
              reg2731 <= (7'h53);
              reg2732 = $signed($unsigned(reg2709));
              reg2733 <= (($unsigned($signed((reg2656 << (8'ha5)))) ^~ $signed((8'h9c))) >>> reg2614[(5'h1b):(4'h9)]);
              reg2734 = reg2710;
            end
          else
            begin
              reg2732 = $signed((reg2726 & (reg2597 >= (wire2473[(4'ha):(4'ha)] ?
                  $signed(reg2646) : reg2579[(5'h15):(5'h10)]))));
              reg2733 <= (-(-(8'ha0)));
              reg2735 <= (reg2671 ?
                  reg2537[(1'h0):(1'h0)] : ($signed(reg2520) ?
                      reg2726 : (|reg2497[(5'h14):(5'h12)])));
            end
          reg2736 = reg2515;
          reg2737 <= reg2493[(4'hd):(2'h2)];
        end
      else
        begin
          if ($signed($unsigned(($signed(wire2470) ? reg2684 : reg2555))))
            begin
              reg2711 = $signed($signed($unsigned((7'h54))));
              reg2714 <= {(~^($unsigned($signed(reg2526)) << ($signed(reg2531) ?
                      $unsigned(reg2545) : (+reg2684))))};
              reg2715 = $signed($signed((-(~^(7'h57)))));
              reg2719 = (^~((7'h51) != reg2641[(3'h4):(2'h3)]));
              reg2721 <= (reg2480 ?
                  reg2660 : ($unsigned($signed(reg2599[(2'h3):(2'h3)])) ?
                      ({reg2674, reg2736[(5'h11):(4'h9)]} ?
                          reg2541[(4'he):(3'h5)] : (-$signed(reg2515))) : {(^reg2698),
                          $unsigned(reg2586[(4'he):(4'he)]),
                          $signed(wire2471)}));
              reg2722 <= reg2703;
            end
          else
            begin
              reg2711 = reg2678;
              reg2714 <= ((($signed($unsigned(reg2486)) <<< $unsigned(reg2520[(5'h16):(4'hf)])) ?
                  (-({reg2545, reg2497, reg2679} ~^ (reg2602 ?
                      reg2654 : reg2649))) : (reg2659 <<< ((reg2734 ?
                      reg2713 : wire2662) << $unsigned(reg2567)))) & reg2671);
              reg2716 <= (reg2615[(1'h1):(1'h0)] >= {{$signed($signed(reg2478))}});
              reg2719 = reg2520[(4'hc):(4'h9)];
              reg2721 <= reg2649[(1'h0):(1'h0)];
              reg2722 <= ((|((~|(reg2528 ? reg2676 : reg2716)) ?
                      (~&(reg2588 ? (8'ha0) : reg2708)) : reg2638)) ?
                  (~|(reg2721[(5'h10):(4'h9)] ?
                      $unsigned((reg2547 <<< reg2604)) : $signed($signed(reg2703)))) : $unsigned(reg2486[(4'hd):(2'h3)]));
            end
          reg2725 = (^reg2555[(2'h3):(1'h1)]);
          if (reg2705)
            begin
              reg2726 <= ($signed((8'hb9)) ?
                  $unsigned(reg2567) : reg2569[(5'h11):(4'h8)]);
              reg2727 <= reg2562;
              reg2729 <= reg2734;
              reg2732 = reg2714;
              reg2733 <= ($signed($unsigned(($signed(reg2541) << (~reg2480)))) <<< (+(reg2497[(5'h16):(5'h15)] ?
                  (7'h46) : ((reg2614 ? (7'h42) : reg2597) ?
                      {reg2507, reg2737, reg2702} : $signed(reg2728)))));
              reg2735 <= ((~^($signed($signed(reg2721)) ?
                  $signed(reg2716) : $unsigned((!reg2693)))) << ($signed($unsigned(reg2729[(1'h0):(1'h0)])) ?
                  $signed((reg2602[(3'h5):(2'h3)] >>> (reg2574 >= reg2707))) : reg2705[(4'h8):(2'h2)]));
              reg2736 = reg2504[(5'h11):(4'he)];
            end
          else
            begin
              reg2728 = $signed(((^~((reg2617 ^~ reg2697) * (&wire2640))) + ((-reg2671[(5'h14):(5'h12)]) ^~ (reg2638[(5'h13):(1'h1)] | (+reg2709)))));
              reg2729 <= reg2542;
              reg2730 <= reg2556[(3'h7):(3'h6)];
              reg2731 <= $signed(((-(reg2720[(3'h4):(1'h0)] ?
                  $unsigned(reg2625) : reg2723)) * {((reg2675 ?
                      reg2678 : reg2544) <<< (~&reg2520)),
                  (7'h49)}));
              reg2733 <= ((($unsigned((^~reg2717)) * ($signed(reg2701) ^~ $signed(reg2510))) >>> reg2678[(2'h3):(2'h2)]) ?
                  $signed(((+(reg2561 ?
                      wire2695 : reg2597)) ~^ wire2474[(4'h8):(1'h1)])) : reg2729[(1'h0):(1'h0)]);
              reg2734 = (~reg2706[(5'h13):(5'h13)]);
              reg2735 <= reg2553[(3'h6):(2'h2)];
            end
          for (forvar2737 = (1'h0); (forvar2737 < (1'h0)); forvar2737 = (forvar2737 + (1'h1)))
            begin
              reg2738 <= reg2719[(3'h5):(1'h1)];
              reg2739 = ($signed({$signed(((8'ha9) < reg2737))}) ?
                  (&{((|reg2726) << {reg2723,
                          reg2562,
                          (7'h53)})}) : ((((8'hb0) ?
                      reg2564 : reg2578) ^ {(&reg2707),
                      (|reg2660)}) ^ $unsigned($unsigned($signed(wire2473)))));
            end
          for (forvar2740 = (1'h0); (forvar2740 < (3'h5)); forvar2740 = (forvar2740 + (1'h1)))
            begin
              reg2741 = (((7'h42) ~^ reg2597) ?
                  ((((~^wire2471) ?
                      (^~reg2713) : (reg2727 ?
                          reg2553 : reg2487)) == {(reg2521 ? reg2728 : (7'h54)),
                      $signed((8'h9d))}) * $unsigned(((^reg2547) != $signed(wire2696)))) : (($signed((reg2693 ?
                          wire2469 : reg2697)) < (reg2537[(1'h1):(1'h0)] == reg2573[(2'h3):(1'h1)])) ?
                      ((reg2671 ~^ ((8'h9e) ?
                          (8'hbf) : reg2654)) != reg2635[(1'h1):(1'h1)]) : {{{(8'hb2),
                                  reg2515,
                                  (8'hbd)},
                              $unsigned(reg2720),
                              reg2731},
                          $signed((reg2520 ^~ reg2531)),
                          (^{reg2583})}));
              reg2742 <= $unsigned($signed(reg2597[(4'he):(4'h9)]));
              reg2743 <= ((~&(reg2679 ? reg2486 : {reg2716})) ?
                  ((|$unsigned((reg2577 ?
                      reg2697 : reg2521))) & (reg2651[(1'h1):(1'h1)] ~^ {(!reg2712)})) : reg2559);
              reg2744 <= $unsigned((~((~^wire2695[(3'h7):(2'h2)]) ?
                  (&(reg2734 ?
                      reg2674 : reg2617)) : $unsigned(reg2564[(5'h12):(5'h11)]))));
              reg2745 = $signed({$unsigned(reg2493[(5'h19):(3'h6)]),
                  ((reg2538 ? {(8'hbc)} : reg2523) ?
                      reg2720[(3'h6):(3'h6)] : $unsigned($signed(reg2732))),
                  ($signed(reg2743[(4'h8):(2'h2)]) <<< (reg2676 << $unsigned(reg2488)))});
              reg2746 <= {(|({{reg2688, reg2638},
                      reg2528[(1'h0):(1'h0)]} * (7'h4f)))};
              reg2747 <= (reg2510 ?
                  reg2709[(4'h8):(1'h0)] : $signed(($signed((reg2708 ?
                      forvar2725 : reg2564)) <<< ($unsigned(reg2706) > reg2531))));
            end
        end
      if ({(({(reg2614 ?
                  reg2562 : reg2641)} > reg2732[(2'h2):(2'h2)]) == reg2634),
          (^~$signed(($signed(reg2493) & $signed(reg2515))))})
        begin
          reg2748 <= ((-reg2646[(4'ha):(4'h9)]) == (reg2671[(2'h2):(2'h2)] ~^ $unsigned(($unsigned((8'hbc)) ?
              reg2577 : ((7'h46) ? reg2590 : reg2716)))));
          reg2749 = reg2526;
        end
      else
        begin
          for (forvar2748 = (1'h0); (forvar2748 < (3'h5)); forvar2748 = (forvar2748 + (1'h1)))
            begin
              reg2750 <= (8'hab);
              reg2751 <= reg2747;
            end
        end
    end
  always
    @(posedge clk) begin
      reg2752 = $unsigned((reg2580[(4'h8):(2'h2)] ~^ (^(wire2469[(2'h2):(1'h1)] ?
          $signed(reg2488) : (reg2544 ? (7'h4d) : (8'hb2))))));
      reg2753 = ((reg2604[(3'h6):(3'h4)] - $unsigned($unsigned((reg2543 != wire2475)))) ?
          reg2538[(4'he):(4'hc)] : reg2731[(3'h7):(1'h1)]);
      for (forvar2754 = (1'h0); (forvar2754 < (3'h4)); forvar2754 = (forvar2754 + (1'h1)))
        begin
          if ($signed((reg2579 - $signed((^wire2662)))))
            begin
              reg2755 = {(~^((~|(reg2531 ^ (8'ha4))) && reg2593[(2'h2):(2'h2)])),
                  $signed(reg2690[(3'h6):(2'h2)])};
              reg2756 = (8'h9e);
              reg2757 <= $unsigned(($unsigned({(^~wire2473),
                  ((8'hbd) <= reg2627),
                  (-reg2590)}) ~^ (reg2706[(3'h6):(1'h0)] ?
                  (!$signed(reg2646)) : $signed($signed((8'hbd))))));
              reg2758 = $signed($unsigned((|(-(reg2487 == reg2675)))));
              reg2759 = ($unsigned(reg2582) ?
                  ($signed(((-reg2574) ?
                      (reg2735 ? reg2510 : reg2586) : {reg2559,
                          reg2614,
                          reg2545})) ^~ (-reg2758)) : (reg2690 ^ {$unsigned((reg2710 ?
                          reg2735 : reg2671)),
                      $unsigned(((7'h4c) == reg2635))}));
              reg2760 = (reg2738[(4'he):(1'h1)] ?
                  ($unsigned($unsigned($signed(wire2471))) ?
                      $unsigned({{reg2685},
                          $unsigned(reg2746),
                          (^~(8'hb5))}) : ({(~reg2729),
                              (reg2528 ? (8'hae) : reg2517)} ?
                          reg2538 : reg2748)) : $signed((8'haa)));
            end
          else
            begin
              reg2757 <= $unsigned($signed($signed(((!reg2480) ^ (8'hae)))));
              reg2758 = reg2583;
              reg2759 = reg2641;
              reg2761 <= {($signed(reg2602[(3'h4):(1'h0)]) ~^ $unsigned((reg2634[(2'h2):(1'h1)] ~^ $unsigned((8'ha5))))),
                  reg2571};
              reg2762 <= $signed(reg2675[(1'h1):(1'h0)]);
            end
          if (((^(~|((~^reg2685) ~^ (!(7'h47))))) <= ((reg2710 < $unsigned(reg2651[(3'h4):(1'h0)])) ?
              wire2470 : ($signed((8'hab)) ?
                  $unsigned(reg2751[(2'h2):(1'h1)]) : ((wire2468 ?
                      reg2723 : reg2760) == reg2561[(3'h6):(3'h6)])))))
            begin
              reg2763 <= {reg2721,
                  (+({((7'h56) == reg2685)} ?
                      ($signed(reg2743) <= $unsigned(reg2761)) : {reg2659,
                          (reg2760 ^ wire2475)})),
                  ((&(~|(~^reg2523))) ~^ (&$signed($signed(reg2702))))};
              reg2764 <= (!({$unsigned(reg2487[(1'h1):(1'h0)])} ?
                  $signed(reg2547[(3'h6):(3'h5)]) : $unsigned($unsigned(reg2493))));
              reg2765 <= reg2526[(4'h8):(3'h4)];
              reg2766 = (|($signed(((~wire2694) >= (^reg2487))) ?
                  (($unsigned((7'h55)) ?
                      (reg2605 ? reg2765 : reg2654) : (reg2564 ?
                          wire2471 : reg2733)) ^~ reg2526) : reg2591));
              reg2767 = ((^~{(8'hb4),
                  reg2495[(1'h0):(1'h0)]}) + ($unsigned($unsigned($unsigned(wire2472))) | $signed({(reg2718 * reg2531),
                  ((7'h57) ^~ reg2605),
                  $signed(reg2583)})));
              reg2768 <= $signed(reg2521[(3'h7):(3'h5)]);
              reg2769 = reg2731;
            end
          else
            begin
              reg2766 = (8'ha2);
              reg2768 <= (reg2484[(5'h13):(5'h13)] ?
                  $unsigned({$unsigned((reg2675 ? (8'hb3) : reg2726)),
                      $unsigned($unsigned((7'h55)))}) : (reg2727[(1'h1):(1'h0)] ^~ reg2651[(3'h4):(2'h3)]));
              reg2770 <= $unsigned({reg2582[(1'h1):(1'h0)],
                  (&reg2484),
                  reg2515[(4'hb):(4'h8)]});
              reg2771 = $unsigned(((reg2588 >>> $signed(reg2561[(3'h7):(2'h3)])) ?
                  {((wire2694 ? reg2656 : reg2638) < reg2578),
                      ($unsigned(wire2470) ? reg2690[(2'h3):(1'h0)] : reg2688),
                      reg2693[(1'h0):(1'h0)]} : ((reg2625 ?
                      (reg2731 ?
                          reg2497 : wire2662) : reg2556[(5'h11):(4'hc)]) ^ $unsigned($unsigned(reg2727)))));
              reg2772 <= ({reg2646,
                  (~&($signed(reg2700) ?
                      $unsigned(reg2727) : {reg2753,
                          reg2561,
                          reg2674}))} ^ $unsigned(reg2660[(5'h11):(3'h7)]));
              reg2773 = $unsigned($unsigned({$unsigned(reg2567)}));
            end
          reg2774 = ((^~{reg2487[(1'h1):(1'h0)]}) << reg2656[(1'h1):(1'h1)]);
          if ((reg2488 ?
              (reg2574[(4'he):(4'h8)] >> (+$unsigned($signed((7'h4f))))) : (!{(~^$signed(forvar2754)),
                  $signed(reg2759)})))
            begin
              reg2775 <= (^$unsigned(reg2771));
            end
          else
            begin
              reg2775 <= {((reg2765 ?
                      {reg2750[(1'h1):(1'h0)],
                          ((7'h4b) ? reg2744 : reg2594),
                          (reg2731 < reg2646)} : $signed((&reg2488))) << (reg2537[(2'h2):(1'h1)] ?
                      reg2605 : (!$unsigned(reg2710))))};
              reg2776 <= $signed($signed((7'h57)));
              reg2777 = (7'h48);
            end
          reg2778 <= {$signed((reg2569[(5'h1a):(2'h2)] >>> {(reg2726 ^~ reg2762),
                  reg2760[(1'h0):(1'h0)]})),
              (~|reg2510[(4'hb):(2'h2)]),
              (reg2567[(5'h13):(1'h1)] >>> $signed((~&(wire2468 ?
                  (8'ha5) : reg2716))))};
          reg2779 <= $unsigned($signed((~|$unsigned(reg2675))));
        end
      reg2780 = {(reg2685 ?
              ((~^$signed(reg2641)) ^~ (~$signed(reg2701))) : ((reg2777 ?
                  wire2469[(2'h2):(2'h2)] : wire2664) <<< (~|$signed(reg2543)))),
          ($unsigned(((reg2582 && reg2704) ?
              $signed(reg2484) : (reg2638 * wire2473))) >>> (!$signed((7'h48)))),
          ((!(~&reg2733[(4'hc):(3'h6)])) - reg2742[(3'h6):(1'h0)])};
      reg2781 <= ($signed(((reg2767 ? $unsigned((7'h43)) : $signed(reg2775)) ?
          ((wire2473 <<< reg2706) ?
              $unsigned(reg2704) : ((8'h9f) ?
                  reg2493 : reg2478)) : (reg2773[(2'h2):(1'h1)] ?
              reg2545 : reg2678))) >>> reg2761);
      if ((wire2469[(3'h5):(2'h2)] ?
          reg2774 : $signed($unsigned((reg2721 >>> (reg2690 <= reg2493))))))
        begin
          reg2782 = (~&(reg2714[(4'h9):(2'h2)] ~^ reg2649));
          reg2783 <= ($unsigned(reg2660) > $signed((^~$unsigned(wire2468))));
          for (forvar2784 = (1'h0); (forvar2784 < (3'h6)); forvar2784 = (forvar2784 + (1'h1)))
            begin
              reg2785 = ((8'ha9) == (~reg2735[(3'h6):(2'h2)]));
              reg2786 <= reg2558;
              reg2787 <= (($unsigned(reg2599[(2'h3):(2'h3)]) ?
                      ({((8'h9f) ^ reg2525)} ?
                          $unsigned((reg2779 ?
                              forvar2754 : reg2557)) : (~reg2779)) : reg2486[(2'h2):(2'h2)]) ?
                  ($signed(reg2591[(5'h15):(4'ha)]) ?
                      $unsigned($unsigned(reg2714)) : $unsigned((~^reg2495[(2'h2):(2'h2)]))) : ((+$signed({(8'hbb)})) >>> (~$signed({reg2688,
                      reg2493}))));
              reg2788 = (~&$signed(($signed(reg2762[(3'h5):(1'h0)]) ?
                  wire2640 : (~&reg2611))));
              reg2789 <= {$unsigned($unsigned(((&reg2762) + {reg2764}))),
                  reg2783,
                  reg2701};
            end
        end
      else
        begin
          for (forvar2782 = (1'h0); (forvar2782 < (1'h0)); forvar2782 = (forvar2782 + (1'h1)))
            begin
              reg2783 <= ($signed((&reg2561)) || (($signed($unsigned(reg2690)) ?
                      (7'h47) : reg2733) ?
                  $signed((7'h55)) : reg2501[(1'h0):(1'h0)]));
              reg2784 = (|(~^(reg2504 ~^ {(reg2646 ? reg2564 : reg2679),
                  reg2746,
                  $unsigned(wire2663)})));
              reg2785 = reg2638[(5'h13):(5'h11)];
              reg2786 <= $unsigned((~((|$unsigned(reg2675)) ~^ $signed(wire2473))));
            end
          if (reg2547[(3'h5):(2'h3)])
            begin
              reg2788 = {$unsigned($unsigned($unsigned((reg2787 << reg2674)))),
                  (~^(|$signed(reg2569)))};
              reg2789 <= ($signed(((7'h51) ~^ reg2504)) ?
                  $unsigned(($signed(reg2613) >> (^~(reg2539 ?
                      reg2558 : reg2582)))) : (7'h56));
              reg2790 <= {(^~(reg2766[(4'hf):(4'hf)] ?
                      reg2478[(2'h3):(2'h2)] : reg2567)),
                  $unsigned(reg2761),
                  reg2520};
              reg2791 = ($unsigned(reg2761[(5'h10):(5'h10)]) ?
                  (~$unsigned($unsigned((reg2764 ?
                      reg2772 : reg2484)))) : $signed($unsigned($unsigned(reg2783))));
              reg2792 <= $unsigned(($signed($unsigned({reg2763,
                      (8'ha1),
                      (8'hbf)})) ?
                  {{(reg2577 >> (8'hb0))},
                      $unsigned($unsigned(reg2722))} : ($unsigned({reg2733,
                      reg2578}) ~^ $signed((-reg2515)))));
              reg2793 = reg2507[(2'h2):(2'h2)];
            end
          else
            begin
              reg2788 = ($signed(((reg2596[(3'h7):(3'h6)] ?
                          (!reg2630) : $signed(reg2768)) ?
                      (reg2668[(5'h14):(4'he)] ?
                          (reg2753 >> reg2594) : (-reg2569)) : ($unsigned((7'h47)) ?
                          (reg2668 - reg2625) : (&reg2768)))) ?
                  (wire2663 || reg2763) : {((8'hb4) ?
                          reg2730[(5'h11):(4'he)] : reg2582[(2'h3):(1'h0)]),
                      reg2789,
                      $signed(reg2758)});
            end
          for (forvar2794 = (1'h0); (forvar2794 < (1'h1)); forvar2794 = (forvar2794 + (1'h1)))
            begin
              reg2795 <= {forvar2782[(4'hd):(4'hc)]};
              reg2796 <= ({reg2510} ?
                  ($signed(reg2795) ?
                      reg2738[(5'h10):(4'hd)] : (&(((8'hba) ~^ (7'h42)) < $unsigned(reg2615)))) : (&((-(|reg2721)) ?
                      ($signed(forvar2782) ?
                          $unsigned(reg2507) : reg2604) : ((+reg2762) ?
                          reg2501 : wire2696))));
              reg2797 <= (!(reg2591 >> (^~((&reg2602) ?
                  (wire2468 ? reg2760 : reg2668) : $unsigned(reg2608)))));
              reg2798 = (reg2515 ?
                  {((~$unsigned(reg2761)) ?
                          $signed($unsigned(reg2613)) : (reg2752[(1'h0):(1'h0)] << reg2674)),
                      $signed($signed((reg2771 ? reg2602 : reg2493))),
                      $signed(reg2627[(2'h2):(1'h0)])} : {{({reg2521,
                                  reg2714,
                                  reg2785} ?
                              $unsigned(reg2596) : wire2640[(5'h16):(3'h4)]),
                          ((reg2722 ? reg2556 : reg2625) ^ (8'h9d))}});
              reg2799 <= reg2544[(2'h3):(1'h1)];
              reg2800 = (^~{(~|(^~wire2696)),
                  reg2504,
                  $unsigned(((&wire2471) ?
                      reg2670[(4'ha):(3'h4)] : {reg2768, reg2759}))});
              reg2801 <= $signed($signed(((((8'hac) << reg2515) ?
                      (reg2608 << reg2729) : {reg2602}) ?
                  $signed((wire2664 ?
                      (7'h53) : reg2634)) : reg2701[(4'hd):(4'hd)])));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1773  (y, clk, wire1778, wire1777, wire1776, wire1775, wire1774);
  output wire [(32'h1c53):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire1778;
  input wire signed [(5'h17):(1'h0)] wire1777;
  input wire signed [(4'h8):(1'h0)] wire1776;
  input wire signed [(5'h1e):(1'h0)] wire1775;
  input wire signed [(5'h10):(1'h0)] wire1774;
  wire [(5'h19):(1'h0)] wire2165;
  wire signed [(5'h16):(1'h0)] wire2078;
  wire signed [(4'hc):(1'h0)] wire2077;
  wire signed [(5'h17):(1'h0)] wire2059;
  wire signed [(5'h16):(1'h0)] wire2015;
  wire signed [(5'h12):(1'h0)] wire2007;
  wire signed [(4'he):(1'h0)] wire2006;
  wire signed [(5'h11):(1'h0)] wire1909;
  wire [(5'h16):(1'h0)] wire1907;
  wire signed [(4'hb):(1'h0)] wire1906;
  wire signed [(4'hd):(1'h0)] wire1905;
  wire [(5'h10):(1'h0)] wire1904;
  wire signed [(4'hf):(1'h0)] wire1810;
  reg [(5'h1e):(1'h0)] reg2194 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2193 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2192 = (1'h0);
  reg [(5'h16):(1'h0)] reg2189 = (1'h0);
  reg [(5'h18):(1'h0)] reg2187 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2183 = (1'h0);
  reg [(5'h19):(1'h0)] reg2182 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2180 = (1'h0);
  reg [(5'h11):(1'h0)] reg2179 = (1'h0);
  reg [(5'h13):(1'h0)] reg2177 = (1'h0);
  reg [(4'h8):(1'h0)] reg2175 = (1'h0);
  reg [(5'h19):(1'h0)] reg2174 = (1'h0);
  reg [(4'h8):(1'h0)] reg2173 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2172 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2168 = (1'h0);
  reg [(4'hc):(1'h0)] reg2167 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2164 = (1'h0);
  reg [(3'h5):(1'h0)] reg2163 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2162 = (1'h0);
  reg [(5'h15):(1'h0)] reg2158 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2156 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2155 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2151 = (1'h0);
  reg [(5'h12):(1'h0)] reg2147 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2146 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2143 = (1'h0);
  reg [(3'h6):(1'h0)] reg2141 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2139 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2137 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2135 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2132 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2130 = (1'h0);
  reg [(5'h11):(1'h0)] reg2127 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2121 = (1'h0);
  reg [(2'h3):(1'h0)] reg2120 = (1'h0);
  reg [(4'ha):(1'h0)] reg2119 = (1'h0);
  reg [(4'hd):(1'h0)] reg2114 = (1'h0);
  reg [(5'h19):(1'h0)] reg2113 = (1'h0);
  reg [(5'h17):(1'h0)] reg2111 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2110 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2108 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2107 = (1'h0);
  reg [(5'h15):(1'h0)] reg2103 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2102 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2100 = (1'h0);
  reg [(5'h11):(1'h0)] reg2097 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2096 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2089 = (1'h0);
  reg [(5'h13):(1'h0)] reg2088 = (1'h0);
  reg [(3'h5):(1'h0)] reg2085 = (1'h0);
  reg [(5'h10):(1'h0)] reg2083 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2082 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2081 = (1'h0);
  reg [(5'h13):(1'h0)] reg2073 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2069 = (1'h0);
  reg [(5'h13):(1'h0)] reg2063 = (1'h0);
  reg [(3'h6):(1'h0)] reg2062 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2058 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2057 = (1'h0);
  reg [(5'h19):(1'h0)] reg2052 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2049 = (1'h0);
  reg [(5'h16):(1'h0)] reg2047 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2044 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2043 = (1'h0);
  reg [(2'h3):(1'h0)] reg2040 = (1'h0);
  reg [(4'hc):(1'h0)] reg2038 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2034 = (1'h0);
  reg [(2'h2):(1'h0)] reg2031 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2030 = (1'h0);
  reg [(4'he):(1'h0)] reg2028 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2022 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2021 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2020 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2019 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2012 = (1'h0);
  reg [(4'hd):(1'h0)] reg2011 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2010 = (1'h0);
  reg [(5'h10):(1'h0)] reg2009 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2004 = (1'h0);
  reg [(4'hf):(1'h0)] reg1997 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2001 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2000 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1993 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1992 = (1'h0);
  reg [(5'h17):(1'h0)] reg1990 = (1'h0);
  reg [(5'h14):(1'h0)] reg1989 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1988 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1987 = (1'h0);
  reg [(4'h8):(1'h0)] reg1985 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1984 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1980 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1978 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1977 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1975 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1972 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1971 = (1'h0);
  reg [(4'he):(1'h0)] reg1970 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1969 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1968 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1966 = (1'h0);
  reg [(5'h10):(1'h0)] reg1965 = (1'h0);
  reg [(3'h5):(1'h0)] reg1961 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1960 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1959 = (1'h0);
  reg [(5'h16):(1'h0)] reg1958 = (1'h0);
  reg [(3'h7):(1'h0)] reg1957 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1955 = (1'h0);
  reg [(5'h13):(1'h0)] reg1953 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1952 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1951 = (1'h0);
  reg [(4'hd):(1'h0)] reg1949 = (1'h0);
  reg [(4'h8):(1'h0)] reg1948 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1947 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1946 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1945 = (1'h0);
  reg [(3'h7):(1'h0)] reg1944 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1942 = (1'h0);
  reg [(5'h12):(1'h0)] reg1941 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1937 = (1'h0);
  reg [(5'h11):(1'h0)] reg1933 = (1'h0);
  reg [(5'h13):(1'h0)] reg1932 = (1'h0);
  reg [(5'h16):(1'h0)] reg1931 = (1'h0);
  reg [(3'h5):(1'h0)] reg1930 = (1'h0);
  reg [(5'h12):(1'h0)] reg1927 = (1'h0);
  reg [(4'h9):(1'h0)] reg1926 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1920 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1917 = (1'h0);
  reg [(5'h12):(1'h0)] reg1916 = (1'h0);
  reg [(5'h18):(1'h0)] reg1914 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1911 = (1'h0);
  reg [(5'h11):(1'h0)] reg1908 = (1'h0);
  reg [(5'h19):(1'h0)] reg1902 = (1'h0);
  reg [(3'h4):(1'h0)] reg1901 = (1'h0);
  reg [(3'h7):(1'h0)] reg1900 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1896 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1895 = (1'h0);
  reg [(5'h10):(1'h0)] reg1894 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1891 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1890 = (1'h0);
  reg [(4'hb):(1'h0)] reg1872 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1889 = (1'h0);
  reg [(5'h17):(1'h0)] reg1885 = (1'h0);
  reg [(2'h3):(1'h0)] reg1884 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1883 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1880 = (1'h0);
  reg [(5'h18):(1'h0)] reg1879 = (1'h0);
  reg [(3'h5):(1'h0)] reg1878 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1877 = (1'h0);
  reg [(5'h12):(1'h0)] reg1876 = (1'h0);
  reg [(4'hf):(1'h0)] reg1874 = (1'h0);
  reg [(4'h9):(1'h0)] reg1873 = (1'h0);
  reg [(5'h17):(1'h0)] reg1870 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1865 = (1'h0);
  reg [(5'h13):(1'h0)] reg1864 = (1'h0);
  reg [(5'h19):(1'h0)] reg1863 = (1'h0);
  reg [(4'he):(1'h0)] reg1859 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1858 = (1'h0);
  reg [(4'hc):(1'h0)] reg1857 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1855 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1854 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1851 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1849 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1811 = (1'h0);
  reg [(5'h11):(1'h0)] reg1840 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1838 = (1'h0);
  reg [(4'hc):(1'h0)] reg1836 = (1'h0);
  reg [(3'h6):(1'h0)] reg1832 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1831 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1824 = (1'h0);
  reg [(4'ha):(1'h0)] reg1822 = (1'h0);
  reg [(5'h18):(1'h0)] reg1821 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1820 = (1'h0);
  reg [(4'hf):(1'h0)] reg1819 = (1'h0);
  reg [(2'h3):(1'h0)] reg1818 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1816 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1814 = (1'h0);
  reg [(4'he):(1'h0)] reg1813 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1807 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1803 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1801 = (1'h0);
  reg [(5'h16):(1'h0)] reg1800 = (1'h0);
  reg [(5'h18):(1'h0)] reg1799 = (1'h0);
  reg [(3'h4):(1'h0)] reg1798 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1797 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1793 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1791 = (1'h0);
  reg [(4'h9):(1'h0)] reg1788 = (1'h0);
  reg [(5'h11):(1'h0)] reg1787 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1786 = (1'h0);
  reg [(4'ha):(1'h0)] reg1785 = (1'h0);
  reg [(4'hc):(1'h0)] reg1783 = (1'h0);
  reg [(5'h16):(1'h0)] reg1782 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2191 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2190 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2188 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2186 = (1'h0);
  reg [(4'he):(1'h0)] reg2185 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2184 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2181 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2178 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2176 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2171 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2170 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2169 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2166 = (1'h0);
  reg [(4'hc):(1'h0)] reg2161 = (1'h0);
  reg [(4'hb):(1'h0)] reg2160 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2159 = (1'h0);
  reg [(3'h7):(1'h0)] reg2157 = (1'h0);
  reg [(5'h19):(1'h0)] reg2154 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2153 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2152 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2150 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2149 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2148 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2145 = (1'h0);
  reg [(4'hb):(1'h0)] reg2144 = (1'h0);
  reg [(3'h7):(1'h0)] reg2142 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2140 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2138 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2136 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2134 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2133 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2131 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2129 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2128 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2126 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2125 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar2124 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2123 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2122 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2118 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2117 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2116 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2115 = (1'h0);
  reg [(5'h18):(1'h0)] reg2104 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2112 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2109 = (1'h0);
  reg [(4'h9):(1'h0)] reg2106 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2105 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar2104 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2101 = (1'h0);
  reg [(5'h18):(1'h0)] reg2099 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2098 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2095 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2094 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2093 = (1'h0);
  reg [(4'hc):(1'h0)] reg2092 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2091 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2090 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2087 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2086 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2084 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2080 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2079 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2076 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2075 = (1'h0);
  reg [(5'h18):(1'h0)] reg2074 = (1'h0);
  reg [(5'h15):(1'h0)] reg2072 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2071 = (1'h0);
  reg [(4'hd):(1'h0)] reg2070 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2068 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2067 = (1'h0);
  reg [(4'hb):(1'h0)] reg2066 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2065 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2064 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2061 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2060 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2056 = (1'h0);
  reg [(3'h4):(1'h0)] reg2055 = (1'h0);
  reg [(5'h15):(1'h0)] reg2054 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2053 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2051 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2050 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2048 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2046 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2045 = (1'h0);
  reg [(5'h12):(1'h0)] reg2042 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2041 = (1'h0);
  reg [(4'h9):(1'h0)] reg2039 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2037 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2036 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2035 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2033 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2032 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2029 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2027 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2026 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2025 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2024 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2023 = (1'h0);
  reg [(5'h15):(1'h0)] reg2018 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar2017 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2016 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2014 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2013 = (1'h0);
  reg [(5'h13):(1'h0)] reg2008 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2005 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2003 = (1'h0);
  reg [(3'h6):(1'h0)] reg2002 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1999 = (1'h0);
  reg [(3'h5):(1'h0)] reg1998 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1997 = (1'h0);
  reg [(5'h19):(1'h0)] reg1996 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1995 = (1'h0);
  reg [(4'he):(1'h0)] reg1994 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1991 = (1'h0);
  reg [(5'h18):(1'h0)] reg1986 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1983 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1982 = (1'h0);
  reg [(5'h15):(1'h0)] reg1981 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1979 = (1'h0);
  reg [(5'h14):(1'h0)] reg1976 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1974 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1973 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1967 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1964 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1938 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1963 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1962 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1956 = (1'h0);
  reg [(5'h17):(1'h0)] reg1954 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1950 = (1'h0);
  reg [(4'ha):(1'h0)] reg1943 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1940 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1939 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1938 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1936 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1935 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1934 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1929 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1928 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1925 = (1'h0);
  reg [(3'h5):(1'h0)] reg1924 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1923 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1922 = (1'h0);
  reg [(2'h3):(1'h0)] reg1921 = (1'h0);
  reg [(3'h6):(1'h0)] reg1919 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1918 = (1'h0);
  reg [(3'h5):(1'h0)] reg1915 = (1'h0);
  reg [(4'hc):(1'h0)] reg1913 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1912 = (1'h0);
  reg [(5'h16):(1'h0)] reg1910 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1903 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1899 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1898 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1897 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1891 = (1'h0);
  reg [(2'h2):(1'h0)] reg1893 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1892 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1881 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1888 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1887 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1886 = (1'h0);
  reg [(5'h14):(1'h0)] reg1882 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1881 = (1'h0);
  reg [(3'h6):(1'h0)] reg1875 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar1872 = (1'h0);
  reg [(5'h17):(1'h0)] reg1871 = (1'h0);
  reg [(4'ha):(1'h0)] reg1869 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1868 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1867 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1866 = (1'h0);
  reg [(5'h14):(1'h0)] reg1862 = (1'h0);
  reg [(5'h15):(1'h0)] reg1861 = (1'h0);
  reg [(4'he):(1'h0)] reg1860 = (1'h0);
  reg [(4'h9):(1'h0)] reg1856 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1853 = (1'h0);
  reg [(3'h6):(1'h0)] reg1852 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1850 = (1'h0);
  reg [(4'hb):(1'h0)] reg1848 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1847 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1846 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1845 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1844 = (1'h0);
  reg [(5'h14):(1'h0)] reg1843 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1842 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1841 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1839 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1837 = (1'h0);
  reg [(5'h19):(1'h0)] reg1835 = (1'h0);
  reg [(4'hf):(1'h0)] reg1834 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1833 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1830 = (1'h0);
  reg [(2'h3):(1'h0)] reg1829 = (1'h0);
  reg [(5'h13):(1'h0)] reg1828 = (1'h0);
  reg [(5'h10):(1'h0)] reg1827 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1826 = (1'h0);
  reg [(4'hd):(1'h0)] reg1825 = (1'h0);
  reg [(2'h2):(1'h0)] reg1823 = (1'h0);
  reg [(5'h10):(1'h0)] reg1817 = (1'h0);
  reg [(5'h16):(1'h0)] reg1815 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1812 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1811 = (1'h0);
  reg [(5'h14):(1'h0)] reg1809 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1808 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1806 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1805 = (1'h0);
  reg [(3'h6):(1'h0)] reg1804 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1802 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1796 = (1'h0);
  reg [(3'h6):(1'h0)] reg1795 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1794 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1792 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1790 = (1'h0);
  reg [(4'h8):(1'h0)] reg1789 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1784 = (1'h0);
  reg [(5'h12):(1'h0)] reg1781 = (1'h0);
  reg [(4'hb):(1'h0)] reg1780 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar1779 = (1'h0);
  assign y = {wire2165,
                 wire2078,
                 wire2077,
                 wire2059,
                 wire2015,
                 wire2007,
                 wire2006,
                 wire1909,
                 wire1907,
                 wire1906,
                 wire1905,
                 wire1904,
                 wire1810,
                 reg2194,
                 reg2193,
                 reg2192,
                 reg2189,
                 reg2187,
                 reg2183,
                 reg2182,
                 reg2180,
                 reg2179,
                 reg2177,
                 reg2175,
                 reg2174,
                 reg2173,
                 reg2172,
                 reg2168,
                 reg2167,
                 reg2164,
                 reg2163,
                 reg2162,
                 reg2158,
                 reg2156,
                 reg2155,
                 reg2151,
                 reg2147,
                 reg2146,
                 reg2143,
                 reg2141,
                 reg2139,
                 reg2137,
                 reg2135,
                 reg2132,
                 reg2130,
                 reg2127,
                 reg2121,
                 reg2120,
                 reg2119,
                 reg2114,
                 reg2113,
                 reg2111,
                 reg2110,
                 reg2108,
                 reg2107,
                 reg2103,
                 reg2102,
                 reg2100,
                 reg2097,
                 reg2096,
                 reg2089,
                 reg2088,
                 reg2085,
                 reg2083,
                 reg2082,
                 reg2081,
                 reg2073,
                 reg2069,
                 reg2063,
                 reg2062,
                 reg2058,
                 reg2057,
                 reg2052,
                 reg2049,
                 reg2047,
                 reg2044,
                 reg2043,
                 reg2040,
                 reg2038,
                 reg2034,
                 reg2031,
                 reg2030,
                 reg2028,
                 reg2022,
                 reg2021,
                 reg2020,
                 reg2019,
                 reg2012,
                 reg2011,
                 reg2010,
                 reg2009,
                 reg2004,
                 reg1997,
                 reg2001,
                 reg2000,
                 reg1993,
                 reg1992,
                 reg1990,
                 reg1989,
                 reg1988,
                 reg1987,
                 reg1985,
                 reg1984,
                 reg1980,
                 reg1978,
                 reg1977,
                 reg1975,
                 reg1972,
                 reg1971,
                 reg1970,
                 reg1969,
                 reg1968,
                 reg1966,
                 reg1965,
                 reg1961,
                 reg1960,
                 reg1959,
                 reg1958,
                 reg1957,
                 reg1955,
                 reg1953,
                 reg1952,
                 reg1951,
                 reg1949,
                 reg1948,
                 reg1947,
                 reg1946,
                 reg1945,
                 reg1944,
                 reg1942,
                 reg1941,
                 reg1937,
                 reg1933,
                 reg1932,
                 reg1931,
                 reg1930,
                 reg1927,
                 reg1926,
                 reg1920,
                 reg1917,
                 reg1916,
                 reg1914,
                 reg1911,
                 reg1908,
                 reg1902,
                 reg1901,
                 reg1900,
                 reg1896,
                 reg1895,
                 reg1894,
                 reg1891,
                 reg1890,
                 reg1872,
                 reg1889,
                 reg1885,
                 reg1884,
                 reg1883,
                 reg1880,
                 reg1879,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1874,
                 reg1873,
                 reg1870,
                 reg1865,
                 reg1864,
                 reg1863,
                 reg1859,
                 reg1858,
                 reg1857,
                 reg1855,
                 reg1854,
                 reg1851,
                 reg1849,
                 reg1811,
                 reg1840,
                 reg1838,
                 reg1836,
                 reg1832,
                 reg1831,
                 reg1824,
                 reg1822,
                 reg1821,
                 reg1820,
                 reg1819,
                 reg1818,
                 reg1816,
                 reg1814,
                 reg1813,
                 reg1807,
                 reg1803,
                 reg1801,
                 reg1800,
                 reg1799,
                 reg1798,
                 reg1797,
                 reg1793,
                 reg1791,
                 reg1788,
                 reg1787,
                 reg1786,
                 reg1785,
                 reg1783,
                 reg1782,
                 reg2191,
                 forvar2190,
                 reg2188,
                 reg2186,
                 reg2185,
                 reg2184,
                 forvar2181,
                 reg2178,
                 forvar2176,
                 reg2171,
                 forvar2170,
                 forvar2169,
                 reg2166,
                 reg2161,
                 reg2160,
                 forvar2159,
                 reg2157,
                 reg2154,
                 reg2153,
                 forvar2152,
                 reg2150,
                 reg2149,
                 reg2148,
                 reg2145,
                 reg2144,
                 reg2142,
                 reg2140,
                 reg2138,
                 forvar2136,
                 reg2134,
                 forvar2133,
                 reg2131,
                 reg2129,
                 reg2128,
                 reg2126,
                 reg2125,
                 forvar2124,
                 reg2123,
                 reg2122,
                 reg2118,
                 reg2117,
                 reg2116,
                 reg2115,
                 reg2104,
                 reg2112,
                 reg2109,
                 reg2106,
                 reg2105,
                 forvar2104,
                 reg2101,
                 reg2099,
                 reg2098,
                 forvar2095,
                 reg2094,
                 forvar2093,
                 reg2092,
                 reg2091,
                 reg2090,
                 forvar2087,
                 forvar2086,
                 reg2084,
                 reg2080,
                 forvar2079,
                 reg2076,
                 reg2075,
                 reg2074,
                 reg2072,
                 forvar2071,
                 reg2070,
                 reg2068,
                 forvar2067,
                 reg2066,
                 reg2065,
                 reg2064,
                 forvar2061,
                 forvar2060,
                 reg2056,
                 reg2055,
                 reg2054,
                 reg2053,
                 reg2051,
                 reg2050,
                 reg2048,
                 reg2046,
                 forvar2045,
                 reg2042,
                 reg2041,
                 reg2039,
                 forvar2037,
                 forvar2036,
                 reg2035,
                 reg2033,
                 reg2032,
                 forvar2029,
                 forvar2027,
                 reg2026,
                 reg2025,
                 forvar2024,
                 reg2023,
                 reg2018,
                 forvar2017,
                 reg2016,
                 reg2014,
                 reg2013,
                 reg2008,
                 reg2005,
                 reg2003,
                 reg2002,
                 reg1999,
                 reg1998,
                 forvar1997,
                 reg1996,
                 reg1995,
                 reg1994,
                 reg1991,
                 reg1986,
                 forvar1983,
                 forvar1982,
                 reg1981,
                 reg1979,
                 reg1976,
                 forvar1974,
                 reg1973,
                 reg1967,
                 forvar1964,
                 forvar1938,
                 reg1963,
                 reg1962,
                 reg1956,
                 reg1954,
                 reg1950,
                 reg1943,
                 reg1940,
                 reg1939,
                 reg1938,
                 forvar1936,
                 reg1935,
                 reg1934,
                 forvar1929,
                 forvar1928,
                 reg1925,
                 reg1924,
                 reg1923,
                 reg1922,
                 reg1921,
                 reg1919,
                 reg1918,
                 reg1915,
                 reg1913,
                 reg1912,
                 reg1910,
                 reg1903,
                 reg1899,
                 forvar1898,
                 forvar1897,
                 forvar1891,
                 reg1893,
                 reg1892,
                 reg1881,
                 reg1888,
                 forvar1887,
                 reg1886,
                 reg1882,
                 forvar1881,
                 reg1875,
                 forvar1872,
                 reg1871,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1862,
                 reg1861,
                 reg1860,
                 reg1856,
                 forvar1853,
                 reg1852,
                 reg1850,
                 reg1848,
                 reg1847,
                 reg1846,
                 reg1845,
                 reg1844,
                 reg1843,
                 reg1842,
                 forvar1841,
                 reg1839,
                 reg1837,
                 reg1835,
                 reg1834,
                 forvar1833,
                 reg1830,
                 reg1829,
                 reg1828,
                 reg1827,
                 reg1826,
                 reg1825,
                 reg1823,
                 reg1817,
                 reg1815,
                 reg1812,
                 forvar1811,
                 reg1809,
                 reg1808,
                 forvar1806,
                 reg1805,
                 reg1804,
                 reg1802,
                 forvar1796,
                 reg1795,
                 forvar1794,
                 reg1792,
                 reg1790,
                 reg1789,
                 reg1784,
                 reg1781,
                 reg1780,
                 forvar1779,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1779 = (1'h0); (forvar1779 < (3'h5)); forvar1779 = (forvar1779 + (1'h1)))
        begin
          reg1780 = ((wire1777[(4'h9):(2'h3)] ?
                  $signed($unsigned(wire1778)) : ((!{wire1776}) >> forvar1779[(4'he):(4'hb)])) ?
              $signed({$unsigned($signed(wire1774)),
                  ($signed((8'hbe)) ?
                      (wire1775 && forvar1779) : $signed(wire1776))}) : $unsigned($unsigned(((~&forvar1779) ?
                  (forvar1779 ? (8'ha9) : forvar1779) : $signed(wire1775)))));
          if (($signed((7'h43)) ?
              ($unsigned({wire1777[(5'h16):(5'h16)]}) ^~ ($signed(wire1778[(5'h12):(1'h0)]) ?
                  wire1777[(5'h12):(4'he)] : wire1777[(4'hb):(3'h4)])) : wire1774[(2'h2):(2'h2)]))
            begin
              reg1781 = (wire1775[(5'h18):(5'h12)] > $signed($signed(((|wire1776) ?
                  $signed(wire1777) : $unsigned(wire1775)))));
            end
          else
            begin
              reg1782 <= (~wire1776);
              reg1783 <= $unsigned(($unsigned($signed($signed(reg1781))) > (forvar1779 ?
                  {(reg1780 ?
                          wire1777 : reg1781)} : $signed($signed(forvar1779)))));
              reg1784 = wire1777;
            end
          reg1785 <= ($signed($signed(wire1775)) ?
              (|$unsigned($signed($signed(forvar1779)))) : $signed(wire1776[(3'h7):(2'h2)]));
          reg1786 <= ($unsigned(wire1774[(3'h7):(2'h2)]) + {({(reg1781 ?
                          wire1774 : reg1780),
                      (!wire1777),
                      {wire1774}} ?
                  wire1776 : (-reg1785[(3'h7):(3'h4)]))});
          if (wire1774[(3'h7):(3'h6)])
            begin
              reg1787 <= reg1785;
              reg1788 <= (8'haa);
            end
          else
            begin
              reg1789 = reg1786[(5'h1e):(4'hb)];
              reg1790 = (reg1789[(1'h0):(1'h0)] ?
                  ({$unsigned(wire1778),
                      $unsigned($unsigned(wire1774))} | (({reg1785,
                      wire1775,
                      reg1787} || $unsigned(reg1789)) == (+(8'hb7)))) : ((~^reg1785) ?
                      (!$signed((8'ha4))) : wire1775));
              reg1791 <= $signed($signed((($unsigned(reg1783) ?
                      reg1782 : reg1788) ?
                  ((reg1786 ? wire1776 : wire1776) ?
                      reg1789[(2'h2):(1'h1)] : $unsigned(forvar1779)) : (+(^~(7'h4a))))));
              reg1792 = ($signed(reg1791) << ((reg1783[(1'h1):(1'h0)] ^~ reg1787) && (+reg1791)));
              reg1793 <= $unsigned((-((!(reg1792 ?
                  forvar1779 : wire1776)) == reg1786)));
            end
        end
      for (forvar1794 = (1'h0); (forvar1794 < (3'h4)); forvar1794 = (forvar1794 + (1'h1)))
        begin
          reg1795 = $signed($unsigned($signed({(reg1793 <= reg1785)})));
          for (forvar1796 = (1'h0); (forvar1796 < (2'h2)); forvar1796 = (forvar1796 + (1'h1)))
            begin
              reg1797 <= $signed($signed((({reg1783} < reg1786[(5'h1c):(4'hf)]) * ((&(8'hbf)) ?
                  reg1791[(4'h8):(3'h5)] : (reg1793 && (7'h53))))));
              reg1798 <= (^~{($signed((reg1792 + forvar1794)) ?
                      $unsigned({(7'h4d)}) : $signed((!forvar1796))),
                  (({reg1786, reg1789, (7'h57)} < (reg1788 ?
                          (8'hac) : reg1789)) ?
                      (+(reg1780 || (7'h55))) : {$unsigned(wire1776)})});
              reg1799 <= (~^forvar1779[(4'hc):(4'hc)]);
              reg1800 <= forvar1794[(5'h16):(5'h12)];
              reg1801 <= $unsigned($signed($unsigned(wire1777)));
              reg1802 = $unsigned((^(~|(forvar1779[(5'h15):(5'h12)] ?
                  $signed(reg1786) : $unsigned(forvar1794)))));
              reg1803 <= $signed((((reg1791 && (7'h43)) - $signed(reg1797)) << (~^(8'haf))));
            end
          reg1804 = (~$signed($signed(reg1783)));
          reg1805 = reg1786[(1'h1):(1'h0)];
          for (forvar1806 = (1'h0); (forvar1806 < (1'h1)); forvar1806 = (forvar1806 + (1'h1)))
            begin
              reg1807 <= reg1786;
            end
          reg1808 = ($unsigned(reg1788[(3'h5):(1'h1)]) << $unsigned($signed(reg1790)));
        end
      reg1809 = reg1782;
    end
  assign wire1810 = $unsigned($unsigned($unsigned($signed(reg1783[(4'hb):(4'h8)]))));
  always
    @(posedge clk) begin
      if ({((!$signed(((8'ha6) ?
              wire1775 : wire1774))) ^~ reg1787[(4'hd):(4'h8)])})
        begin
          for (forvar1811 = (1'h0); (forvar1811 < (3'h6)); forvar1811 = (forvar1811 + (1'h1)))
            begin
              reg1812 = (reg1799 ?
                  $unsigned((^$signed($signed(wire1810)))) : (^(({reg1799} ?
                          (wire1777 ? reg1798 : reg1788) : (reg1791 ?
                              (8'ha2) : wire1778)) ?
                      ($unsigned(reg1807) ?
                          (reg1791 ?
                              reg1799 : forvar1811) : $signed(reg1785)) : (8'hbf))));
              reg1813 <= (($unsigned({$unsigned(wire1810),
                      ((7'h42) ? reg1787 : (8'ha6))}) ?
                  ((wire1810[(3'h4):(2'h3)] ^~ (reg1799 ?
                      reg1788 : (8'ha7))) ~^ $unsigned(wire1776[(1'h1):(1'h1)])) : reg1797[(4'hc):(4'hb)]) << (reg1798 ?
                  ({reg1782, (reg1807 ? reg1800 : reg1797)} ?
                      $unsigned((^~(7'h45))) : ((wire1777 - reg1791) ?
                          forvar1811[(4'ha):(4'h9)] : wire1810[(2'h2):(1'h1)])) : reg1807[(4'hb):(1'h0)]));
              reg1814 <= ((((((8'ha1) != wire1774) ?
                          (reg1798 <= reg1801) : (wire1777 ?
                              wire1776 : reg1787)) >= ($signed((7'h4d)) ?
                          wire1777[(4'hc):(3'h5)] : (~(8'h9f)))) ?
                      wire1776 : {{reg1803, (reg1807 | reg1791), {reg1807}}}) ?
                  {($signed((&wire1810)) ?
                          $signed(((7'h54) ?
                              wire1777 : reg1782)) : {$signed((8'h9c))}),
                      $unsigned($unsigned((!reg1783)))} : ({$unsigned((~|reg1785)),
                      ({reg1807} ?
                          reg1787[(4'h9):(3'h6)] : {(7'h4b)})} * (&($signed(reg1786) & wire1810[(4'hf):(4'hd)]))));
              reg1815 = (^~wire1778[(1'h1):(1'h1)]);
              reg1816 <= reg1801;
            end
          if (reg1807)
            begin
              reg1817 = (|reg1800);
              reg1818 <= (reg1801[(4'hc):(3'h6)] ?
                  (^$signed((|(^~reg1785)))) : {(|($unsigned(reg1815) + (reg1803 >>> reg1785))),
                      {$unsigned($signed((7'h4c))), (8'hb3)}});
              reg1819 <= ($signed(reg1816) > (!reg1793[(1'h1):(1'h0)]));
              reg1820 <= {{(reg1785[(1'h0):(1'h0)] || ($signed(reg1793) > (&reg1797))),
                      ($signed((reg1799 | reg1814)) ?
                          (~|(forvar1811 > reg1816)) : reg1782),
                      $signed(((|forvar1811) && $signed((8'ha3))))}};
              reg1821 <= $signed($unsigned(forvar1811));
              reg1822 <= $signed(($signed(((reg1797 ? (7'h44) : reg1786) ?
                      $signed(reg1799) : (7'h47))) ?
                  reg1812[(3'h6):(2'h2)] : (reg1821[(2'h3):(1'h0)] ?
                      ((reg1819 ?
                          (7'h41) : reg1812) >>> (+reg1803)) : (reg1801 ?
                          (wire1810 >>> reg1797) : (forvar1811 * reg1791)))));
            end
          else
            begin
              reg1818 <= reg1818;
              reg1819 <= (({$signed($signed(reg1815))} << ($signed({(7'h4f)}) ?
                      (+(reg1818 ?
                          reg1785 : reg1822)) : $signed((reg1798 || (8'hbe))))) ?
                  reg1785[(3'h5):(1'h0)] : (~|reg1817[(4'he):(4'hb)]));
              reg1820 <= reg1786[(5'h1f):(4'h8)];
              reg1823 = reg1820;
              reg1824 <= (~^reg1801[(5'h1d):(4'hb)]);
              reg1825 = $signed((({(wire1774 ?
                          reg1803 : reg1818)} > reg1813[(2'h3):(2'h2)]) ?
                  $unsigned($unsigned($signed(reg1807))) : reg1783[(4'hc):(4'hb)]));
            end
          if ($unsigned((reg1801[(4'hc):(4'h8)] ?
              reg1814 : ($unsigned($unsigned(reg1798)) + $unsigned((reg1798 ?
                  reg1818 : wire1774))))))
            begin
              reg1826 = reg1820[(5'h14):(3'h7)];
              reg1827 = (reg1782[(4'hb):(1'h0)] > ((~^reg1814[(4'hc):(3'h7)]) << $unsigned(($unsigned(reg1817) ?
                  $signed(reg1816) : reg1825[(3'h4):(2'h3)]))));
              reg1828 = reg1813[(1'h1):(1'h1)];
              reg1829 = ((~$signed(reg1815[(3'h6):(3'h5)])) - $unsigned(reg1816));
              reg1830 = ($signed($signed(reg1803[(4'hb):(3'h6)])) ?
                  (($unsigned({reg1823}) <<< reg1791) != ((~|reg1786) <<< ((reg1823 ?
                      (7'h53) : reg1782) + reg1814))) : $unsigned(reg1785[(3'h4):(3'h4)]));
              reg1831 <= reg1787[(4'hb):(4'ha)];
            end
          else
            begin
              reg1826 = (~^$signed((reg1801 | wire1776[(3'h7):(1'h1)])));
              reg1831 <= ($signed(reg1800[(3'h5):(3'h5)]) < wire1776);
            end
          reg1832 <= $unsigned(({$unsigned((reg1782 ? (8'hae) : reg1818)),
                  (reg1800[(4'h9):(2'h2)] + (&reg1830))} ?
              {reg1825[(3'h7):(3'h5)]} : $unsigned((((7'h41) >> (8'hbd)) != (7'h52)))));
          for (forvar1833 = (1'h0); (forvar1833 < (3'h6)); forvar1833 = (forvar1833 + (1'h1)))
            begin
              reg1834 = ($signed($signed(reg1819)) + $unsigned(wire1777));
              reg1835 = $unsigned(((&$unsigned($signed(reg1813))) != reg1813));
              reg1836 <= reg1797[(5'h1c):(4'h8)];
              reg1837 = reg1812;
              reg1838 <= (~&((reg1814 || ((reg1820 ?
                      wire1810 : reg1830) ^~ (8'hb6))) ?
                  reg1826[(4'hb):(3'h6)] : {$unsigned(((7'h47) <= reg1834))}));
              reg1839 = {((((reg1793 == reg1822) >>> (|reg1801)) + (~^{reg1800,
                      (8'hbf),
                      wire1777})) * (wire1776[(2'h3):(2'h2)] ?
                      reg1827 : (reg1819[(2'h3):(2'h3)] ?
                          $unsigned(reg1831) : reg1814))),
                  (($unsigned(reg1816[(5'h10):(4'ha)]) & (!$unsigned(wire1777))) ?
                      (~|($signed(reg1837) ^ $signed(reg1799))) : reg1834[(1'h0):(1'h0)])};
              reg1840 <= reg1829;
            end
          for (forvar1841 = (1'h0); (forvar1841 < (2'h3)); forvar1841 = (forvar1841 + (1'h1)))
            begin
              reg1842 = {(reg1840 | $unsigned(wire1778)),
                  reg1836,
                  $unsigned((($unsigned(reg1814) << (reg1791 ?
                      reg1801 : reg1815)) ^ (^~reg1820[(5'h1b):(4'hc)])))};
              reg1843 = {(($signed($signed(reg1836)) > $signed(reg1812[(4'hb):(4'h8)])) ?
                      ((|(reg1819 ^~ reg1831)) ~^ $signed(wire1774)) : reg1838),
                  wire1778[(3'h4):(2'h2)],
                  {$unsigned((-(reg1797 <= reg1831))),
                      (~reg1819[(4'h8):(3'h4)]),
                      $unsigned($unsigned((reg1798 - reg1842)))}};
              reg1844 = (reg1827 - (({reg1819} ?
                  ((8'hb6) >> reg1843[(2'h3):(2'h3)]) : reg1782[(4'hf):(2'h3)]) >> ((^~{reg1798,
                  reg1788}) ^~ {$unsigned(reg1821), (~&reg1799)})));
              reg1845 = ($unsigned((reg1837 ~^ reg1837[(4'ha):(4'h9)])) ?
                  {(reg1814[(4'hf):(2'h2)] ?
                          $unsigned(reg1840) : reg1791[(5'h14):(4'he)])} : reg1830[(5'h15):(5'h11)]);
              reg1846 = ($unsigned($unsigned(($signed(reg1829) ?
                  reg1814[(4'hb):(1'h1)] : {(8'hb7),
                      reg1827,
                      wire1775}))) && ((7'h58) ?
                  (reg1803 > $unsigned($unsigned(reg1814))) : (~&({(8'h9c),
                      reg1836} == (&reg1801)))));
              reg1847 = ($signed((reg1839 ?
                      $signed((reg1787 >> (8'hbd))) : {((8'hae) ^ reg1826)})) ?
                  ({reg1817} || $unsigned((((8'ha8) ^~ reg1785) << reg1823[(2'h2):(1'h1)]))) : ({reg1822,
                      ($unsigned(wire1775) != (reg1813 ?
                          reg1835 : reg1843))} >= reg1807));
            end
          reg1848 = $unsigned((~(-reg1832)));
        end
      else
        begin
          reg1811 <= (reg1835 == ($unsigned((reg1783[(3'h7):(3'h4)] <<< {wire1775,
                  reg1839})) ?
              {((wire1775 ? reg1845 : (7'h42)) ?
                      reg1846[(4'hf):(4'h9)] : $signed(forvar1841)),
                  ((reg1819 ? reg1843 : reg1837) ~^ (reg1836 ?
                      reg1797 : reg1787)),
                  $signed(reg1823)} : $signed($unsigned(reg1791[(4'he):(4'h9)]))));
          reg1813 <= reg1831;
          reg1815 = ((+(((reg1832 ? reg1819 : wire1774) ?
                      $unsigned((8'h9e)) : (reg1785 - reg1811)) ?
                  (&(-(8'ha7))) : reg1783)) ?
              reg1835 : reg1820);
          reg1816 <= reg1834;
          reg1817 = ((~($unsigned((+reg1811)) + reg1835[(5'h10):(4'he)])) ?
              $signed(reg1816) : (($signed($unsigned(wire1810)) ?
                      ((|reg1834) ?
                          {reg1829,
                              reg1785,
                              (8'ha3)} : (reg1814 << reg1837)) : {(reg1813 <<< reg1825),
                          (^~(7'h4a))}) ?
                  reg1829 : $signed($signed($signed(reg1815)))));
        end
      reg1849 <= reg1838[(5'h1a):(5'h10)];
      reg1850 = (^~($unsigned($signed(reg1801)) ?
          $unsigned((wire1810 | $signed(forvar1833))) : reg1800[(1'h1):(1'h0)]));
      reg1851 <= {(^(((~&(7'h46)) ^~ $unsigned(reg1839)) >= reg1822[(3'h4):(2'h3)]))};
    end
  always
    @(posedge clk) begin
      reg1852 = (~^((reg1822 < $unsigned({(7'h49)})) ?
          (~^{reg1785[(3'h6):(2'h2)]}) : (($signed(reg1807) != reg1814[(4'hb):(2'h3)]) * $signed(reg1787[(3'h5):(3'h4)]))));
      for (forvar1853 = (1'h0); (forvar1853 < (2'h3)); forvar1853 = (forvar1853 + (1'h1)))
        begin
          reg1854 <= (($signed((reg1836 ?
              (+reg1793) : (reg1788 ?
                  reg1797 : (7'h52)))) & ($signed((reg1820 || reg1849)) ?
              $unsigned(reg1851) : $unsigned(reg1820))) >>> $unsigned({reg1782,
              $signed((~|reg1800))}));
          reg1855 <= $signed($unsigned((~&((~&reg1820) > (|(8'hb0))))));
          reg1856 = $unsigned((^reg1852[(2'h3):(1'h0)]));
          if ({wire1777[(3'h5):(1'h0)],
              $signed($unsigned($signed((~|reg1838))))})
            begin
              reg1857 <= (-(7'h45));
            end
          else
            begin
              reg1857 <= (~|reg1855);
              reg1858 <= {$signed((8'hb4)),
                  (^((((8'hbf) ? reg1852 : (7'h46)) != $unsigned(reg1832)) ?
                      (reg1786 ?
                          (reg1791 >> (7'h51)) : $signed(reg1840)) : $unsigned(reg1813[(4'hb):(2'h2)]))),
                  (^reg1816[(5'h15):(4'h8)])};
              reg1859 <= reg1816;
              reg1860 = reg1832[(3'h4):(2'h3)];
              reg1861 = ($unsigned(reg1832) ?
                  $unsigned(reg1785) : $unsigned(($signed($unsigned((7'h49))) <= {$unsigned((7'h44)),
                      $unsigned(reg1836)})));
            end
          reg1862 = (~^wire1778[(4'ha):(1'h0)]);
        end
      if (reg1840[(4'h8):(3'h5)])
        begin
          if (reg1854)
            begin
              reg1863 <= ($unsigned(reg1831[(2'h2):(2'h2)]) | ($signed({$signed(wire1810),
                      wire1774[(4'hd):(4'hb)]}) ?
                  ($unsigned((reg1798 ^ (8'hbc))) * $unsigned({reg1782,
                      reg1855})) : wire1810));
              reg1864 <= $signed((reg1811[(1'h1):(1'h0)] ?
                  ((((8'hac) ?
                      reg1851 : wire1777) <<< (8'hb7)) ^~ (((8'hb3) >= reg1859) ?
                      $signed(reg1824) : (|reg1855))) : {(~&$signed(wire1776)),
                      (reg1849[(3'h6):(2'h3)] ?
                          $unsigned(reg1816) : {reg1788, reg1857}),
                      (^~(!reg1819))}));
              reg1865 <= ((8'hb8) > reg1787);
              reg1866 = ((reg1807[(1'h0):(1'h0)] ?
                  (~|(~reg1862[(4'hf):(4'h9)])) : $unsigned({{(8'hb0)},
                      reg1816[(5'h11):(5'h10)],
                      {(7'h42),
                          reg1818}})) - $signed($signed($unsigned((reg1860 >> (7'h49))))));
              reg1867 = reg1865;
              reg1868 = ({(reg1819 & $signed(reg1818)),
                      $unsigned($signed(reg1852[(3'h4):(2'h2)])),
                      reg1799} ?
                  reg1786 : (((^~$signed(reg1852)) ?
                          $signed((8'hba)) : (!(~^(8'hac)))) ?
                      reg1783[(4'ha):(4'ha)] : wire1776[(3'h4):(2'h3)]));
              reg1869 = (~|$signed(($signed(((8'had) ? reg1800 : reg1840)) ?
                  $signed((reg1857 ? (8'hbf) : reg1811)) : ({(7'h47), (8'hac)} ?
                      reg1791[(5'h10):(4'hb)] : (^reg1793)))));
            end
          else
            begin
              reg1866 = (+(+(~&$signed({reg1787, reg1814, wire1778}))));
              reg1870 <= ($unsigned($unsigned(reg1868[(1'h0):(1'h0)])) && {$unsigned($signed(reg1863[(1'h1):(1'h1)])),
                  wire1777[(5'h17):(1'h1)]});
            end
          reg1871 = {((reg1818[(1'h1):(1'h1)] ?
                  (&((7'h55) >= (8'h9c))) : {$signed(reg1820)}) ~^ reg1861),
              {(reg1798[(1'h1):(1'h1)] <= (-(~reg1855))),
                  (|(reg1854[(4'hf):(1'h1)] - reg1813[(3'h5):(3'h5)]))}};
          for (forvar1872 = (1'h0); (forvar1872 < (1'h0)); forvar1872 = (forvar1872 + (1'h1)))
            begin
              reg1873 <= ($unsigned($signed(reg1856)) ?
                  (~^((((7'h57) ? reg1866 : reg1787) >>> (reg1860 != reg1860)) ?
                      $unsigned((reg1861 ^~ reg1861)) : (reg1867[(1'h1):(1'h0)] + $signed(reg1862)))) : (~(&$signed($unsigned(reg1813)))));
              reg1874 <= $signed(reg1856);
              reg1875 = (~{reg1874, (wire1778[(3'h4):(2'h2)] <= wire1810)});
              reg1876 <= $signed($unsigned(((((8'hb8) ?
                  reg1798 : reg1851) >= (reg1860 ?
                  reg1799 : reg1800)) >> (reg1787[(4'ha):(4'h8)] ^ (reg1821 + reg1816)))));
              reg1877 <= reg1868[(1'h0):(1'h0)];
              reg1878 <= $signed(reg1860);
            end
          reg1879 <= (reg1782 > $signed($unsigned(wire1810)));
          reg1880 <= (7'h54);
          for (forvar1881 = (1'h0); (forvar1881 < (2'h2)); forvar1881 = (forvar1881 + (1'h1)))
            begin
              reg1882 = ($signed(reg1859[(4'h9):(1'h0)]) ?
                  reg1854 : (~&{((reg1836 ?
                          (8'ha2) : reg1876) & $unsigned(reg1866))}));
              reg1883 <= (reg1869 ~^ $unsigned(((reg1868 ?
                  (reg1800 + reg1813) : (~reg1879)) ~^ reg1818[(1'h1):(1'h1)])));
              reg1884 <= ((+($unsigned((reg1870 ? reg1798 : (8'h9d))) ?
                  {reg1859[(3'h6):(3'h6)]} : $unsigned((|reg1879)))) - {forvar1853,
                  ($signed((reg1797 ?
                      reg1793 : forvar1872)) * reg1813[(4'hc):(3'h5)]),
                  reg1786});
              reg1885 <= ($signed(reg1822[(3'h5):(2'h3)]) ?
                  $signed(reg1836[(4'hc):(1'h1)]) : forvar1872[(1'h0):(1'h0)]);
              reg1886 = {((^~((reg1858 * reg1798) ?
                          $unsigned(reg1785) : (reg1880 >>> forvar1872))) ?
                      (($signed(reg1862) <<< $signed(reg1879)) ?
                          reg1785[(4'h9):(4'h8)] : $unsigned((reg1856 ?
                              reg1885 : forvar1853))) : ((((8'haf) > forvar1872) + (reg1865 ?
                          reg1885 : forvar1881)) == reg1859[(3'h4):(3'h4)])),
                  ({$signed((reg1878 ? reg1803 : reg1874)),
                      (((8'hb8) >>> reg1798) ?
                          reg1793[(4'hd):(4'hc)] : {reg1838, reg1861}),
                      ((reg1875 >= reg1882) ?
                          {(7'h51), wire1776} : (reg1878 ?
                              reg1869 : reg1783))} || $signed({$unsigned(reg1854),
                      $signed(reg1788)})),
                  ((8'haf) && $unsigned(((^reg1803) ?
                      (reg1832 ? reg1824 : (7'h4c)) : $unsigned(reg1854))))};
            end
          for (forvar1887 = (1'h0); (forvar1887 < (1'h1)); forvar1887 = (forvar1887 + (1'h1)))
            begin
              reg1888 = $unsigned((+(reg1836[(3'h7):(3'h6)] ?
                  {((8'hbe) || reg1870),
                      (reg1861 ~^ reg1883),
                      reg1879[(2'h3):(2'h2)]} : (^~reg1801))));
              reg1889 <= $signed(reg1824[(1'h1):(1'h1)]);
            end
        end
      else
        begin
          reg1866 = (($unsigned($signed((^(8'ha0)))) << $unsigned((wire1810[(1'h0):(1'h0)] ?
              $unsigned(reg1836) : (+(7'h4d))))) << (8'ha7));
          if (($unsigned(reg1871) ? (^~reg1860[(4'he):(3'h4)]) : reg1868))
            begin
              reg1867 = {(~^($signed(reg1873) == (!(|(8'hbe))))),
                  {(wire1810 | reg1803[(4'h9):(3'h4)]),
                      $unsigned((~^reg1855)),
                      (reg1807 ? $unsigned((8'ha1)) : (|{wire1777, reg1821}))}};
              reg1870 <= ($signed(reg1874) == {$signed(reg1787)});
              reg1871 = $unsigned($unsigned($unsigned({reg1800})));
              reg1872 <= $unsigned(reg1832[(2'h2):(2'h2)]);
            end
          else
            begin
              reg1870 <= {(reg1816[(5'h17):(5'h16)] ?
                      {$signed(((8'ha1) ? reg1869 : reg1840)),
                          (~&$signed(reg1851)),
                          $unsigned($signed(reg1788))} : {reg1882[(5'h10):(1'h1)]}),
                  (reg1855[(4'h9):(1'h1)] ?
                      ((^~reg1849[(2'h3):(1'h0)]) ?
                          wire1778 : ($signed(reg1871) ?
                              {reg1787,
                                  reg1849,
                                  (7'h49)} : $signed(reg1863))) : ($unsigned($unsigned(reg1885)) <= reg1838))};
              reg1871 = $signed((~^reg1868[(1'h1):(1'h0)]));
              reg1872 <= $unsigned(((^~$unsigned((reg1814 ?
                  reg1862 : reg1885))) || ($signed($signed(reg1782)) ?
                  (((8'hb7) ?
                      reg1861 : reg1876) ~^ reg1857) : (reg1786[(4'hf):(4'h9)] >= $unsigned(reg1793)))));
              reg1875 = (~^(!{$unsigned((^~forvar1887))}));
            end
          reg1881 = $signed($unsigned((!((&reg1849) ?
              reg1862[(2'h2):(1'h0)] : (~reg1882)))));
          reg1883 <= $unsigned((~&((reg1882[(3'h6):(1'h1)] | (reg1861 ^~ reg1882)) ~^ $signed(reg1831[(1'h0):(1'h0)]))));
        end
      if ((^((|reg1868) ? {reg1872} : reg1885)))
        begin
          reg1890 <= (-(8'hb0));
          reg1891 <= $unsigned((!({reg1840[(5'h11):(1'h1)],
              reg1803} >> reg1877[(3'h5):(2'h3)])));
          if ($unsigned({$unsigned(((reg1855 ? reg1860 : (8'hb6)) ?
                  reg1862[(4'h9):(1'h1)] : reg1783[(2'h3):(1'h1)]))}))
            begin
              reg1892 = (^~(~^reg1886[(5'h10):(3'h5)]));
              reg1893 = reg1864[(5'h10):(2'h2)];
            end
          else
            begin
              reg1894 <= $signed(reg1814[(4'hf):(4'ha)]);
              reg1895 <= {reg1813,
                  (((^~(reg1820 ? reg1797 : reg1782)) ?
                          $unsigned((~^forvar1872)) : $unsigned(reg1857)) ?
                      $signed(reg1858[(3'h5):(3'h4)]) : (^$unsigned(((8'hbf) | reg1874)))),
                  ((reg1873[(4'h8):(1'h1)] && {(!reg1881),
                      {reg1884, reg1881}}) ^~ ($signed((reg1881 ?
                          forvar1887 : wire1776)) ?
                      $signed((|reg1893)) : ($unsigned(reg1814) == ((8'ha6) ?
                          reg1869 : reg1889))))};
              reg1896 <= (reg1816 ?
                  (wire1778[(4'hc):(3'h7)] & $unsigned($unsigned(((8'hba) ?
                      reg1820 : reg1819)))) : (reg1893 >> (reg1788 ?
                      reg1811[(1'h1):(1'h0)] : {{reg1877, (8'hbe), reg1854}})));
            end
        end
      else
        begin
          reg1890 <= $unsigned(reg1836[(3'h6):(1'h0)]);
          for (forvar1891 = (1'h0); (forvar1891 < (1'h0)); forvar1891 = (forvar1891 + (1'h1)))
            begin
              reg1892 = reg1880[(1'h1):(1'h0)];
            end
          reg1893 = (~|$signed((reg1797 << $signed((^reg1831)))));
          reg1894 <= (~^(!$signed((!(wire1778 <<< reg1875)))));
        end
      for (forvar1897 = (1'h0); (forvar1897 < (2'h2)); forvar1897 = (forvar1897 + (1'h1)))
        begin
          for (forvar1898 = (1'h0); (forvar1898 < (1'h0)); forvar1898 = (forvar1898 + (1'h1)))
            begin
              reg1899 = reg1896[(5'h13):(3'h5)];
              reg1900 <= {$signed({($signed(reg1793) ?
                          (reg1869 - reg1872) : reg1859),
                      $signed($signed(reg1875)),
                      ({(8'hb1)} ? (~^reg1876) : (reg1858 >>> reg1875))})};
              reg1901 <= $signed((!$signed($signed($signed(reg1854)))));
              reg1902 <= $unsigned(reg1797);
              reg1903 = reg1803;
            end
        end
    end
  assign wire1904 = ($unsigned((+reg1877)) ?
                        $signed(reg1801) : ($signed(reg1851) ?
                            ({$signed((7'h50)),
                                (|reg1857),
                                reg1819[(4'hf):(4'h8)]} | {(reg1824 + reg1901),
                                reg1864,
                                reg1824[(1'h1):(1'h1)]}) : ((wire1778[(4'h9):(2'h3)] >> $unsigned(reg1878)) ~^ wire1777)));
  assign wire1905 = reg1864[(5'h10):(3'h4)];
  assign wire1906 = $signed(wire1810);
  assign wire1907 = (^$signed((-$signed((reg1840 ? reg1878 : (7'h42))))));
  always
    @(posedge clk) begin
      reg1908 <= (reg1818[(2'h3):(2'h2)] && ((reg1880[(1'h1):(1'h0)] ^ reg1786) <= $signed(((^reg1865) ?
          $unsigned(reg1864) : (reg1901 << reg1864)))));
    end
  assign wire1909 = $unsigned($signed((((reg1885 || reg1880) ?
                            reg1803[(3'h6):(1'h1)] : (~^reg1849)) ?
                        $signed((&wire1777)) : ((reg1857 <= reg1836) ?
                            $signed(wire1907) : $unsigned((8'ha3))))));
  always
    @(posedge clk) begin
      if ($unsigned((reg1816[(3'h4):(1'h1)] ?
          {(reg1876 ? reg1884 : reg1876[(4'hd):(1'h0)])} : $signed(reg1873))))
        begin
          reg1910 = reg1891[(3'h6):(1'h0)];
          reg1911 <= $signed((reg1879 | (8'h9e)));
          reg1912 = $unsigned(reg1877[(3'h4):(2'h3)]);
          reg1913 = $signed(((reg1811[(1'h1):(1'h0)] ?
                  $signed($signed((7'h45))) : (reg1851 ?
                      $unsigned(reg1890) : reg1786[(5'h1c):(5'h11)])) ?
              wire1909 : $unsigned((reg1801[(4'hd):(1'h0)] && wire1775[(5'h10):(4'hc)]))));
          reg1914 <= $unsigned(({{reg1902[(5'h19):(5'h18)], $signed(wire1810)},
              (+$unsigned((8'hb3)))} | {((reg1894 | reg1877) ?
                  (8'ha9) : (~&reg1787))}));
          reg1915 = {reg1785,
              (reg1851[(3'h5):(2'h3)] ?
                  ($signed($unsigned(reg1857)) + (reg1891[(4'ha):(3'h6)] <= (wire1810 ?
                      wire1777 : reg1819))) : ($unsigned($unsigned(reg1901)) ^ $unsigned((~wire1810))))};
        end
      else
        begin
          if ($signed($signed({$unsigned((reg1884 || wire1774))})))
            begin
              reg1910 = $unsigned(({{reg1822[(4'ha):(3'h4)],
                      (reg1878 ? reg1832 : reg1914),
                      (~reg1831)},
                  $signed($unsigned(reg1859))} & (^$signed((~^(8'hbb))))));
              reg1912 = $unsigned($unsigned((reg1798 <= reg1824)));
              reg1914 <= ($unsigned(reg1803[(4'hf):(2'h2)]) >= (reg1857[(3'h4):(2'h3)] <<< ($unsigned($unsigned(reg1788)) >= wire1904[(4'hc):(3'h6)])));
              reg1915 = $signed(reg1801[(1'h1):(1'h0)]);
              reg1916 <= $unsigned($unsigned($unsigned($signed(reg1813[(4'ha):(1'h0)]))));
              reg1917 <= reg1891;
              reg1918 = $unsigned((^$signed($signed((^~reg1782)))));
            end
          else
            begin
              reg1910 = $unsigned((reg1816 ?
                  reg1787 : $unsigned(reg1787[(2'h2):(1'h0)])));
            end
          if ({reg1911[(4'h9):(2'h2)]})
            begin
              reg1919 = reg1791;
              reg1920 <= reg1858;
              reg1921 = $signed(($unsigned((^~(7'h41))) & $signed($unsigned({reg1910,
                  reg1895}))));
              reg1922 = $signed($unsigned(wire1905));
              reg1923 = ($unsigned((7'h44)) >> (7'h57));
              reg1924 = wire1904;
              reg1925 = reg1911;
            end
          else
            begin
              reg1919 = ((&{wire1778[(3'h6):(1'h1)],
                      $unsigned(wire1907),
                      $unsigned(reg1803[(1'h1):(1'h1)])}) ?
                  $signed((((|reg1813) ?
                          (reg1880 ? reg1895 : reg1908) : (reg1917 ?
                              reg1902 : reg1919)) ?
                      reg1797 : reg1819)) : (((^(reg1849 ~^ reg1921)) ?
                      (reg1798[(1'h1):(1'h0)] && (8'h9e)) : (~^(wire1776 && wire1907))) || (&($unsigned(reg1891) ?
                      (~&wire1905) : reg1885[(5'h11):(3'h6)]))));
              reg1921 = ({((^~(8'hbe)) ?
                      reg1797 : ($unsigned(reg1877) ?
                          ((8'h9e) <<< reg1917) : wire1905))} != (^((^~wire1776) <= $signed($signed(reg1908)))));
              reg1926 <= ($signed({{$unsigned(reg1878), reg1890},
                      reg1807[(2'h3):(2'h3)],
                      (^~wire1907[(1'h0):(1'h0)])}) ?
                  ({reg1914[(4'hb):(3'h7)], reg1878[(3'h4):(1'h0)]} ?
                      reg1821 : $unsigned({(reg1801 ? reg1920 : reg1822),
                          (&reg1900),
                          (7'h42)})) : reg1821[(5'h12):(2'h3)]);
            end
          reg1927 <= reg1824[(2'h3):(2'h3)];
        end
      for (forvar1928 = (1'h0); (forvar1928 < (1'h1)); forvar1928 = (forvar1928 + (1'h1)))
        begin
          for (forvar1929 = (1'h0); (forvar1929 < (2'h3)); forvar1929 = (forvar1929 + (1'h1)))
            begin
              reg1930 <= (reg1902 >>> ((reg1914[(1'h1):(1'h1)] ^ (~&(~|reg1872))) < ($unsigned((~|reg1786)) ?
                  (~&reg1787) : $signed($signed(reg1820)))));
              reg1931 <= $signed(((|reg1801[(5'h16):(5'h10)]) ^~ (!(8'ha5))));
              reg1932 <= $signed((wire1904[(5'h10):(3'h7)] | reg1917));
              reg1933 <= $unsigned({$unsigned(reg1788),
                  ($unsigned((forvar1929 ? reg1920 : (8'hb5))) >= ({reg1890,
                      reg1786,
                      forvar1929} << ((8'ha3) ? reg1822 : reg1832))),
                  reg1858[(3'h5):(3'h5)]});
              reg1934 = (-$unsigned(forvar1929[(1'h0):(1'h0)]));
            end
          reg1935 = (reg1831[(1'h0):(1'h0)] <<< $unsigned(reg1916));
          for (forvar1936 = (1'h0); (forvar1936 < (1'h1)); forvar1936 = (forvar1936 + (1'h1)))
            begin
              reg1937 <= reg1822[(4'ha):(3'h5)];
            end
        end
      if ((8'ha0))
        begin
          if ((-$unsigned(reg1838[(1'h1):(1'h1)])))
            begin
              reg1938 = {(8'hb7)};
              reg1939 = ((+(($signed(reg1813) ?
                  $unsigned(forvar1929) : reg1797) >= $unsigned($signed(reg1831)))) | $signed((~^reg1819[(1'h1):(1'h0)])));
              reg1940 = reg1854;
              reg1941 <= $signed((+{$unsigned({(8'hb0), (7'h4a), reg1854}),
                  (reg1930[(1'h1):(1'h0)] ?
                      $signed(reg1939) : reg1838[(5'h1e):(5'h1c)]),
                  $signed($signed(reg1786))}));
              reg1942 <= $unsigned($unsigned(((8'ha3) >>> (7'h54))));
              reg1943 = reg1864;
            end
          else
            begin
              reg1938 = reg1865[(3'h6):(1'h1)];
              reg1939 = $unsigned((wire1777[(3'h4):(1'h1)] ?
                  ($unsigned((wire1776 || reg1914)) ^~ ({reg1939,
                          reg1942,
                          reg1883} ?
                      (~&(7'h4d)) : reg1818[(1'h1):(1'h1)])) : ($unsigned((^~wire1778)) ?
                      (reg1801 ?
                          reg1884[(2'h3):(2'h3)] : wire1810[(3'h6):(1'h0)]) : ((wire1909 == (8'hba)) && (reg1896 || reg1818)))));
              reg1940 = reg1782;
              reg1941 <= ($unsigned($unsigned((8'hbc))) <= ($unsigned(reg1821) >= reg1913[(2'h3):(2'h2)]));
              reg1943 = reg1890[(3'h4):(2'h3)];
              reg1944 <= (wire1777[(2'h3):(2'h2)] ?
                  {(~|((reg1799 ? (7'h53) : reg1896) ?
                          reg1801[(1'h1):(1'h0)] : $signed(reg1939)))} : ($unsigned(((~&(8'ha3)) | reg1923)) >>> {($signed(reg1849) > reg1787[(4'hf):(4'hc)]),
                      ($signed(reg1849) ? $unsigned(reg1943) : (~reg1783))}));
            end
          if ((reg1840[(4'hd):(2'h2)] ?
              $signed((~|(|$signed(reg1896)))) : (((reg1920 ?
                          (reg1799 << (7'h47)) : {wire1906, wire1905}) ?
                      (reg1890[(2'h3):(2'h3)] == reg1927) : $signed((reg1894 * reg1935))) ?
                  reg1858[(5'h12):(2'h2)] : $unsigned(((+reg1873) ?
                      (~&wire1810) : (|reg1914))))))
            begin
              reg1945 <= $signed($unsigned((^(reg1863[(1'h1):(1'h1)] | reg1944[(3'h7):(2'h2)]))));
              reg1946 <= (reg1910[(5'h15):(1'h1)] >> {reg1914,
                  $unsigned(($unsigned(wire1906) ?
                      reg1821 : reg1800[(5'h12):(1'h0)]))});
              reg1947 <= reg1924[(3'h4):(3'h4)];
              reg1948 <= (wire1777[(4'hb):(3'h4)] != wire1775);
              reg1949 <= ((reg1943[(3'h4):(3'h4)] + ((wire1810 ?
                  {reg1945,
                      reg1786,
                      reg1782} : $signed((7'h56))) & ((7'h4e) == reg1832[(2'h3):(2'h3)]))) ~^ $signed((reg1948 ?
                  reg1818[(2'h2):(1'h1)] : {(reg1921 ^ reg1822)})));
              reg1950 = (($signed(reg1883[(5'h10):(3'h6)]) ^~ $unsigned({(!reg1807),
                  $signed(reg1912)})) != {($unsigned(reg1917[(4'hd):(4'hc)]) + $signed((^~reg1811)))});
            end
          else
            begin
              reg1950 = reg1910[(5'h16):(4'he)];
            end
          if ($signed(($unsigned(((7'h53) >> (~^reg1940))) != (^($unsigned(reg1900) ^ {wire1904})))))
            begin
              reg1951 <= {({reg1924,
                      ((wire1810 << reg1800) ?
                          reg1798 : (reg1797 ? (7'h48) : reg1948)),
                      $signed(reg1949)} == $unsigned((reg1832 > reg1924[(3'h5):(2'h2)])))};
              reg1952 <= (reg1885[(2'h2):(1'h1)] ?
                  $unsigned(($signed((reg1831 >>> reg1924)) ?
                      ($signed(reg1908) ~^ ((8'hb7) ?
                          reg1872 : wire1776)) : ({forvar1936,
                          reg1912} >> $signed(reg1786)))) : (reg1859[(1'h1):(1'h0)] ?
                      $signed({$unsigned(reg1883),
                          (wire1775 ? reg1818 : (7'h4b)),
                          (reg1919 * reg1913)}) : {$signed((^~reg1935))}));
              reg1953 <= $signed(reg1785);
              reg1954 = {reg1793[(5'h1a):(5'h13)],
                  ($signed(($unsigned(reg1923) ?
                          reg1943 : $unsigned((8'ha3)))) ?
                      ($unsigned((|reg1923)) || reg1807) : {wire1904,
                          ((wire1777 ? reg1944 : reg1900) ?
                              $unsigned(reg1921) : ((7'h56) <<< reg1858)),
                          {(reg1944 >>> reg1821), $unsigned((7'h54))}})};
              reg1955 <= reg1872;
            end
          else
            begin
              reg1951 <= $signed((^reg1937));
              reg1954 = (^~($signed($unsigned($unsigned(reg1814))) ?
                  ($signed(reg1822) ?
                      ((7'h56) + (reg1895 ?
                          reg1854 : reg1925)) : {((7'h52) >>> reg1912)}) : $signed(reg1836[(4'hc):(2'h3)])));
            end
          if ($signed($signed($signed($unsigned($signed(reg1880))))))
            begin
              reg1956 = reg1814;
              reg1957 <= reg1916;
              reg1958 <= $unsigned(reg1955);
            end
          else
            begin
              reg1957 <= (&$signed((|(reg1807 ^~ reg1945))));
              reg1958 <= ($signed((reg1798[(1'h1):(1'h0)] ?
                      reg1870[(5'h14):(5'h10)] : $signed({reg1836,
                          wire1776}))) ?
                  (((~|reg1912[(1'h0):(1'h0)]) - ((reg1889 ?
                          (8'ha2) : reg1955) ?
                      (&reg1939) : $unsigned(reg1816))) >> forvar1928) : wire1775[(5'h13):(3'h6)]);
              reg1959 <= (reg1894[(5'h10):(4'ha)] ?
                  (reg1954 != $signed($unsigned($signed((7'h53))))) : {(-($unsigned(reg1957) == reg1919[(2'h2):(2'h2)])),
                      reg1877[(4'he):(4'h9)]});
              reg1960 <= $signed((reg1877[(1'h1):(1'h0)] << (~(+$unsigned(reg1900)))));
              reg1961 <= $unsigned((~(+$unsigned($unsigned(reg1803)))));
              reg1962 = (reg1788 < reg1931);
              reg1963 = (8'ha0);
            end
        end
      else
        begin
          for (forvar1938 = (1'h0); (forvar1938 < (1'h1)); forvar1938 = (forvar1938 + (1'h1)))
            begin
              reg1939 = $unsigned((reg1921 ?
                  ($unsigned($unsigned(reg1814)) ?
                      $unsigned((forvar1928 < reg1925)) : reg1951[(3'h6):(2'h3)]) : (!($signed((7'h49)) ?
                      reg1933[(1'h0):(1'h0)] : {(7'h44), reg1889, (7'h44)}))));
              reg1941 <= ($unsigned(($signed(reg1870[(4'hd):(4'hd)]) ?
                      (8'h9c) : $unsigned({reg1911, reg1831}))) ?
                  $unsigned($signed($signed(reg1858[(2'h3):(1'h0)]))) : reg1950);
              reg1942 <= {reg1945[(2'h2):(2'h2)],
                  $unsigned(($signed({reg1927, wire1777, reg1872}) ?
                      ((~|reg1857) ?
                          ((8'hb8) ?
                              forvar1928 : reg1818) : (~|reg1858)) : $unsigned($signed(wire1810))))};
              reg1944 <= reg1885[(4'h9):(3'h7)];
              reg1950 = (^~reg1962[(2'h3):(1'h0)]);
            end
          if ((~|reg1854[(4'hf):(4'hd)]))
            begin
              reg1951 <= (((reg1962 || ($signed(reg1900) ?
                  reg1798 : {reg1921,
                      reg1949,
                      (8'ha0)})) | $unsigned(($signed(reg1951) > (reg1801 * (7'h49))))) - (reg1915 ?
                  $signed(reg1912[(4'hd):(3'h6)]) : (~($unsigned((7'h40)) ?
                      (reg1807 ? reg1800 : (8'ha2)) : (^reg1962)))));
              reg1954 = ($signed(($unsigned({(7'h52), reg1948}) == (^~(reg1894 ?
                  reg1952 : (8'hb9))))) - ({wire1776, $unsigned((~|wire1905))} ?
                  reg1884[(1'h1):(1'h1)] : {reg1857}));
              reg1956 = (+{{$unsigned(reg1910[(3'h7):(3'h6)])}});
            end
          else
            begin
              reg1951 <= $unsigned(reg1786[(5'h17):(1'h0)]);
              reg1952 <= $unsigned($unsigned({reg1916, reg1854, reg1923}));
              reg1953 <= ($unsigned(reg1921[(1'h0):(1'h0)]) ?
                  (8'ha3) : reg1797[(5'h16):(4'h8)]);
              reg1954 = ($signed((reg1799 >>> reg1838[(4'h8):(3'h6)])) <= $signed(reg1859[(3'h7):(1'h0)]));
            end
          reg1957 <= reg1787;
        end
      if (($signed($signed((reg1915 ?
          (8'hab) : (reg1849 ? (8'hbd) : reg1925)))) ^ reg1854))
        begin
          for (forvar1964 = (1'h0); (forvar1964 < (1'h0)); forvar1964 = (forvar1964 + (1'h1)))
            begin
              reg1965 <= reg1941[(4'hf):(1'h1)];
              reg1966 <= reg1961[(3'h4):(1'h1)];
              reg1967 = {reg1819[(3'h6):(1'h1)],
                  ((~{reg1896, $signed(wire1906), $unsigned(reg1949)}) ?
                      $signed($unsigned($unsigned(reg1959))) : ((~&$signed(reg1965)) ~^ reg1793[(5'h17):(4'hd)]))};
              reg1968 <= reg1849;
              reg1969 <= (reg1849[(3'h7):(3'h5)] ?
                  reg1782 : reg1832[(1'h0):(1'h0)]);
              reg1970 <= reg1818;
              reg1971 <= $unsigned($unsigned((~^(~^(~^reg1807)))));
            end
          reg1972 <= (^~$signed((($unsigned((8'hba)) ?
              (7'h42) : $signed((7'h53))) == (|reg1932))));
        end
      else
        begin
          for (forvar1964 = (1'h0); (forvar1964 < (3'h6)); forvar1964 = (forvar1964 + (1'h1)))
            begin
              reg1965 <= $signed((^(~^{(reg1958 + reg1855)})));
              reg1966 <= (~(({(reg1801 ? (7'h42) : reg1813),
                      reg1946[(3'h5):(3'h4)]} ?
                  ((reg1872 ^~ reg1807) ?
                      wire1909[(4'hb):(3'h6)] : {reg1858,
                          wire1775,
                          (7'h48)}) : reg1917[(5'h15):(3'h7)]) != (((reg1896 <= reg1785) + (reg1791 ~^ wire1906)) ?
                  ((reg1952 ? reg1872 : reg1894) ?
                      (reg1924 < reg1970) : {reg1889,
                          reg1958,
                          reg1951}) : $unsigned($unsigned(reg1851)))));
              reg1967 = forvar1936;
              reg1968 <= {$signed($signed({(reg1968 >>> reg1820)})),
                  $signed((reg1854 ^~ reg1917[(5'h16):(5'h13)]))};
            end
          reg1969 <= (((((reg1949 ? forvar1936 : reg1787) ?
                      reg1800[(3'h4):(1'h1)] : (|(8'hb1))) ?
                  $unsigned($unsigned(reg1901)) : ((reg1822 <<< reg1880) * reg1941[(4'h9):(4'h9)])) ?
              (^$signed((!reg1793))) : $unsigned(($unsigned(reg1971) ?
                  reg1945[(5'h10):(4'he)] : $signed(reg1945)))) == $signed((~|$signed((~reg1949)))));
          reg1973 = reg1960;
          for (forvar1974 = (1'h0); (forvar1974 < (3'h6)); forvar1974 = (forvar1974 + (1'h1)))
            begin
              reg1975 <= $unsigned({reg1970[(4'ha):(4'h9)]});
              reg1976 = reg1970;
              reg1977 <= reg1913;
              reg1978 <= ($unsigned((($unsigned(reg1910) ?
                          (~&reg1976) : {reg1923, reg1824, wire1909}) ?
                      (7'h4d) : $signed((reg1799 + reg1791)))) ?
                  $unsigned($unsigned(reg1876[(5'h11):(2'h2)])) : $unsigned(($signed($signed(reg1914)) ~^ reg1901)));
              reg1979 = $unsigned(reg1967);
              reg1980 <= $signed(reg1917[(4'hf):(4'h9)]);
            end
        end
      reg1981 = (&(&$signed((^~(reg1966 * reg1863)))));
      for (forvar1982 = (1'h0); (forvar1982 < (2'h2)); forvar1982 = (forvar1982 + (1'h1)))
        begin
          for (forvar1983 = (1'h0); (forvar1983 < (3'h5)); forvar1983 = (forvar1983 + (1'h1)))
            begin
              reg1984 <= $signed(reg1970);
              reg1985 <= {{(~reg1957)}};
              reg1986 = reg1879[(4'ha):(3'h6)];
              reg1987 <= reg1836[(4'hc):(4'hb)];
              reg1988 <= $signed((~&$signed(reg1783)));
              reg1989 <= $signed(($signed(reg1956) ^~ $signed((reg1942[(2'h2):(2'h2)] == (reg1946 - (7'h40))))));
            end
          reg1990 <= reg1877[(4'h8):(3'h7)];
          reg1991 = {reg1931, ((forvar1964 || $unsigned(reg1840)) < reg1820)};
          reg1992 <= $signed(reg1863);
          reg1993 <= $signed($signed($unsigned($signed($unsigned((8'hb3))))));
        end
      if (reg1787[(4'hb):(4'h9)])
        begin
          reg1994 = $signed(((reg1884 ?
              $unsigned({reg1987}) : reg1954) >= reg1782));
          reg1995 = $signed($unsigned($signed((7'h58))));
          reg1996 = $unsigned({reg1798});
          for (forvar1997 = (1'h0); (forvar1997 < (1'h0)); forvar1997 = (forvar1997 + (1'h1)))
            begin
              reg1998 = $signed((reg1922 ?
                  ({$unsigned(reg1865)} ?
                      (~&$unsigned((8'hb6))) : {$unsigned(reg1915),
                          ((7'h41) * wire1907),
                          forvar1928[(3'h7):(2'h3)]}) : $signed($signed(reg1941))));
              reg1999 = $signed((~&reg1883[(5'h19):(3'h5)]));
              reg2000 <= {reg1935};
            end
          reg2001 <= reg1939[(5'h11):(4'he)];
          reg2002 = reg1947;
          reg2003 = $unsigned(reg1901[(2'h2):(1'h0)]);
        end
      else
        begin
          if (((reg1836[(4'h8):(2'h2)] ?
                  (~$unsigned((|reg1967))) : (&($unsigned(reg1911) - (reg1902 ?
                      reg1884 : reg2000)))) ?
              ((($signed(reg1920) ?
                      (reg1799 ? reg1840 : (8'hb1)) : (+(8'hbc))) ?
                  reg1988 : $signed((reg1961 > reg1791))) == reg1832) : (({$unsigned((8'had)),
                          (reg1890 ? (7'h45) : reg1883),
                          (reg1838 == reg1820)} ?
                      (8'h9f) : $signed((reg1857 == reg1884))) ?
                  $signed(reg1786) : (reg1895[(2'h2):(2'h2)] * reg1876))))
            begin
              reg1997 <= reg1932[(3'h7):(3'h6)];
              reg1998 = reg1910;
            end
          else
            begin
              reg1997 <= (reg1953 * (($signed($unsigned(reg1975)) ?
                      ($signed((8'hba)) ?
                          reg1949 : forvar1936[(5'h11):(1'h1)]) : $unsigned((reg1916 == reg1901))) ?
                  (8'hb2) : reg1851));
              reg2000 <= reg1894[(4'h8):(3'h5)];
              reg2001 <= ((8'ha1) || wire1774);
              reg2002 = reg1926[(3'h4):(2'h3)];
              reg2003 = $unsigned(reg1798[(1'h0):(1'h0)]);
              reg2004 <= ($unsigned(reg1876) ?
                  ($unsigned(((reg1883 ~^ reg1940) > (reg1787 || reg1991))) ?
                      $signed((~&reg1991[(4'hd):(4'h8)])) : ((7'h50) ?
                          reg1855[(4'h8):(4'h8)] : $unsigned({reg1891,
                              (7'h50),
                              (8'h9f)}))) : $unsigned($unsigned({reg1836[(4'hb):(2'h2)]})));
            end
          reg2005 = $signed(reg1975);
        end
    end
  assign wire2006 = {(+(reg1872 & ((reg1908 < reg1832) ?
                            $signed(reg1941) : ((8'ha7) ? (7'h49) : reg1945)))),
                        (~^(reg1984 + {$unsigned(reg1824),
                            (reg1855 ? reg1785 : reg1945)}))};
  assign wire2007 = ((wire1774 << (($signed(reg1908) ?
                        $signed(reg2001) : reg1788[(3'h6):(2'h2)]) > {$signed((8'ha8)),
                        reg1877[(1'h1):(1'h0)],
                        $unsigned(wire1777)})) ^~ {((|reg1980) && ($signed(wire1777) ?
                            (reg1968 ?
                                reg1851 : reg1972) : $unsigned(reg1840))),
                        $unsigned(((reg1785 & (7'h49)) ?
                            $signed((8'hb6)) : reg1884))});
  always
    @(posedge clk) begin
      reg2008 = ($signed((-reg1957[(2'h2):(1'h1)])) - (~^(reg1902 ?
          $unsigned(reg1857) : ($signed(reg1966) && ((7'h43) - reg1953)))));
      reg2009 <= ($unsigned((reg1896[(5'h10):(2'h3)] >> $signed(reg1889[(5'h16):(5'h12)]))) == ((reg1908[(4'he):(4'hb)] << (((8'hb8) ?
                  (8'haa) : reg1916) ?
              (8'hb0) : $unsigned(reg1987))) ?
          reg1927 : reg1989[(4'hd):(4'hc)]));
      reg2010 <= (^$unsigned(reg1783[(4'hb):(3'h6)]));
      reg2011 <= $signed($unsigned(((wire1776[(3'h5):(2'h3)] >= reg1908) ?
          $signed({reg1859, wire2007}) : (7'h49))));
      reg2012 <= (wire2006[(4'hd):(2'h3)] ^ ((($signed(reg1785) >= reg1857) & (^{reg1863,
          reg1932})) << (~|reg1855)));
      reg2013 = $unsigned((!($unsigned((~|reg1937)) * $unsigned($unsigned(reg1969)))));
      if ($signed({$unsigned(reg1894[(3'h6):(1'h0)]), reg1872[(1'h1):(1'h1)]}))
        begin
          reg2014 = $unsigned(($signed(wire2007[(4'hc):(3'h6)]) ?
              reg1949 : {((reg1959 ? reg1838 : reg1883) ? (-reg1926) : (7'h51)),
                  reg1927[(3'h5):(3'h4)],
                  reg1820}));
        end
      else
        begin
          reg2014 = reg1955;
        end
    end
  assign wire2015 = ($unsigned(reg1914) ?
                        (reg1880 ?
                            (7'h51) : $signed(((reg1896 ?
                                (8'hab) : reg1836) << {reg1953,
                                (7'h4c),
                                (7'h41)}))) : $unsigned({(8'hac),
                            reg1836,
                            {reg1859[(3'h4):(1'h0)], reg1894, (^reg1955)}}));
  always
    @(posedge clk) begin
      reg2016 = reg1955;
      for (forvar2017 = (1'h0); (forvar2017 < (1'h1)); forvar2017 = (forvar2017 + (1'h1)))
        begin
          if ((reg1820 ?
              (~&$signed(reg1814)) : $signed((+{{reg1819, reg1865},
                  reg2016,
                  reg1873}))))
            begin
              reg2018 = (reg1840[(4'hd):(1'h1)] | ({$signed($signed(reg1883)),
                  (8'ha5)} & $unsigned((^~{reg1931, reg1931, reg1797}))));
            end
          else
            begin
              reg2019 <= reg1968;
              reg2020 <= reg1972[(5'h12):(3'h6)];
            end
          reg2021 <= reg1874[(4'ha):(4'h9)];
        end
      reg2022 <= wire2015;
    end
  always
    @(posedge clk) begin
      reg2023 = (($unsigned((~&wire1810)) ?
          ($unsigned((7'h52)) ?
              $signed($signed(reg1894)) : reg1870) : ($signed((reg1914 ?
                  reg1953 : reg1854)) ?
              ((reg2010 ^~ (8'hbb)) & reg2000) : reg1854[(5'h10):(4'he)])) >= ($signed({{wire1907,
              reg2009}}) != (((~&reg1890) == (reg1872 ? (7'h56) : reg2012)) ?
          {reg1831[(4'h8):(1'h1)]} : $unsigned((~wire1777)))));
      for (forvar2024 = (1'h0); (forvar2024 < (3'h4)); forvar2024 = (forvar2024 + (1'h1)))
        begin
          reg2025 = $unsigned($unsigned((+($unsigned(reg1958) <<< (reg1990 & reg1952)))));
          reg2026 = $signed(($signed(reg1946) ?
              {($unsigned(reg1863) * reg1870)} : (reg2025 ?
                  {$unsigned(reg1977), (~reg1783)} : ((reg1984 ?
                          wire2007 : (7'h4b)) ?
                      {wire1774} : $signed(reg1970)))));
        end
      for (forvar2027 = (1'h0); (forvar2027 < (3'h5)); forvar2027 = (forvar2027 + (1'h1)))
        begin
          reg2028 <= (~|(((^~$signed(reg1970)) ?
                  wire1810 : $unsigned((reg1961 >> reg1926))) ?
              $signed($unsigned(reg2023)) : (wire1909 ?
                  reg1977 : reg1958[(2'h3):(2'h3)])));
          for (forvar2029 = (1'h0); (forvar2029 < (1'h0)); forvar2029 = (forvar2029 + (1'h1)))
            begin
              reg2030 <= (~|{$unsigned({(reg1824 + reg1822),
                      (reg1813 | reg1822),
                      $unsigned(reg1865)}),
                  $unsigned({reg1941[(4'hd):(4'hb)]}),
                  (-$unsigned(reg1863[(4'h9):(3'h7)]))});
              reg2031 <= reg1865[(1'h1):(1'h0)];
              reg2032 = (|(~&reg1917[(5'h18):(3'h4)]));
              reg2033 = reg1840;
              reg2034 <= (reg1944 + reg1896[(1'h0):(1'h0)]);
            end
        end
      reg2035 = reg1813;
      for (forvar2036 = (1'h0); (forvar2036 < (3'h4)); forvar2036 = (forvar2036 + (1'h1)))
        begin
          for (forvar2037 = (1'h0); (forvar2037 < (1'h0)); forvar2037 = (forvar2037 + (1'h1)))
            begin
              reg2038 <= reg1824;
              reg2039 = {(reg1958[(4'hf):(2'h2)] ? reg1908 : reg1958),
                  (wire1907 ?
                      ((^~(reg1895 <<< reg2031)) ?
                          (reg2025 ?
                              ((8'ha8) ?
                                  reg2030 : reg1946) : (~^(7'h4d))) : ((reg1993 ?
                                  (8'ha6) : reg1902) ?
                              reg1858[(4'hb):(1'h1)] : $unsigned(forvar2029))) : reg1959),
                  reg1814[(3'h6):(1'h0)]};
              reg2040 <= {(&$unsigned((^reg1879[(4'he):(4'hd)]))),
                  {{forvar2029[(2'h3):(1'h1)], $signed($unsigned(reg2031))},
                      reg2035[(4'ha):(4'h9)],
                      {reg1807, $unsigned(((8'h9d) != reg1854))}}};
              reg2041 = ($signed($signed($signed(reg2004))) ?
                  (reg1873[(3'h6):(1'h1)] ?
                      $signed($signed($signed(wire1777))) : $signed($unsigned({reg1801}))) : (|reg1811));
              reg2042 = reg1807[(1'h0):(1'h0)];
              reg2043 <= (({({(8'ha4), (7'h57), reg1821} ?
                          (reg1997 >= reg1942) : (reg1793 >>> reg1993)),
                      $signed($unsigned(reg1819))} << (((reg2001 ?
                              reg1911 : (8'hb5)) ?
                          $signed(reg1799) : (+wire2006)) ?
                      $signed((&(8'ha9))) : (reg1980[(5'h15):(5'h12)] ?
                          (forvar2037 <<< reg2035) : (7'h44)))) ?
                  reg1874[(4'he):(4'hc)] : $signed({($signed(reg1788) ?
                          $signed((7'h41)) : (reg1917 ? reg1873 : reg1849))}));
              reg2044 <= (|reg1799);
            end
          for (forvar2045 = (1'h0); (forvar2045 < (1'h0)); forvar2045 = (forvar2045 + (1'h1)))
            begin
              reg2046 = (reg2033[(4'h9):(3'h6)] ?
                  $signed($unsigned((^~(|reg1975)))) : reg2030[(2'h3):(1'h0)]);
              reg2047 <= (reg1858 ^~ reg1859);
            end
          reg2048 = reg1917;
          reg2049 <= (^((^($signed(reg2038) != wire1810[(4'hb):(3'h7)])) != $signed(($unsigned(reg1785) - $unsigned(reg1911)))));
          if ($signed($unsigned(wire1905[(1'h1):(1'h1)])))
            begin
              reg2050 = $unsigned((~(8'hb2)));
              reg2051 = (reg1821[(5'h13):(4'hd)] ^ $signed($signed($unsigned(wire2007[(3'h5):(2'h2)]))));
              reg2052 <= wire2015;
              reg2053 = reg1948[(2'h3):(2'h3)];
            end
          else
            begin
              reg2050 = reg1920;
              reg2052 <= reg1941;
              reg2053 = ((~($signed(reg1785) ?
                      reg2034[(4'hc):(2'h3)] : reg2023)) ?
                  $unsigned(((-$signed(reg1832)) ?
                      $unsigned((reg1840 < reg2039)) : (&(+reg1965)))) : {reg1947[(4'h8):(2'h2)]});
              reg2054 = reg2038;
              reg2055 = $signed($unsigned($unsigned((reg2038 ?
                  reg1813 : $signed(reg1879)))));
              reg2056 = reg1870[(3'h7):(3'h6)];
            end
        end
      reg2057 <= {{reg1914[(2'h2):(1'h0)], reg1787[(4'he):(4'h8)]}, (7'h44)};
      reg2058 <= reg1798[(2'h2):(1'h0)];
    end
  assign wire2059 = ($unsigned($signed(reg1975)) == $unsigned($signed(((reg1813 ?
                            (8'hbf) : reg2001) ?
                        $signed(reg2038) : ((8'haf) ? reg1985 : wire1907)))));
  always
    @(posedge clk) begin
      for (forvar2060 = (1'h0); (forvar2060 < (3'h4)); forvar2060 = (forvar2060 + (1'h1)))
        begin
          for (forvar2061 = (1'h0); (forvar2061 < (2'h3)); forvar2061 = (forvar2061 + (1'h1)))
            begin
              reg2062 <= (+$unsigned(($signed($unsigned(wire1905)) ?
                  $unsigned(reg1993) : $unsigned({reg1865,
                      reg1891,
                      reg1911}))));
              reg2063 <= {reg2062[(2'h3):(1'h0)],
                  (7'h4b),
                  $unsigned(((reg1807 ?
                      (reg1945 ?
                          (7'h4d) : reg1930) : (~|reg2038)) & ((reg1813 + reg1819) && reg2028)))};
              reg2064 = (~$unsigned($signed((8'hb9))));
              reg2065 = (~|($unsigned(((+wire1775) ?
                      (reg1785 >> reg1969) : $unsigned(reg2057))) ?
                  (!(^~reg2047)) : (8'hab)));
            end
          reg2066 = $signed($signed((~^(|$signed(reg2044)))));
          for (forvar2067 = (1'h0); (forvar2067 < (2'h2)); forvar2067 = (forvar2067 + (1'h1)))
            begin
              reg2068 = (~^reg1926[(4'h9):(2'h2)]);
              reg2069 <= $unsigned($unsigned(forvar2067[(2'h3):(1'h1)]));
              reg2070 = (~&((~&reg1980) | $unsigned(reg1997[(3'h5):(1'h0)])));
            end
          for (forvar2071 = (1'h0); (forvar2071 < (1'h0)); forvar2071 = (forvar2071 + (1'h1)))
            begin
              reg2072 = {(~((^(reg1970 || reg1916)) ?
                      ((reg1791 <<< (8'ha6)) ^ (reg1946 ?
                          reg1798 : reg1836)) : $unsigned((reg1858 ?
                          forvar2060 : reg1948)))),
                  $signed((reg2065[(4'he):(2'h3)] >= $signed($unsigned(reg1930)))),
                  (reg1989[(4'h9):(3'h7)] ?
                      ((reg1932[(4'h9):(4'h9)] ?
                          $signed(wire2059) : (reg1971 ?
                              reg2052 : reg1993)) && ($unsigned(reg1966) ?
                          wire1778[(1'h0):(1'h0)] : (reg1977 >>> (8'ha3)))) : (wire1774[(2'h3):(2'h2)] ?
                          reg2012[(3'h7):(3'h4)] : wire1778[(1'h1):(1'h1)]))};
              reg2073 <= {(-(8'had))};
              reg2074 = reg1864[(4'hf):(4'hb)];
              reg2075 = (~^reg1801);
              reg2076 = (reg1970 <<< reg1891[(2'h2):(1'h1)]);
            end
        end
    end
  assign wire2077 = reg1800[(5'h12):(2'h2)];
  assign wire2078 = $unsigned((({$signed(wire2077)} < ((wire2015 ?
                            reg1797 : reg2019) > (reg2063 ?
                            wire2077 : reg1978))) ?
                        (reg1889 >>> reg1894[(4'he):(4'ha)]) : (($unsigned((8'h9d)) ~^ wire2015[(2'h2):(1'h1)]) ?
                            {(!reg2028),
                                (~^wire2077)} : wire1777[(3'h7):(3'h7)])));
  always
    @(posedge clk) begin
      for (forvar2079 = (1'h0); (forvar2079 < (1'h1)); forvar2079 = (forvar2079 + (1'h1)))
        begin
          if (reg1872)
            begin
              reg2080 = $signed($signed($unsigned(($signed(reg1787) || $unsigned(reg1831)))));
              reg2081 <= reg2031;
              reg2082 <= (8'hba);
              reg2083 <= $unsigned($unsigned(reg2004[(4'he):(4'hc)]));
              reg2084 = reg1966[(5'h12):(4'h8)];
              reg2085 <= reg1811;
            end
          else
            begin
              reg2080 = $unsigned((reg1895 ?
                  ($signed($signed(reg1944)) >= reg1878) : $signed($unsigned((reg1814 ^~ reg1941)))));
              reg2081 <= $signed(($unsigned(reg1840[(4'hf):(1'h1)]) < (reg1946[(3'h6):(3'h5)] ?
                  (!(|(8'ha1))) : reg2010[(5'h15):(1'h0)])));
              reg2082 <= $signed((((|(^~reg2082)) ?
                      ((~&reg1937) >= $signed(reg1819)) : wire1810) ?
                  $unsigned(((|reg2052) * $signed(reg1831))) : $unsigned(((|reg1952) ?
                      ((7'h4d) + reg1896) : (~^reg1874)))));
              reg2083 <= {((reg1873[(4'h8):(4'h8)] ?
                      (+$signed(reg1955)) : ($signed(reg1803) <<< ((8'hb1) >= reg1877))) && reg1971)};
            end
        end
      for (forvar2086 = (1'h0); (forvar2086 < (3'h4)); forvar2086 = (forvar2086 + (1'h1)))
        begin
          for (forvar2087 = (1'h0); (forvar2087 < (1'h0)); forvar2087 = (forvar2087 + (1'h1)))
            begin
              reg2088 <= ($unsigned({{(reg1917 || (8'hb7)), (~&reg1945)},
                  {(wire1775 + reg1980)},
                  reg1858[(4'hc):(4'h8)]}) > $signed(reg1800[(1'h1):(1'h0)]));
              reg2089 <= $unsigned($signed(reg1793[(1'h1):(1'h0)]));
              reg2090 = (((wire2006[(3'h4):(1'h1)] + $unsigned($unsigned(reg1987))) ^ reg2020[(5'h18):(4'h8)]) ?
                  reg1824 : (((reg1926[(3'h4):(2'h3)] * (reg2084 > wire1778)) ~^ {(reg1793 - reg1873),
                      $unsigned((8'hbb)),
                      reg1920}) - $signed($signed($signed(reg1997)))));
              reg2091 = reg1944;
            end
          reg2092 = (^~$unsigned(($signed((!reg1889)) || (reg2081[(4'h9):(1'h1)] ?
              {reg1977, reg2049, reg2085} : (reg1782 << reg2031)))));
          for (forvar2093 = (1'h0); (forvar2093 < (1'h0)); forvar2093 = (forvar2093 + (1'h1)))
            begin
              reg2094 = reg1978[(2'h2):(2'h2)];
            end
          for (forvar2095 = (1'h0); (forvar2095 < (1'h1)); forvar2095 = (forvar2095 + (1'h1)))
            begin
              reg2096 <= wire2077[(3'h4):(2'h2)];
              reg2097 <= (~|reg2011);
              reg2098 = reg1927;
              reg2099 = reg2090;
              reg2100 <= {(reg2019[(1'h1):(1'h1)] || $unsigned((~&(reg2000 - reg2098)))),
                  ({(reg1854[(4'he):(1'h0)] ?
                          {reg2049, (8'hb5)} : reg2080[(3'h6):(2'h2)]),
                      (~^$unsigned(reg1953)),
                      ((reg2020 >>> reg1984) ?
                          $unsigned(reg1797) : reg1927)} >> (reg1971 ?
                      (((8'ha4) ?
                          reg1984 : reg2052) != (8'ha7)) : (reg2073 != $signed(reg2092))))};
              reg2101 = ((|(reg2062 - $signed({reg1858,
                  reg2019,
                  reg1859}))) ^~ ($signed(((-reg1840) ?
                      (reg1863 ^~ reg1993) : (~|reg1960))) ?
                  reg1821[(4'hb):(3'h5)] : reg2088[(5'h11):(3'h6)]));
            end
        end
      if ($unsigned((((reg1820[(5'h18):(5'h10)] ?
              (!reg1798) : wire1775[(3'h5):(1'h0)]) <= reg1811) ?
          reg1947[(3'h6):(3'h6)] : ($signed({reg2100,
              reg1997}) <= (|(&reg1838))))))
        begin
          reg2102 <= $unsigned($signed(reg2082[(5'h1c):(1'h0)]));
          reg2103 <= (($unsigned(($signed(reg1987) ?
                  reg1969[(5'h16):(5'h11)] : $unsigned(reg1785))) <<< $unsigned(reg1900)) ?
              (^$unsigned(((!reg2099) > (reg1971 - forvar2086)))) : (7'h45));
          for (forvar2104 = (1'h0); (forvar2104 < (2'h3)); forvar2104 = (forvar2104 + (1'h1)))
            begin
              reg2105 = reg2012;
              reg2106 = $unsigned($unsigned($signed((+(!reg2040)))));
              reg2107 <= reg1955[(5'h13):(3'h7)];
            end
          reg2108 <= ($unsigned($signed({reg1800, reg1930, $signed(reg1863)})) ?
              (8'h9e) : reg1997);
          if ({(~$unsigned(reg1877[(2'h3):(2'h2)])),
              reg1951[(3'h6):(2'h3)],
              (!($signed($unsigned(wire1777)) || $signed(reg1877[(5'h11):(4'hd)])))})
            begin
              reg2109 = $signed((reg2030 * reg2012[(3'h7):(3'h4)]));
              reg2110 <= (-$unsigned(({{(8'ha1), reg1953},
                      (-reg2107),
                      {(8'hba)}} ?
                  $signed(reg2089) : {$signed(reg2040), {reg1953, reg2062}})));
              reg2111 <= reg2084;
            end
          else
            begin
              reg2109 = (-reg1958[(3'h6):(3'h6)]);
              reg2112 = reg1889[(5'h1b):(2'h3)];
            end
        end
      else
        begin
          if ((~^reg2001))
            begin
              reg2104 = (8'haf);
              reg2107 <= ((~|(((reg1813 >> reg1824) | $unsigned(reg1788)) < (!{reg1908,
                      reg1803}))) ?
                  (^{$unsigned((reg1874 ?
                          (8'ha6) : reg1946))}) : (reg1863 - $signed(($signed((7'h48)) ?
                      {(7'h56)} : ((8'hb5) ^~ reg1786)))));
              reg2109 = ({(reg1798[(2'h2):(2'h2)] >>> ((reg1836 && reg1831) ?
                      {(8'ha1),
                          reg1849} : $signed(reg2111)))} != reg1786[(4'hf):(3'h4)]);
              reg2112 = $unsigned({(+((^reg1891) & (reg2044 + (8'hb8)))),
                  reg2097});
              reg2113 <= forvar2087;
            end
          else
            begin
              reg2102 <= $unsigned((($unsigned(reg1832[(3'h5):(1'h1)]) ?
                      $signed((reg1878 ? (8'h9d) : reg1975)) : reg1948) ?
                  reg1953 : reg2103[(3'h7):(2'h3)]));
              reg2104 = reg2104;
              reg2107 <= $signed($signed((7'h56)));
            end
          if (($unsigned(wire1905) ?
              wire1774[(4'hb):(1'h0)] : {((&$signed(wire2078)) >> ((reg2089 != reg1992) ?
                      (&reg2010) : (reg2069 ? reg1798 : reg2103))),
                  (|reg1884)}))
            begin
              reg2114 <= reg1890;
              reg2115 = reg2069;
              reg2116 = reg1968[(2'h3):(2'h3)];
              reg2117 = wire1909;
              reg2118 = (!(($signed((reg1863 ^ reg1916)) ?
                      reg1877[(5'h12):(4'h9)] : ((reg1985 ? reg2073 : reg2108) ?
                          (~&reg1836) : (|reg2113))) ?
                  reg2107 : $signed($signed(((7'h4f) || reg2069)))));
              reg2119 <= ($signed(reg1864) ?
                  {$signed({reg1980[(5'h15):(5'h11)], $unsigned(reg2004)}),
                      ($unsigned($signed((7'h4d))) ?
                          wire2077[(3'h7):(3'h5)] : reg2098[(1'h1):(1'h0)]),
                      reg1984[(5'h13):(1'h1)]} : ((($unsigned(reg2010) * (reg2022 ?
                          reg1797 : reg1874)) ?
                      (8'ha8) : reg1818[(1'h1):(1'h0)]) >= {($unsigned(reg2009) ^ (reg1787 ?
                          reg2043 : reg1977)),
                      reg1914,
                      ($unsigned((8'hb1)) >>> (|reg2011))}));
            end
          else
            begin
              reg2114 <= $unsigned({((reg1927 >>> ((8'hb5) ?
                          reg1902 : reg2081)) ?
                      ($unsigned(reg2069) ?
                          forvar2093[(3'h7):(3'h5)] : $unsigned(reg2062)) : reg1822[(4'h9):(3'h7)]),
                  $signed($unsigned(reg2090[(4'ha):(4'h9)])),
                  (reg1798[(2'h3):(1'h1)] ?
                      reg2052 : (reg1993[(5'h10):(4'hd)] ?
                          (reg1941 < reg2116) : reg1783[(4'h8):(1'h1)]))});
              reg2115 = (8'ha9);
              reg2119 <= {(reg1946[(5'h14):(5'h14)] && (((reg1902 ?
                          reg1965 : reg1916) ?
                      reg1977 : {reg1947, reg2118, reg1997}) <= reg1984)),
                  {(!reg1955[(5'h11):(4'hf)]), reg2021[(2'h3):(2'h3)]},
                  ((+reg1931) ?
                      ($signed($unsigned((7'h50))) && ((8'h9e) > $signed((8'hb5)))) : ({(reg1890 ?
                                  wire2007 : reg1849),
                              {reg2073},
                              wire1909[(2'h2):(1'h1)]} ?
                          (^~(reg1968 ? reg1816 : (8'ha1))) : (reg1821 ?
                              ((7'h4a) ? reg2110 : reg2096) : (|reg1947))))};
              reg2120 <= (8'haf);
              reg2121 <= reg1889[(2'h3):(2'h3)];
              reg2122 = reg1920;
            end
          reg2123 = (reg1874[(2'h3):(1'h1)] ?
              $signed($unsigned(({(8'h9d),
                  reg2121} < reg2092))) : $unsigned(reg1855[(4'h9):(2'h2)]));
          for (forvar2124 = (1'h0); (forvar2124 < (3'h4)); forvar2124 = (forvar2124 + (1'h1)))
            begin
              reg2125 = $signed((((reg2115 ?
                      $signed(forvar2079) : (reg2028 ?
                          reg1984 : (8'ha0))) == reg2123) ?
                  $unsigned(((reg1851 || reg2062) << (reg2028 - reg2122))) : (~^reg1953[(4'h9):(2'h3)])));
              reg2126 = reg2021[(2'h2):(2'h2)];
              reg2127 <= $unsigned(reg2117[(3'h7):(3'h6)]);
              reg2128 = (~^reg1822[(2'h3):(1'h0)]);
              reg2129 = reg1813;
              reg2130 <= ($signed(reg2111[(4'h8):(3'h4)]) < ((reg1945 & $signed((reg1971 || reg2097))) ?
                  reg1838[(4'h9):(2'h2)] : $signed(((~|(8'h9f)) | (&reg1870)))));
            end
          reg2131 = (^$signed((~&reg1874)));
        end
    end
  always
    @(posedge clk) begin
      reg2132 <= $signed(({reg2047[(4'hd):(1'h0)]} ?
          (~(reg1793 > reg2110[(1'h1):(1'h1)])) : $unsigned($unsigned($unsigned(reg1863)))));
      for (forvar2133 = (1'h0); (forvar2133 < (1'h1)); forvar2133 = (forvar2133 + (1'h1)))
        begin
          reg2134 = {$signed($unsigned(reg1818[(2'h2):(1'h0)])),
              reg1800,
              reg1885};
          reg2135 <= wire2077[(3'h4):(1'h0)];
          for (forvar2136 = (1'h0); (forvar2136 < (3'h5)); forvar2136 = (forvar2136 + (1'h1)))
            begin
              reg2137 <= ({(&$signed($signed(reg1859))),
                      reg2127[(5'h10):(3'h4)]} ?
                  wire1778[(4'he):(3'h6)] : {reg1890[(4'h8):(1'h0)]});
              reg2138 = ($signed(reg1816[(5'h11):(4'hf)]) ?
                  (~|(|$unsigned({reg1980,
                      reg1972,
                      (8'ha6)}))) : (((reg1937 > $signed(reg1863)) ?
                      reg2011 : (~^(reg2057 ?
                          (7'h40) : reg1895))) * ((+(&reg1889)) ?
                      ((reg1969 ? reg1873 : wire1774) ?
                          {(7'h43),
                              wire2015} : $signed(forvar2136)) : reg2097)));
              reg2139 <= (&reg1931[(5'h14):(4'hb)]);
              reg2140 = reg1933;
              reg2141 <= ($signed((({(7'h4d), (8'hbc)} ?
                          reg1791[(4'hc):(2'h2)] : (reg1970 ?
                              reg1977 : wire1907)) ?
                      ($signed(reg1990) > {(8'hbc)}) : (^~reg1787[(3'h4):(1'h0)]))) ?
                  $unsigned(reg1966[(5'h10):(5'h10)]) : $signed(wire1774));
              reg2142 = (^(~|$signed($unsigned($signed(wire1778)))));
              reg2143 <= (~&(wire2077[(4'h9):(2'h2)] ?
                  ($signed($signed(reg1859)) ^~ ((^~reg2119) | $signed(reg2043))) : (reg2020 - (!((8'h9c) ?
                      reg1787 : reg2088)))));
            end
          reg2144 = reg2009[(4'hd):(2'h2)];
          if ($signed(wire1810))
            begin
              reg2145 = (reg2139[(4'hf):(3'h5)] ?
                  reg1970 : ($unsigned((~|$unsigned(reg1873))) && $signed($unsigned((wire1907 ^ wire2078)))));
              reg2146 <= $unsigned($unsigned($unsigned($signed($signed(reg2083)))));
              reg2147 <= (^(reg2000 ?
                  $unsigned($signed(((7'h56) <<< reg1966))) : (~&(~|(reg2085 ?
                      (8'hb5) : reg2019)))));
              reg2148 = reg1855;
              reg2149 = (~$signed((reg2063 >>> $unsigned($signed((8'hac))))));
              reg2150 = (~$signed(reg2081));
              reg2151 <= (((8'hb9) ?
                      $signed(reg2083) : reg2127[(3'h6):(2'h2)]) ?
                  (~&$unsigned({(wire2006 ^ (7'h58)),
                      reg2147,
                      (-wire1778)})) : forvar2136[(3'h4):(1'h1)]);
            end
          else
            begin
              reg2145 = $signed((7'h43));
              reg2146 <= ($signed(($unsigned($signed(reg1985)) ?
                      $unsigned({reg1816}) : (^~$unsigned(reg1920)))) ?
                  wire1810[(3'h5):(2'h2)] : $signed((((reg1865 ?
                          (8'hb2) : reg2137) * (reg2028 ? (8'had) : reg1908)) ?
                      $unsigned((reg2069 + (8'hb9))) : reg2038[(4'h8):(2'h3)])));
              reg2147 <= (^~($unsigned((~|(reg1908 ? (8'hb0) : reg2149))) ?
                  (reg2040[(2'h2):(1'h1)] - (8'ha6)) : $signed((reg2142 ?
                      (reg1811 ? reg2149 : reg1941) : {(7'h55)}))));
              reg2148 = $signed($signed((reg2028 - reg1793)));
              reg2149 = reg1949[(3'h7):(3'h4)];
              reg2151 <= ($unsigned((reg1816[(4'he):(1'h0)] - ($unsigned((7'h50)) << wire1774[(3'h4):(2'h2)]))) ?
                  {({reg1933} ?
                          $unsigned((reg1814 != reg1948)) : ($unsigned(reg1971) || (reg1872 << reg2148)))} : (reg1816 | reg1858));
            end
          for (forvar2152 = (1'h0); (forvar2152 < (3'h4)); forvar2152 = (forvar2152 + (1'h1)))
            begin
              reg2153 = (reg2148[(2'h2):(1'h0)] ?
                  (-wire1774) : $unsigned($signed(reg2057)));
              reg2154 = {{reg2069[(2'h3):(1'h0)], reg1961[(3'h5):(2'h2)]},
                  ($signed({$signed(reg1988),
                          ((7'h42) ? reg1859 : reg1785),
                          reg2147}) ?
                      (!reg2052) : $unsigned(((wire1909 | reg1859) + $signed(reg2063)))),
                  (reg1880 ?
                      reg2134[(2'h3):(2'h2)] : $signed((!(reg1970 ?
                          (8'hb1) : reg1946))))};
              reg2155 <= ((|(reg1960[(1'h1):(1'h0)] <= wire1904[(4'hc):(1'h0)])) == reg2081[(3'h4):(2'h2)]);
              reg2156 <= wire1774;
              reg2157 = (reg2009[(4'ha):(3'h6)] ?
                  (reg2062 ^~ ($unsigned(((8'haa) ? reg1902 : reg1876)) ?
                      (^~(reg2130 ?
                          (8'hb7) : reg1799)) : (reg2000[(5'h11):(4'h9)] >>> $signed(reg1791)))) : reg1883);
              reg2158 <= (((((reg1978 ? reg1933 : reg1863) ?
                      $unsigned((7'h45)) : reg2021[(2'h3):(1'h1)]) ?
                  $signed(wire1775[(5'h1a):(2'h2)]) : ({reg1836} ?
                      (reg2044 ? reg1872 : reg2114) : {reg2030,
                          reg1970,
                          reg1944})) < ($signed((reg1857 >= (8'ha5))) ~^ (~&$unsigned(reg2038)))) ~^ $signed(($signed((reg1948 ?
                  reg1961 : reg1980)) ^ ($signed((7'h4b)) | reg1874))));
            end
        end
      for (forvar2159 = (1'h0); (forvar2159 < (2'h2)); forvar2159 = (forvar2159 + (1'h1)))
        begin
          if ($signed(reg1980))
            begin
              reg2160 = ($signed((|(^$unsigned(reg2149)))) ?
                  (((-$unsigned(reg1911)) || $unsigned($unsigned(wire1906))) * reg1908) : $unsigned({reg1932[(1'h1):(1'h0)]}));
              reg2161 = reg1988[(4'ha):(1'h1)];
            end
          else
            begin
              reg2160 = $signed($unsigned($unsigned({reg2156[(3'h4):(3'h4)]})));
              reg2162 <= reg1937[(5'h1d):(5'h16)];
            end
          reg2163 <= $signed($unsigned($unsigned($unsigned(reg2004[(5'h18):(4'he)]))));
          reg2164 <= (&($unsigned(($signed(wire2078) + (~&reg1800))) > (~(reg1993[(5'h17):(5'h15)] ?
              reg1872[(4'h8):(4'h8)] : $unsigned((7'h53))))));
        end
    end
  assign wire2165 = reg1840;
  always
    @(posedge clk) begin
      reg2166 = (8'ha8);
      reg2167 <= (reg1832[(3'h4):(1'h1)] ?
          reg1836[(4'h9):(3'h6)] : ({(~^$signed(reg1783)),
              (reg1811 ?
                  (-reg2162) : (reg2011 ?
                      reg1977 : reg1914))} == (reg1874 >= {{reg2049, reg1814},
              (reg2121 ? reg1927 : reg1927),
              reg1916})));
      reg2168 <= $signed(reg1818[(1'h0):(1'h0)]);
      for (forvar2169 = (1'h0); (forvar2169 < (1'h1)); forvar2169 = (forvar2169 + (1'h1)))
        begin
          for (forvar2170 = (1'h0); (forvar2170 < (3'h5)); forvar2170 = (forvar2170 + (1'h1)))
            begin
              reg2171 = reg1884[(2'h2):(2'h2)];
              reg2172 <= (^~$signed($signed(reg2030[(3'h5):(2'h2)])));
            end
          reg2173 <= reg2130[(5'h10):(5'h10)];
          reg2174 <= $unsigned(reg2028[(1'h1):(1'h1)]);
          reg2175 <= (reg1872[(1'h0):(1'h0)] << reg2103[(4'hb):(4'hb)]);
          for (forvar2176 = (1'h0); (forvar2176 < (3'h6)); forvar2176 = (forvar2176 + (1'h1)))
            begin
              reg2177 <= (reg2100 | reg2110);
              reg2178 = $signed({$unsigned((reg1857 != $unsigned(reg1959)))});
              reg2179 <= (((reg2178 ?
                  ((|reg1879) != (reg1931 * reg1959)) : ((~^reg2163) ?
                      $unsigned(reg1811) : reg1785[(3'h4):(2'h2)])) & wire2006[(1'h1):(1'h0)]) == (&(reg2031 + $signed((8'ha7)))));
            end
          reg2180 <= $signed($unsigned(reg2173));
          for (forvar2181 = (1'h0); (forvar2181 < (3'h6)); forvar2181 = (forvar2181 + (1'h1)))
            begin
              reg2182 <= $unsigned((reg2088 > ({$signed(reg2172)} ?
                  ($unsigned((7'h45)) + (reg2057 ?
                      reg2114 : reg1865)) : reg1836[(3'h6):(3'h5)])));
              reg2183 <= reg2114;
              reg2184 = ({$signed({reg2141[(3'h5):(3'h5)],
                          ((8'hb3) - (8'hb8))}),
                      $unsigned($unsigned(reg2052))} ?
                  reg2151 : reg2096[(4'h8):(3'h7)]);
              reg2185 = ((+((!((7'h53) ?
                      reg2047 : reg2168)) | {$signed(reg1937),
                      (reg1966 ? reg1782 : reg2162)})) ?
                  $signed((+reg2058)) : ({$signed($unsigned(reg2127)),
                      ((reg1824 >> reg2028) != $signed(reg2171))} - $signed(reg1917[(5'h11):(5'h11)])));
              reg2186 = {reg2009[(3'h4):(1'h0)],
                  $signed({$unsigned((reg2097 ? reg2069 : reg2147))}),
                  (reg2085 ? reg1814 : reg1955)};
            end
        end
      reg2187 <= $signed(((($unsigned(reg2100) ?
                  reg1937 : (reg1997 ? wire2059 : reg1797)) ?
              (8'ha3) : ((~|reg1990) - {reg1883})) ?
          reg2021 : reg2044));
      if ($unsigned((~&reg2158[(1'h0):(1'h0)])))
        begin
          reg2188 = {(($signed({(8'hb4), reg2063, reg1811}) ?
                      (&reg1970[(4'hc):(4'hc)]) : reg2146[(3'h5):(2'h2)]) ?
                  (((wire1775 <<< reg2030) >>> reg1916) ?
                      (reg2180[(5'h17):(1'h0)] ?
                          $signed(reg2004) : (8'hb6)) : reg1873) : (({reg2127} ?
                      ((7'h43) ?
                          reg1980 : reg2139) : reg2132[(4'h8):(1'h1)]) == ($signed(reg2182) ?
                      (!reg1880) : wire1909[(5'h10):(3'h4)]))),
              $unsigned({reg2166[(3'h7):(2'h3)],
                  ($unsigned(reg2100) ?
                      $unsigned(wire2165) : (reg1896 > (8'ha8)))})};
          reg2189 <= (8'hac);
          for (forvar2190 = (1'h0); (forvar2190 < (1'h0)); forvar2190 = (forvar2190 + (1'h1)))
            begin
              reg2191 = $signed($unsigned(reg2096));
              reg2192 <= $unsigned($unsigned($unsigned(({reg1891,
                      reg1951,
                      reg1961} ?
                  (reg2010 + (8'hbd)) : $unsigned(reg2147)))));
              reg2193 <= $signed(($signed(reg1971[(3'h5):(1'h1)]) < reg1814));
              reg2194 <= reg2121[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg2188 = {{reg2194},
              $unsigned(((8'hab) ?
                  {(~&reg2030),
                      reg1811,
                      (reg1877 ? reg2021 : reg1797)} : reg2069[(4'hb):(3'h7)])),
              (+(~|(~^{reg1965})))};
          reg2189 <= $signed(((reg2177[(4'hc):(3'h5)] - {$signed(reg2022),
                  {wire2059},
                  $unsigned(reg2139)}) ?
              (reg1947[(4'ha):(3'h5)] * ($signed(reg1977) < (reg1945 && reg2179))) : reg2155[(5'h1d):(4'he)]));
          for (forvar2190 = (1'h0); (forvar2190 < (3'h5)); forvar2190 = (forvar2190 + (1'h1)))
            begin
              reg2192 <= $unsigned({$signed(wire1774[(4'h8):(2'h2)]), reg1807});
            end
          reg2193 <= reg2121[(4'he):(2'h2)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1376
#(parameter param1769 = (~(~|((8'hb7) ? (+(~^(8'hbd))) : ((|(8'had)) ? {(7'h4d), (8'hb7)} : ((7'h50) * (8'hbf)))))))
(y, clk, wire1381, wire1380, wire1379, wire1378, wire1377);
  output wire [(32'h1a96):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire1381;
  input wire signed [(5'h13):(1'h0)] wire1380;
  input wire [(5'h1f):(1'h0)] wire1379;
  input wire signed [(4'ha):(1'h0)] wire1378;
  input wire signed [(4'hf):(1'h0)] wire1377;
  wire signed [(4'hf):(1'h0)] wire1764;
  wire [(5'h18):(1'h0)] wire1763;
  wire [(5'h1a):(1'h0)] wire1762;
  wire [(5'h17):(1'h0)] wire1761;
  wire [(4'hd):(1'h0)] wire1760;
  wire signed [(4'hb):(1'h0)] wire1669;
  wire signed [(3'h7):(1'h0)] wire1668;
  wire [(5'h11):(1'h0)] wire1648;
  wire [(4'hb):(1'h0)] wire1647;
  wire [(5'h1d):(1'h0)] wire1585;
  wire [(4'hf):(1'h0)] wire1584;
  wire [(5'h1a):(1'h0)] wire1583;
  wire [(5'h1a):(1'h0)] wire1567;
  wire [(5'h1b):(1'h0)] wire1566;
  wire signed [(2'h2):(1'h0)] wire1462;
  wire [(5'h1a):(1'h0)] wire1461;
  wire signed [(3'h4):(1'h0)] wire1460;
  wire signed [(5'h12):(1'h0)] wire1422;
  reg signed [(2'h2):(1'h0)] reg1766 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1759 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1758 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1755 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1752 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1748 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1747 = (1'h0);
  reg [(5'h17):(1'h0)] reg1746 = (1'h0);
  reg [(3'h4):(1'h0)] reg1744 = (1'h0);
  reg [(3'h5):(1'h0)] reg1743 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1742 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1740 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1739 = (1'h0);
  reg [(3'h5):(1'h0)] reg1734 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1733 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1732 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1730 = (1'h0);
  reg [(5'h18):(1'h0)] reg1726 = (1'h0);
  reg [(3'h7):(1'h0)] reg1721 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1720 = (1'h0);
  reg [(5'h12):(1'h0)] reg1719 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1717 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1716 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1715 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1714 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1713 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1712 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1711 = (1'h0);
  reg [(5'h19):(1'h0)] reg1710 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1709 = (1'h0);
  reg [(5'h12):(1'h0)] reg1708 = (1'h0);
  reg [(5'h14):(1'h0)] reg1705 = (1'h0);
  reg [(4'hd):(1'h0)] reg1704 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1702 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1700 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1698 = (1'h0);
  reg [(2'h3):(1'h0)] reg1697 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1695 = (1'h0);
  reg [(4'ha):(1'h0)] reg1690 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1689 = (1'h0);
  reg [(5'h18):(1'h0)] reg1688 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1687 = (1'h0);
  reg [(3'h7):(1'h0)] reg1685 = (1'h0);
  reg [(5'h15):(1'h0)] reg1683 = (1'h0);
  reg [(5'h15):(1'h0)] reg1682 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1681 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1678 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1673 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1671 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1670 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1663 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1662 = (1'h0);
  reg [(3'h7):(1'h0)] reg1661 = (1'h0);
  reg [(5'h15):(1'h0)] reg1660 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1658 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1652 = (1'h0);
  reg [(4'h8):(1'h0)] reg1650 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1645 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1644 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1622 = (1'h0);
  reg [(5'h11):(1'h0)] reg1643 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1642 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1641 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1639 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1637 = (1'h0);
  reg [(5'h11):(1'h0)] reg1633 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1631 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1630 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1626 = (1'h0);
  reg [(4'hc):(1'h0)] reg1625 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1624 = (1'h0);
  reg [(5'h14):(1'h0)] reg1623 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1619 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1617 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1614 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1613 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1611 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1608 = (1'h0);
  reg [(4'hc):(1'h0)] reg1607 = (1'h0);
  reg [(5'h12):(1'h0)] reg1606 = (1'h0);
  reg [(4'he):(1'h0)] reg1604 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1601 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1600 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1599 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1598 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1595 = (1'h0);
  reg [(5'h12):(1'h0)] reg1593 = (1'h0);
  reg [(4'h8):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1591 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1590 = (1'h0);
  reg [(5'h12):(1'h0)] reg1589 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1588 = (1'h0);
  reg [(5'h19):(1'h0)] reg1582 = (1'h0);
  reg [(3'h5):(1'h0)] reg1581 = (1'h0);
  reg [(2'h3):(1'h0)] reg1577 = (1'h0);
  reg [(5'h19):(1'h0)] reg1576 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1575 = (1'h0);
  reg [(4'ha):(1'h0)] reg1573 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1572 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1568 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1565 = (1'h0);
  reg [(4'he):(1'h0)] reg1564 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1563 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1561 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1560 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1559 = (1'h0);
  reg [(2'h3):(1'h0)] reg1556 = (1'h0);
  reg [(5'h16):(1'h0)] reg1553 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1552 = (1'h0);
  reg [(5'h11):(1'h0)] reg1550 = (1'h0);
  reg [(5'h18):(1'h0)] reg1544 = (1'h0);
  reg [(3'h6):(1'h0)] reg1547 = (1'h0);
  reg [(5'h12):(1'h0)] reg1546 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1545 = (1'h0);
  reg [(5'h14):(1'h0)] reg1534 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1531 = (1'h0);
  reg [(4'hb):(1'h0)] reg1529 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1528 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1525 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1524 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1521 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1520 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1516 = (1'h0);
  reg [(4'hd):(1'h0)] reg1515 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1514 = (1'h0);
  reg [(4'ha):(1'h0)] reg1512 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1507 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1502 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1510 = (1'h0);
  reg [(5'h18):(1'h0)] reg1509 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1508 = (1'h0);
  reg [(3'h7):(1'h0)] reg1505 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1504 = (1'h0);
  reg [(3'h4):(1'h0)] reg1501 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1500 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1497 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1496 = (1'h0);
  reg [(4'he):(1'h0)] reg1493 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1491 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1489 = (1'h0);
  reg [(4'hd):(1'h0)] reg1487 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1486 = (1'h0);
  reg [(5'h15):(1'h0)] reg1485 = (1'h0);
  reg [(4'he):(1'h0)] reg1483 = (1'h0);
  reg [(3'h7):(1'h0)] reg1481 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1479 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1478 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1474 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1473 = (1'h0);
  reg [(2'h2):(1'h0)] reg1472 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1470 = (1'h0);
  reg [(3'h6):(1'h0)] reg1467 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1465 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1464 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1463 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1458 = (1'h0);
  reg [(3'h4):(1'h0)] reg1456 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1454 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1453 = (1'h0);
  reg [(4'h8):(1'h0)] reg1452 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1451 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1447 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1446 = (1'h0);
  reg [(5'h11):(1'h0)] reg1445 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1444 = (1'h0);
  reg [(4'hd):(1'h0)] reg1441 = (1'h0);
  reg [(3'h4):(1'h0)] reg1425 = (1'h0);
  reg [(3'h5):(1'h0)] reg1440 = (1'h0);
  reg [(5'h16):(1'h0)] reg1439 = (1'h0);
  reg [(5'h12):(1'h0)] reg1436 = (1'h0);
  reg [(5'h14):(1'h0)] reg1435 = (1'h0);
  reg [(5'h16):(1'h0)] reg1432 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1431 = (1'h0);
  reg [(4'h9):(1'h0)] reg1430 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1428 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1427 = (1'h0);
  reg [(5'h18):(1'h0)] reg1426 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1415 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1414 = (1'h0);
  reg [(4'h9):(1'h0)] reg1412 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1411 = (1'h0);
  reg [(4'hf):(1'h0)] reg1406 = (1'h0);
  reg [(5'h10):(1'h0)] reg1397 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1393 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1391 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1388 = (1'h0);
  reg [(5'h10):(1'h0)] reg1386 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1385 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1768 = (1'h0);
  reg [(5'h14):(1'h0)] reg1767 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1765 = (1'h0);
  reg [(4'ha):(1'h0)] reg1757 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1756 = (1'h0);
  reg [(5'h14):(1'h0)] reg1754 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1753 = (1'h0);
  reg [(4'hb):(1'h0)] reg1751 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1750 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1749 = (1'h0);
  reg [(3'h5):(1'h0)] reg1745 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1741 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1738 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1737 = (1'h0);
  reg [(5'h11):(1'h0)] reg1736 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1735 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1731 = (1'h0);
  reg [(3'h5):(1'h0)] reg1729 = (1'h0);
  reg [(5'h12):(1'h0)] reg1728 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1727 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1725 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1724 = (1'h0);
  reg [(3'h4):(1'h0)] reg1723 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1722 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1718 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1707 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1706 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1693 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1692 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1703 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1701 = (1'h0);
  reg [(3'h7):(1'h0)] reg1699 = (1'h0);
  reg [(4'hd):(1'h0)] reg1696 = (1'h0);
  reg [(5'h13):(1'h0)] reg1694 = (1'h0);
  reg [(2'h2):(1'h0)] reg1693 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1692 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1691 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1686 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1684 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1680 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1679 = (1'h0);
  reg [(4'hd):(1'h0)] reg1677 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1676 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1675 = (1'h0);
  reg [(3'h6):(1'h0)] reg1674 = (1'h0);
  reg [(4'h8):(1'h0)] reg1672 = (1'h0);
  reg [(4'hd):(1'h0)] reg1667 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1666 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1665 = (1'h0);
  reg [(4'h8):(1'h0)] reg1664 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1659 = (1'h0);
  reg [(5'h11):(1'h0)] reg1657 = (1'h0);
  reg [(5'h19):(1'h0)] reg1656 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1655 = (1'h0);
  reg [(4'ha):(1'h0)] reg1654 = (1'h0);
  reg [(5'h11):(1'h0)] reg1653 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1651 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1649 = (1'h0);
  reg [(5'h17):(1'h0)] reg1646 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1640 = (1'h0);
  reg [(4'he):(1'h0)] forvar1638 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1636 = (1'h0);
  reg [(4'ha):(1'h0)] reg1635 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1634 = (1'h0);
  reg [(4'hd):(1'h0)] reg1632 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1629 = (1'h0);
  reg [(2'h3):(1'h0)] reg1628 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1627 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1622 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1621 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1602 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1620 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1618 = (1'h0);
  reg [(5'h15):(1'h0)] reg1616 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1615 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1612 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1610 = (1'h0);
  reg [(5'h15):(1'h0)] reg1609 = (1'h0);
  reg [(4'ha):(1'h0)] reg1605 = (1'h0);
  reg [(4'hc):(1'h0)] reg1603 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1602 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1597 = (1'h0);
  reg [(4'ha):(1'h0)] reg1596 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1594 = (1'h0);
  reg [(3'h4):(1'h0)] reg1587 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1586 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1580 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1579 = (1'h0);
  reg [(5'h17):(1'h0)] reg1578 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1574 = (1'h0);
  reg [(5'h18):(1'h0)] reg1571 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1570 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1569 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1562 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1558 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1557 = (1'h0);
  reg [(5'h15):(1'h0)] reg1555 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1554 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1551 = (1'h0);
  reg [(2'h2):(1'h0)] reg1549 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1548 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1544 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1543 = (1'h0);
  reg [(5'h15):(1'h0)] reg1542 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1541 = (1'h0);
  reg [(5'h19):(1'h0)] reg1540 = (1'h0);
  reg [(4'ha):(1'h0)] reg1539 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1538 = (1'h0);
  reg [(5'h16):(1'h0)] reg1537 = (1'h0);
  reg [(4'hf):(1'h0)] reg1536 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1535 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1533 = (1'h0);
  reg [(4'ha):(1'h0)] reg1532 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1523 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1522 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1519 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1530 = (1'h0);
  reg [(2'h3):(1'h0)] reg1527 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1526 = (1'h0);
  reg [(4'hb):(1'h0)] reg1523 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1522 = (1'h0);
  reg [(5'h12):(1'h0)] reg1519 = (1'h0);
  reg [(4'hb):(1'h0)] reg1518 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1517 = (1'h0);
  reg [(5'h13):(1'h0)] reg1513 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1511 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1507 = (1'h0);
  reg [(4'hf):(1'h0)] reg1506 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1503 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1502 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1499 = (1'h0);
  reg [(4'hc):(1'h0)] reg1498 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1495 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1494 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1492 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1490 = (1'h0);
  reg [(5'h12):(1'h0)] reg1488 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1488 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1484 = (1'h0);
  reg [(4'h9):(1'h0)] reg1482 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1480 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1477 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1476 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1475 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1471 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1469 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1468 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1466 = (1'h0);
  reg [(4'he):(1'h0)] reg1459 = (1'h0);
  reg [(3'h7):(1'h0)] reg1457 = (1'h0);
  reg [(5'h16):(1'h0)] reg1455 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1450 = (1'h0);
  reg [(4'ha):(1'h0)] reg1449 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1448 = (1'h0);
  reg [(4'hd):(1'h0)] reg1443 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1442 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1438 = (1'h0);
  reg [(4'ha):(1'h0)] reg1437 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1434 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1433 = (1'h0);
  reg [(4'hb):(1'h0)] reg1429 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1425 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1424 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1423 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1421 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1420 = (1'h0);
  reg [(5'h17):(1'h0)] reg1419 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1418 = (1'h0);
  reg [(4'hb):(1'h0)] reg1417 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1416 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1413 = (1'h0);
  reg [(3'h4):(1'h0)] reg1410 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1409 = (1'h0);
  reg [(5'h10):(1'h0)] reg1408 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1407 = (1'h0);
  reg [(3'h6):(1'h0)] reg1405 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1404 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1403 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1402 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1401 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1400 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1399 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1398 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1396 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1395 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1394 = (1'h0);
  reg [(5'h14):(1'h0)] reg1392 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1390 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1389 = (1'h0);
  reg [(4'hd):(1'h0)] reg1387 = (1'h0);
  reg [(5'h19):(1'h0)] reg1384 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1383 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1382 = (1'h0);
  assign y = {wire1764,
                 wire1763,
                 wire1762,
                 wire1761,
                 wire1760,
                 wire1669,
                 wire1668,
                 wire1648,
                 wire1647,
                 wire1585,
                 wire1584,
                 wire1583,
                 wire1567,
                 wire1566,
                 wire1462,
                 wire1461,
                 wire1460,
                 wire1422,
                 reg1766,
                 reg1759,
                 reg1758,
                 reg1755,
                 reg1752,
                 reg1748,
                 reg1747,
                 reg1746,
                 reg1744,
                 reg1743,
                 reg1742,
                 reg1740,
                 reg1739,
                 reg1734,
                 reg1733,
                 reg1732,
                 reg1730,
                 reg1726,
                 reg1721,
                 reg1720,
                 reg1719,
                 reg1717,
                 reg1716,
                 reg1715,
                 reg1714,
                 reg1713,
                 reg1712,
                 reg1711,
                 reg1710,
                 reg1709,
                 reg1708,
                 reg1705,
                 reg1704,
                 reg1702,
                 reg1700,
                 reg1698,
                 reg1697,
                 reg1695,
                 reg1690,
                 reg1689,
                 reg1688,
                 reg1687,
                 reg1685,
                 reg1683,
                 reg1682,
                 reg1681,
                 reg1678,
                 reg1673,
                 reg1671,
                 reg1670,
                 reg1663,
                 reg1662,
                 reg1661,
                 reg1660,
                 reg1658,
                 reg1652,
                 reg1650,
                 reg1645,
                 reg1644,
                 reg1622,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1639,
                 reg1637,
                 reg1633,
                 reg1631,
                 reg1630,
                 reg1626,
                 reg1625,
                 reg1624,
                 reg1623,
                 reg1619,
                 reg1617,
                 reg1614,
                 reg1613,
                 reg1611,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1604,
                 reg1601,
                 reg1600,
                 reg1599,
                 reg1598,
                 reg1595,
                 reg1593,
                 reg1592,
                 reg1591,
                 reg1590,
                 reg1589,
                 reg1588,
                 reg1582,
                 reg1581,
                 reg1577,
                 reg1576,
                 reg1575,
                 reg1573,
                 reg1572,
                 reg1568,
                 reg1565,
                 reg1564,
                 reg1563,
                 reg1561,
                 reg1560,
                 reg1559,
                 reg1556,
                 reg1553,
                 reg1552,
                 reg1550,
                 reg1544,
                 reg1547,
                 reg1546,
                 reg1545,
                 reg1534,
                 reg1531,
                 reg1529,
                 reg1528,
                 reg1525,
                 reg1524,
                 reg1521,
                 reg1520,
                 reg1516,
                 reg1515,
                 reg1514,
                 reg1512,
                 reg1507,
                 reg1502,
                 reg1510,
                 reg1509,
                 reg1508,
                 reg1505,
                 reg1504,
                 reg1501,
                 reg1500,
                 reg1497,
                 reg1496,
                 reg1493,
                 reg1491,
                 reg1489,
                 reg1487,
                 reg1486,
                 reg1485,
                 reg1483,
                 reg1481,
                 reg1479,
                 reg1478,
                 reg1474,
                 reg1473,
                 reg1472,
                 reg1470,
                 reg1467,
                 reg1465,
                 reg1464,
                 reg1463,
                 reg1458,
                 reg1456,
                 reg1454,
                 reg1453,
                 reg1452,
                 reg1451,
                 reg1447,
                 reg1446,
                 reg1445,
                 reg1444,
                 reg1441,
                 reg1425,
                 reg1440,
                 reg1439,
                 reg1436,
                 reg1435,
                 reg1432,
                 reg1431,
                 reg1430,
                 reg1428,
                 reg1427,
                 reg1426,
                 reg1415,
                 reg1414,
                 reg1412,
                 reg1411,
                 reg1406,
                 reg1397,
                 reg1393,
                 reg1391,
                 reg1388,
                 reg1386,
                 reg1385,
                 reg1768,
                 reg1767,
                 forvar1765,
                 reg1757,
                 reg1756,
                 reg1754,
                 forvar1753,
                 reg1751,
                 forvar1750,
                 reg1749,
                 reg1745,
                 forvar1741,
                 reg1738,
                 reg1737,
                 reg1736,
                 forvar1735,
                 reg1731,
                 reg1729,
                 reg1728,
                 forvar1727,
                 reg1725,
                 forvar1724,
                 reg1723,
                 reg1722,
                 reg1718,
                 forvar1707,
                 forvar1706,
                 forvar1693,
                 reg1692,
                 reg1703,
                 forvar1701,
                 reg1699,
                 reg1696,
                 reg1694,
                 reg1693,
                 forvar1692,
                 reg1691,
                 reg1686,
                 reg1684,
                 reg1680,
                 reg1679,
                 reg1677,
                 reg1676,
                 reg1675,
                 reg1674,
                 reg1672,
                 reg1667,
                 reg1666,
                 reg1665,
                 reg1664,
                 reg1659,
                 reg1657,
                 reg1656,
                 reg1655,
                 reg1654,
                 reg1653,
                 reg1651,
                 reg1649,
                 reg1646,
                 reg1640,
                 forvar1638,
                 forvar1636,
                 reg1635,
                 reg1634,
                 reg1632,
                 reg1629,
                 reg1628,
                 reg1627,
                 forvar1622,
                 reg1621,
                 reg1602,
                 reg1620,
                 forvar1618,
                 reg1616,
                 reg1615,
                 reg1612,
                 reg1610,
                 reg1609,
                 reg1605,
                 reg1603,
                 forvar1602,
                 reg1597,
                 reg1596,
                 reg1594,
                 reg1587,
                 forvar1586,
                 reg1580,
                 reg1579,
                 reg1578,
                 reg1574,
                 reg1571,
                 reg1570,
                 forvar1569,
                 reg1562,
                 forvar1558,
                 reg1557,
                 reg1555,
                 reg1554,
                 reg1551,
                 reg1549,
                 reg1548,
                 forvar1544,
                 reg1543,
                 reg1542,
                 reg1541,
                 reg1540,
                 reg1539,
                 reg1538,
                 reg1537,
                 reg1536,
                 reg1535,
                 forvar1533,
                 reg1532,
                 forvar1523,
                 reg1522,
                 forvar1519,
                 reg1530,
                 reg1527,
                 reg1526,
                 reg1523,
                 forvar1522,
                 reg1519,
                 reg1518,
                 reg1517,
                 reg1513,
                 forvar1511,
                 forvar1507,
                 reg1506,
                 reg1503,
                 forvar1502,
                 forvar1499,
                 reg1498,
                 forvar1495,
                 reg1494,
                 reg1492,
                 reg1490,
                 reg1488,
                 forvar1488,
                 reg1484,
                 reg1482,
                 reg1480,
                 reg1477,
                 forvar1476,
                 reg1475,
                 reg1471,
                 reg1469,
                 forvar1468,
                 reg1466,
                 reg1459,
                 reg1457,
                 reg1455,
                 forvar1450,
                 reg1449,
                 forvar1448,
                 reg1443,
                 reg1442,
                 reg1438,
                 reg1437,
                 reg1434,
                 reg1433,
                 reg1429,
                 forvar1425,
                 reg1424,
                 reg1423,
                 reg1421,
                 reg1420,
                 reg1419,
                 reg1418,
                 reg1417,
                 reg1416,
                 reg1413,
                 reg1410,
                 reg1409,
                 reg1408,
                 reg1407,
                 reg1405,
                 reg1404,
                 forvar1403,
                 reg1402,
                 forvar1401,
                 reg1400,
                 reg1399,
                 reg1398,
                 reg1396,
                 forvar1395,
                 reg1394,
                 reg1392,
                 reg1390,
                 reg1389,
                 reg1387,
                 reg1384,
                 reg1383,
                 forvar1382,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned(($unsigned($unsigned(((8'hae) == wire1377))) ?
          $unsigned($signed($unsigned(wire1378))) : ($signed({wire1381}) <<< (-(wire1378 ?
              wire1381 : (8'hbf)))))))
        begin
          for (forvar1382 = (1'h0); (forvar1382 < (3'h4)); forvar1382 = (forvar1382 + (1'h1)))
            begin
              reg1383 = $signed((!((wire1377 ?
                  {wire1377} : wire1379) > wire1378[(4'h8):(3'h5)])));
            end
        end
      else
        begin
          for (forvar1382 = (1'h0); (forvar1382 < (3'h5)); forvar1382 = (forvar1382 + (1'h1)))
            begin
              reg1383 = ((({$signed(wire1379),
                              (wire1381 ~^ wire1379),
                              {wire1378, (7'h4e), (8'had)}} ?
                          ((wire1380 != wire1380) * (wire1377 > (7'h57))) : ($signed(wire1379) ?
                              $unsigned(wire1378) : (wire1380 ?
                                  wire1381 : forvar1382))) ?
                      (-reg1383) : ((|(wire1381 <<< wire1378)) ?
                          wire1377[(4'he):(4'hc)] : wire1377)) ?
                  (^wire1377[(4'hb):(4'ha)]) : wire1381[(3'h6):(3'h6)]);
              reg1384 = ((-wire1378[(1'h1):(1'h0)]) ?
                  reg1383[(3'h7):(2'h3)] : forvar1382);
              reg1385 <= ((wire1381 >>> ($unsigned((wire1380 - wire1377)) ?
                      forvar1382[(4'h9):(2'h2)] : ($unsigned(forvar1382) ?
                          $signed((8'ha2)) : $unsigned(wire1380)))) ?
                  $unsigned(($signed((~|(7'h40))) != $unsigned($unsigned(wire1379)))) : {(wire1378[(4'h9):(2'h3)] != (8'hbf))});
            end
          if ((^~(({$unsigned(wire1378)} - (7'h40)) == ((wire1380 > {(7'h47)}) & ((forvar1382 && wire1378) ?
              wire1378[(1'h0):(1'h0)] : wire1380)))))
            begin
              reg1386 <= $signed((wire1380[(4'ha):(3'h6)] ?
                  ({wire1377,
                      $unsigned(reg1385),
                      (wire1379 * (8'hbc))} >= ((~&wire1381) ^~ $signed(reg1384))) : ($signed($unsigned(wire1380)) ?
                      $unsigned({forvar1382}) : $signed((wire1379 | wire1380)))));
              reg1387 = $unsigned(reg1384);
              reg1388 <= $signed((wire1377[(4'hd):(4'h8)] >= (&(~$signed(reg1383)))));
              reg1389 = ($unsigned(wire1379[(5'h18):(4'hc)]) ^~ (&$unsigned($unsigned($signed(reg1387)))));
              reg1390 = (forvar1382[(4'hd):(4'h8)] ?
                  $unsigned({$signed($unsigned(reg1384))}) : (~&$unsigned($unsigned(forvar1382))));
              reg1391 <= $signed(({reg1383[(5'h12):(5'h12)],
                      wire1377[(4'h9):(4'h8)],
                      $unsigned((reg1384 >> wire1378))} ?
                  wire1381[(1'h0):(1'h0)] : (wire1379 ?
                      wire1379[(5'h11):(4'hf)] : $unsigned(wire1381[(1'h0):(1'h0)]))));
              reg1392 = {(wire1381 < {(+(reg1389 << (7'h4f))), (~reg1389)}),
                  ((^{reg1387[(3'h6):(3'h6)]}) | $signed(($unsigned(wire1377) >>> $signed((8'hba))))),
                  ($signed(reg1383) ?
                      (((reg1386 ~^ reg1387) >= ((7'h50) ?
                              reg1390 : forvar1382)) ?
                          (wire1377 && (reg1388 ?
                              (7'h46) : wire1379)) : $unsigned($signed(reg1385))) : $signed((reg1383[(3'h4):(3'h4)] ?
                          (-wire1377) : (reg1387 ? reg1391 : reg1386))))};
            end
          else
            begin
              reg1386 <= $unsigned((wire1381 | $unsigned(reg1387[(4'h9):(1'h0)])));
              reg1387 = ((~^{(wire1381 ? reg1389 : reg1383[(5'h12):(3'h6)]),
                  $unsigned(reg1383)}) ^~ (&(~|$signed($signed(reg1390)))));
              reg1388 <= $unsigned(($unsigned(((reg1386 ? reg1391 : reg1384) ?
                      reg1391[(3'h6):(3'h5)] : reg1387)) ?
                  (~wire1381[(3'h5):(3'h4)]) : reg1383[(1'h1):(1'h0)]));
              reg1391 <= (+(8'had));
              reg1393 <= (~(~^(&wire1377[(2'h2):(1'h1)])));
              reg1394 = $signed($signed(reg1387[(4'hc):(1'h1)]));
            end
          for (forvar1395 = (1'h0); (forvar1395 < (1'h1)); forvar1395 = (forvar1395 + (1'h1)))
            begin
              reg1396 = (((|{(^reg1389), (wire1379 + reg1384)}) ?
                      ($unsigned((reg1391 ? reg1391 : reg1388)) ?
                          {(reg1387 ^ reg1394),
                              $unsigned(wire1378),
                              (-forvar1395)} : (~^reg1383[(3'h4):(3'h4)])) : $signed(($signed(wire1378) ?
                          $unsigned(wire1381) : {reg1390, (8'hb7), reg1389}))) ?
                  {(~&$signed($signed((7'h57))))} : (($unsigned({reg1385,
                      (7'h47)}) == $unsigned($signed(reg1393))) ~^ (!wire1377)));
            end
          reg1397 <= $signed((wire1377[(2'h3):(2'h3)] ?
              reg1396 : $signed((7'h46))));
          reg1398 = (^~(8'hae));
          reg1399 = reg1390[(3'h6):(3'h6)];
          reg1400 = (~|reg1390);
        end
      for (forvar1401 = (1'h0); (forvar1401 < (2'h2)); forvar1401 = (forvar1401 + (1'h1)))
        begin
          reg1402 = $unsigned(reg1393[(2'h3):(2'h2)]);
          for (forvar1403 = (1'h0); (forvar1403 < (1'h1)); forvar1403 = (forvar1403 + (1'h1)))
            begin
              reg1404 = reg1393[(1'h0):(1'h0)];
              reg1405 = reg1400;
              reg1406 <= ((^~((^(reg1400 ?
                      reg1391 : wire1380)) & {$signed(forvar1403)})) ?
                  reg1389[(4'h9):(2'h2)] : $signed($unsigned(($signed(reg1404) ?
                      ((8'ha3) - reg1400) : $signed((8'ha9))))));
              reg1407 = reg1390;
              reg1408 = ((!(~&{(~^(8'had)),
                  ((8'hb5) ? reg1394 : (8'hb8)),
                  $signed((7'h56))})) & (reg1407[(5'h14):(4'h8)] ?
                  forvar1382[(3'h5):(1'h1)] : (-wire1380[(4'ha):(3'h7)])));
            end
          reg1409 = forvar1401[(5'h1c):(5'h13)];
          if ($unsigned($unsigned(($signed(reg1406[(2'h2):(1'h0)]) >>> $signed($signed(reg1387))))))
            begin
              reg1410 = ((~|(reg1397 == $unsigned((reg1406 ?
                      reg1409 : wire1378)))) ?
                  wire1378 : {wire1379[(1'h0):(1'h0)], (reg1409 ^ (7'h56))});
              reg1411 <= ((reg1409 ?
                      (((reg1407 ^~ reg1397) ?
                          (reg1409 ?
                              reg1410 : reg1383) : {forvar1382}) <= ((reg1391 - reg1404) ?
                          reg1394 : (reg1408 - forvar1382))) : (wire1378 ?
                          $signed((reg1396 ? reg1410 : wire1378)) : ((reg1397 ?
                              (7'h4b) : wire1381) << (wire1381 ?
                              reg1391 : (7'h57))))) ?
                  reg1408 : ($unsigned((~^{wire1379, forvar1401, forvar1382})) ?
                      reg1386[(4'hc):(3'h7)] : (-(reg1404 != $signed(forvar1403)))));
              reg1412 <= (forvar1401[(5'h1d):(2'h2)] ?
                  reg1405[(1'h1):(1'h1)] : (^~(!reg1392[(3'h5):(2'h2)])));
              reg1413 = $unsigned($unsigned($signed(((reg1412 ?
                      (7'h44) : reg1383) ?
                  (^reg1398) : (wire1381 > wire1377)))));
              reg1414 <= $signed(reg1385);
              reg1415 <= (reg1393 ?
                  (7'h49) : ($signed($signed({reg1390, (8'hb5), reg1383})) ?
                      (7'h40) : $unsigned(reg1399)));
            end
          else
            begin
              reg1411 <= reg1386;
              reg1413 = (reg1391[(1'h1):(1'h1)] ?
                  ((reg1390 ?
                      reg1404 : reg1396) - reg1394[(1'h0):(1'h0)]) : $signed((wire1381 ?
                      reg1404 : reg1388[(3'h4):(1'h0)])));
              reg1416 = $signed(($unsigned((~^$unsigned(reg1393))) != (reg1411 ^~ {reg1404})));
              reg1417 = forvar1401;
              reg1418 = {reg1400,
                  (~|(({reg1391, forvar1403, (7'h58)} ?
                          (reg1396 ~^ reg1392) : $unsigned(reg1396)) ?
                      $signed(reg1387[(4'h8):(3'h6)]) : (^reg1384))),
                  reg1390[(2'h2):(1'h1)]};
              reg1419 = (+forvar1401[(5'h1a):(5'h13)]);
            end
          reg1420 = $signed($signed((8'haf)));
        end
      reg1421 = $unsigned($signed($unsigned(($unsigned(forvar1401) - (reg1419 ?
          reg1408 : reg1411)))));
    end
  assign wire1422 = wire1380;
  always
    @(posedge clk) begin
      reg1423 = wire1378[(3'h7):(3'h5)];
      reg1424 = $signed((-wire1422));
      if ((reg1393 + (~|({(reg1414 ^ wire1381)} && (~^$unsigned(reg1423))))))
        begin
          for (forvar1425 = (1'h0); (forvar1425 < (1'h1)); forvar1425 = (forvar1425 + (1'h1)))
            begin
              reg1426 <= ((~|$signed(($signed(reg1412) ~^ (reg1385 ~^ reg1397)))) | $signed((wire1422 ?
                  reg1391[(2'h2):(1'h1)] : forvar1425[(4'h8):(2'h3)])));
              reg1427 <= wire1378[(1'h1):(1'h1)];
              reg1428 <= $signed(reg1397);
              reg1429 = ({reg1427[(5'h15):(3'h4)],
                  ($unsigned((^~reg1424)) ? wire1422 : (!$signed(wire1422))),
                  $signed($unsigned($signed((8'hab))))} >= (reg1426[(5'h18):(5'h15)] >>> (^$unsigned((reg1428 ^~ reg1428)))));
              reg1430 <= (reg1393[(4'he):(3'h7)] ? (8'hab) : (-(~wire1380)));
              reg1431 <= $unsigned($signed({reg1423}));
            end
          if (wire1377)
            begin
              reg1432 <= (~reg1430);
              reg1433 = (~(8'ha8));
            end
          else
            begin
              reg1433 = ($signed($signed($unsigned($unsigned(reg1424)))) ?
                  (+$unsigned(((&reg1427) ?
                      ((8'ha4) ? reg1429 : (8'ha3)) : (reg1414 ?
                          reg1428 : reg1406)))) : $unsigned(($unsigned($unsigned(reg1423)) >>> (wire1377[(3'h6):(1'h0)] & ((7'h45) & reg1388)))));
              reg1434 = reg1414;
              reg1435 <= wire1380;
              reg1436 <= $signed(((($unsigned(wire1380) != $signed(wire1378)) >= ((+reg1424) != $unsigned(reg1435))) ^ $unsigned(reg1432)));
              reg1437 = {{$unsigned($signed((~^reg1385)))}};
              reg1438 = reg1385[(4'hb):(3'h4)];
              reg1439 <= $signed($signed((reg1437 | reg1412[(4'h8):(3'h7)])));
            end
          reg1440 <= (reg1385 & reg1428[(5'h13):(1'h1)]);
        end
      else
        begin
          if ({$unsigned((^~((reg1414 ~^ (8'hb0)) <= reg1415[(1'h0):(1'h0)])))})
            begin
              reg1425 <= reg1437[(2'h2):(2'h2)];
              reg1426 <= $unsigned((~&({(~reg1386),
                      (reg1425 ? reg1435 : (8'ha7)),
                      $signed((7'h57))} ?
                  (~&$unsigned((8'hae))) : $unsigned((~&reg1423)))));
              reg1427 <= (reg1423 - {{$signed($unsigned(reg1414)),
                      {(reg1393 ? reg1431 : reg1438), (reg1433 << reg1435)}},
                  ($signed($unsigned(reg1397)) && reg1414[(5'h18):(4'hb)])});
              reg1429 = reg1433;
              reg1430 <= ({(7'h40)} || {forvar1425[(3'h6):(1'h0)],
                  ((~&(reg1434 ? reg1385 : reg1428)) ?
                      $signed(wire1380[(4'hf):(4'h9)]) : (~$unsigned((7'h49)))),
                  (8'ha4)});
              reg1433 = $unsigned({reg1415[(5'h18):(5'h16)]});
              reg1435 <= (reg1425[(2'h2):(1'h1)] ?
                  ((8'hb6) >= (~^$unsigned(((7'h57) ?
                      reg1415 : reg1440)))) : ($unsigned($unsigned(reg1397)) >> ($unsigned($unsigned((7'h4f))) >= $unsigned(reg1430[(3'h6):(3'h6)]))));
            end
          else
            begin
              reg1429 = (~|$unsigned(({(~reg1425),
                  reg1429[(2'h2):(2'h2)]} >>> wire1378[(4'h8):(3'h4)])));
              reg1433 = {reg1427[(3'h7):(3'h5)],
                  ((^~wire1380[(3'h7):(3'h7)]) << $unsigned($signed({wire1378})))};
              reg1435 <= reg1435;
              reg1437 = $unsigned(((((forvar1425 ? wire1378 : wire1381) ?
                      $signed(wire1377) : (reg1430 ? reg1431 : (7'h4b))) ?
                  ($unsigned(forvar1425) + (!reg1434)) : (8'h9e)) ~^ (({reg1431} == $signed(reg1434)) < reg1414[(5'h18):(5'h12)])));
            end
          if (reg1437[(4'h9):(2'h2)])
            begin
              reg1439 <= wire1381[(3'h5):(2'h2)];
              reg1440 <= $unsigned({reg1432,
                  ($unsigned($unsigned(reg1433)) - (reg1386[(4'hd):(3'h4)] ?
                      wire1422 : reg1436)),
                  (|(reg1424 || $unsigned(reg1436)))});
              reg1441 <= (((&($unsigned((8'hbf)) ?
                      (reg1430 != reg1397) : reg1432[(5'h11):(4'hd)])) ~^ (~^reg1426)) ?
                  ($signed((~&$unsigned(reg1426))) ~^ $signed($unsigned((-reg1397)))) : $signed($unsigned({((8'hb2) ?
                          forvar1425 : reg1386),
                      reg1393[(5'h10):(3'h4)],
                      reg1429[(3'h5):(3'h4)]})));
              reg1442 = ({$signed(reg1412),
                  ($unsigned((wire1378 ? reg1437 : reg1435)) ?
                      $signed($unsigned((7'h47))) : $signed(reg1411[(5'h19):(5'h11)])),
                  {reg1431[(1'h0):(1'h0)],
                      reg1386[(3'h6):(1'h1)]}} ^ ($unsigned($unsigned((reg1385 ?
                      reg1430 : (7'h45)))) ?
                  $unsigned($unsigned((wire1378 ?
                      reg1412 : reg1429))) : (((~^reg1411) ?
                      (~|reg1434) : (wire1381 ?
                          reg1439 : wire1422)) <= $signed((8'hb6)))));
              reg1443 = {reg1437[(1'h0):(1'h0)]};
            end
          else
            begin
              reg1439 <= reg1434;
              reg1442 = $unsigned(reg1437);
              reg1443 = (reg1397 >= {(wire1422[(4'h9):(3'h4)] & reg1432),
                  ($unsigned($unsigned(reg1414)) & (^$signed(reg1443))),
                  $signed(((^reg1397) ?
                      {reg1438, reg1441, forvar1425} : $signed(reg1439)))});
              reg1444 <= {({$unsigned((reg1429 ? reg1442 : (7'h55))),
                          $unsigned(reg1435)} ?
                      reg1436[(3'h7):(2'h3)] : {$unsigned((reg1423 ?
                              reg1439 : reg1434)),
                          $signed((reg1442 ? reg1441 : wire1381)),
                          {reg1443,
                              (reg1423 ? reg1406 : reg1391),
                              (^reg1393)}}),
                  ((^~reg1433) ?
                      {((7'h4b) << $signed(reg1393)),
                          ((reg1443 != reg1436) ?
                              reg1414 : reg1430)} : {(~^reg1426[(5'h15):(5'h12)]),
                          ($unsigned(wire1378) != $signed((7'h50)))})};
              reg1445 <= $unsigned({$unsigned(reg1434),
                  $signed({reg1443, (8'ha0)}),
                  wire1380[(3'h7):(3'h6)]});
              reg1446 <= $signed(reg1424[(4'ha):(3'h6)]);
            end
          reg1447 <= ($unsigned($signed($signed($signed(reg1429)))) << reg1439[(4'hf):(3'h7)]);
          for (forvar1448 = (1'h0); (forvar1448 < (1'h1)); forvar1448 = (forvar1448 + (1'h1)))
            begin
              reg1449 = wire1422[(2'h3):(2'h3)];
            end
          for (forvar1450 = (1'h0); (forvar1450 < (1'h0)); forvar1450 = (forvar1450 + (1'h1)))
            begin
              reg1451 <= $signed($signed({(reg1414 < reg1388[(1'h0):(1'h0)]),
                  (^(~&wire1378))}));
              reg1452 <= {$unsigned($unsigned($signed($signed(reg1397)))),
                  (($unsigned($signed(reg1385)) & (-(&(7'h4a)))) ?
                      $unsigned(reg1427) : wire1380)};
              reg1453 <= (reg1449 ^ {((7'h56) ?
                      reg1452 : $unsigned((reg1391 ? reg1432 : (8'h9c)))),
                  (reg1445 ? reg1406 : $unsigned(reg1442)),
                  $unsigned($unsigned(reg1406))});
            end
          if ({$signed(reg1393),
              ($signed(((forvar1450 == wire1380) - reg1432[(5'h10):(4'hc)])) ?
                  $unsigned(((-(7'h44)) + $signed(reg1432))) : $signed(((reg1427 < reg1432) ?
                      (-reg1424) : wire1381[(3'h4):(3'h4)]))),
              reg1428})
            begin
              reg1454 <= ((8'haa) >= wire1379[(5'h18):(5'h15)]);
              reg1455 = $unsigned(reg1426[(5'h16):(4'hd)]);
            end
          else
            begin
              reg1454 <= reg1443;
              reg1456 <= reg1433[(2'h3):(1'h0)];
              reg1457 = {((~&$signed({reg1432})) ?
                      reg1437 : {(wire1377 ? (reg1426 >>> reg1412) : {(8'hac)}),
                          reg1412}),
                  $signed(($unsigned($unsigned((8'had))) ?
                      {((7'h42) ? reg1391 : (8'hb5)),
                          {forvar1450, reg1451}} : (reg1393 ?
                          (reg1455 ? reg1438 : forvar1448) : (~&reg1438)))),
                  (^~$signed((!$signed((7'h48)))))};
              reg1458 <= ($signed($unsigned((^~forvar1450))) ?
                  reg1434[(5'h14):(5'h12)] : {reg1440[(3'h4):(1'h0)]});
            end
        end
      reg1459 = wire1379[(3'h7):(3'h7)];
    end
  assign wire1460 = $unsigned($signed($signed(reg1426)));
  assign wire1461 = $unsigned((8'hb2));
  assign wire1462 = $signed(reg1435[(5'h10):(5'h10)]);
  always
    @(posedge clk) begin
      if (reg1427)
        begin
          reg1463 <= $signed(wire1381[(2'h3):(2'h2)]);
          reg1464 <= {$unsigned(({((8'hac) && reg1432),
                  $signed(reg1406)} >= {$signed(reg1463)})),
              (~&$unsigned(reg1440[(2'h2):(1'h0)]))};
          reg1465 <= $unsigned($signed($unsigned(((reg1435 << reg1393) || (+reg1452)))));
        end
      else
        begin
          reg1466 = reg1391[(4'h8):(3'h7)];
          reg1467 <= $signed(reg1406[(2'h2):(1'h0)]);
          for (forvar1468 = (1'h0); (forvar1468 < (1'h1)); forvar1468 = (forvar1468 + (1'h1)))
            begin
              reg1469 = (($signed((~&(reg1435 ?
                  reg1453 : reg1430))) != $unsigned(reg1406[(3'h7):(1'h0)])) + {(~^$signed((reg1464 != reg1440)))});
              reg1470 <= (($signed(reg1452[(2'h2):(1'h0)]) + $signed($unsigned($signed(reg1414)))) ?
                  $signed($unsigned(((+wire1460) ?
                      (reg1385 + reg1452) : $signed(reg1463)))) : ((~^{(!reg1456),
                      reg1452[(1'h1):(1'h1)]}) * (((reg1426 ?
                          reg1444 : wire1422) ?
                      reg1435 : $signed(reg1456)) < ({reg1432,
                          reg1430,
                          wire1378} ?
                      (reg1445 ?
                          wire1379 : (7'h51)) : reg1469[(5'h15):(3'h7)]))));
              reg1471 = (-$unsigned(($signed({reg1439,
                  reg1432}) && wire1381[(1'h1):(1'h0)])));
              reg1472 <= $unsigned((((((8'hbd) ^~ (8'ha6)) ?
                  (forvar1468 ?
                      reg1464 : reg1414) : reg1467) == $unsigned((reg1453 ?
                  reg1431 : (8'ha4)))) ~^ reg1466[(3'h7):(2'h3)]));
              reg1473 <= reg1444[(4'h9):(3'h6)];
              reg1474 <= {((^$signed($unsigned(reg1456))) ?
                      $signed(({(8'hb7)} >>> reg1445)) : (7'h52)),
                  {({{reg1463, reg1412, reg1445},
                          {reg1412, reg1435, reg1467},
                          $signed(reg1471)} << ((7'h46) ?
                          (reg1385 ? reg1452 : (7'h4f)) : wire1462)),
                      $signed($signed(reg1473)),
                      $signed((~$signed(reg1430)))}};
            end
          reg1475 = (~((-((~|reg1458) ?
                  ((7'h58) * wire1381) : $unsigned(reg1458))) ?
              (reg1430[(3'h4):(3'h4)] >= $signed((reg1469 ~^ reg1451))) : ($unsigned(reg1456) - ($unsigned(reg1397) >= (^~wire1461)))));
          for (forvar1476 = (1'h0); (forvar1476 < (2'h3)); forvar1476 = (forvar1476 + (1'h1)))
            begin
              reg1477 = (!(^~(reg1414 != reg1453)));
              reg1478 <= reg1414[(5'h19):(4'h8)];
            end
          reg1479 <= $signed($signed((^(^~(reg1444 ? wire1381 : reg1397)))));
        end
      if ($signed(reg1463[(3'h4):(2'h2)]))
        begin
          if ($unsigned((^~$unsigned(((wire1378 ?
              reg1393 : reg1386) | reg1393[(4'he):(3'h4)])))))
            begin
              reg1480 = {reg1393[(1'h1):(1'h1)]};
              reg1481 <= $unsigned((((reg1471 ?
                      (reg1469 ? reg1414 : (7'h48)) : (reg1458 ~^ reg1386)) ?
                  {(reg1436 >> reg1451),
                      (reg1393 ?
                          (8'ha3) : reg1397)} : (&(^~reg1479))) >= reg1393));
              reg1482 = ($signed(reg1479) ^~ reg1430);
              reg1483 <= (~$unsigned($unsigned((~&(reg1469 >> reg1385)))));
              reg1484 = ((8'ha5) && $signed(reg1427[(1'h1):(1'h0)]));
              reg1485 <= (($signed({$unsigned(reg1397),
                  $signed(reg1436)}) >>> $signed(((reg1453 ?
                      reg1388 : (8'haf)) ?
                  $signed((8'hab)) : $unsigned(reg1484)))) || $signed((-$unsigned((-reg1479)))));
              reg1486 <= ((|(wire1380 && (8'hbd))) ?
                  reg1388[(3'h7):(3'h5)] : ($signed((reg1432[(4'h8):(2'h2)] <<< reg1456[(1'h0):(1'h0)])) ?
                      ((+(!(8'hb8))) + (~|reg1444[(2'h2):(1'h1)])) : (~$signed(reg1456[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg1481 <= reg1393[(5'h13):(3'h4)];
              reg1482 = reg1471;
              reg1483 <= reg1430[(3'h4):(1'h1)];
              reg1484 = reg1415[(5'h1b):(3'h7)];
            end
          reg1487 <= ((~^reg1426[(5'h14):(4'hf)]) ?
              ({reg1447[(4'h8):(2'h3)],
                  (~^reg1467[(3'h5):(1'h1)])} >>> $signed($signed((reg1480 ?
                  wire1378 : reg1446)))) : ($unsigned((^~(reg1414 ?
                  wire1379 : reg1439))) ~^ wire1461[(5'h13):(2'h3)]));
          for (forvar1488 = (1'h0); (forvar1488 < (3'h4)); forvar1488 = (forvar1488 + (1'h1)))
            begin
              reg1489 <= {$signed((^{(wire1377 | reg1485),
                      (reg1478 * wire1422),
                      $signed((7'h4a))})),
                  reg1480[(3'h5):(1'h1)]};
            end
        end
      else
        begin
          reg1481 <= reg1472;
          reg1483 <= (($signed(((^~(8'hbb)) <= (~^reg1411))) >= (~^($unsigned(reg1445) ?
              (^reg1484) : reg1478[(1'h1):(1'h0)]))) >= wire1380);
          if ((8'ha1))
            begin
              reg1485 <= (($signed((^{reg1391, reg1469})) ?
                  (|(!{reg1473})) : (((|reg1444) + (8'h9c)) * ((reg1464 * reg1406) ?
                      (reg1385 ?
                          reg1385 : reg1445) : reg1427[(4'he):(4'ha)]))) > (((|$signed(wire1377)) ?
                  (&(reg1425 ? wire1460 : reg1412)) : (reg1472 ?
                      $unsigned(reg1412) : reg1472[(2'h2):(1'h1)])) & reg1456));
              reg1486 <= $signed({($signed({reg1445, reg1412}) >>> {{(8'had),
                          (8'had)},
                      (reg1431 << wire1377)}),
                  {(~$signed(reg1393)), $signed(reg1412)},
                  ($unsigned($unsigned(reg1414)) ?
                      $unsigned($signed(reg1456)) : (~&$signed(reg1465)))});
              reg1488 = $signed($signed($signed((-reg1458[(5'h12):(3'h5)]))));
              reg1490 = reg1445;
              reg1491 <= $unsigned(reg1463);
            end
          else
            begin
              reg1484 = $signed($signed(reg1481));
              reg1488 = ($signed((reg1456[(2'h3):(2'h2)] & ($signed(reg1481) ?
                  reg1414 : $signed(reg1427)))) << reg1475[(2'h2):(1'h1)]);
              reg1490 = reg1470[(4'hb):(4'hb)];
              reg1492 = (~^reg1485[(4'h9):(3'h7)]);
              reg1493 <= reg1477[(4'h8):(3'h6)];
            end
          reg1494 = (!reg1385);
          for (forvar1495 = (1'h0); (forvar1495 < (1'h0)); forvar1495 = (forvar1495 + (1'h1)))
            begin
              reg1496 <= reg1458;
              reg1497 <= $signed(reg1479);
              reg1498 = ($unsigned({($unsigned(reg1488) ?
                          $signed(reg1431) : $unsigned(wire1379)),
                      reg1478}) ?
                  reg1471[(3'h7):(1'h0)] : ($unsigned(($signed(reg1485) != (^~reg1482))) ?
                      (~&((8'hb8) & reg1393[(4'he):(4'h8)])) : (reg1463[(5'h10):(4'ha)] ?
                          $signed(forvar1488[(1'h0):(1'h0)]) : $unsigned(reg1489[(4'hf):(4'hb)]))));
            end
          for (forvar1499 = (1'h0); (forvar1499 < (3'h4)); forvar1499 = (forvar1499 + (1'h1)))
            begin
              reg1500 <= $signed((reg1474[(5'h18):(4'ha)] << $signed(reg1435[(5'h12):(1'h0)])));
              reg1501 <= ($signed((~^{$signed(reg1463),
                      forvar1499[(3'h4):(2'h3)]})) ?
                  reg1482[(2'h3):(2'h2)] : reg1386);
            end
        end
      if ((reg1393 + $signed($signed(reg1439))))
        begin
          for (forvar1502 = (1'h0); (forvar1502 < (2'h2)); forvar1502 = (forvar1502 + (1'h1)))
            begin
              reg1503 = reg1411[(3'h7):(3'h5)];
              reg1504 <= {($signed(((~reg1464) | (reg1385 ?
                      reg1490 : reg1479))) * reg1431[(5'h14):(2'h2)]),
                  ($signed(reg1498) ?
                      (-{reg1486[(4'hf):(3'h7)]}) : (~&$signed((reg1483 ~^ reg1385))))};
              reg1505 <= (&({(reg1440[(3'h5):(2'h2)] ?
                          $signed((8'ha4)) : (reg1480 ?
                              reg1385 : forvar1476))} ?
                  $signed(((reg1446 ? reg1391 : reg1504) ?
                      (reg1441 == (8'hb6)) : wire1462[(1'h0):(1'h0)])) : (reg1494 ?
                      (!(reg1483 ?
                          reg1458 : reg1447)) : (+reg1441[(3'h6):(3'h4)]))));
              reg1506 = reg1386;
            end
          for (forvar1507 = (1'h0); (forvar1507 < (2'h2)); forvar1507 = (forvar1507 + (1'h1)))
            begin
              reg1508 <= $unsigned((~reg1440));
              reg1509 <= reg1447[(3'h6):(2'h2)];
              reg1510 <= (({$signed($signed(reg1426)),
                          ((reg1469 ~^ reg1467) <= $unsigned(reg1406))} ?
                      $signed({(reg1454 ? wire1379 : reg1498),
                          $signed(reg1428)}) : ($unsigned(reg1483) ?
                          $unsigned($signed((8'hb4))) : reg1445[(4'h8):(2'h3)])) ?
                  reg1430[(3'h4):(2'h2)] : forvar1476);
            end
        end
      else
        begin
          reg1502 <= reg1487;
          reg1504 <= wire1461;
          reg1506 = (~&wire1380[(4'h9):(3'h6)]);
          reg1507 <= reg1501[(3'h4):(2'h2)];
        end
      if ($unsigned($unsigned((~(reg1439[(1'h1):(1'h0)] <= $signed(reg1482))))))
        begin
          for (forvar1511 = (1'h0); (forvar1511 < (1'h1)); forvar1511 = (forvar1511 + (1'h1)))
            begin
              reg1512 <= $unsigned($unsigned($signed(({wire1422,
                  forvar1495} >>> (reg1500 ? reg1440 : reg1478)))));
              reg1513 = (~|forvar1495);
              reg1514 <= (~(^~$unsigned(reg1440)));
              reg1515 <= {$unsigned({$unsigned(reg1428)}),
                  {{reg1477}, reg1435, reg1474},
                  reg1485[(3'h4):(3'h4)]};
            end
          reg1516 <= (reg1515 != (7'h45));
          if ($unsigned($signed($unsigned(($unsigned(reg1503) >> (~|reg1411))))))
            begin
              reg1517 = ($unsigned($signed((reg1492 ?
                      $unsigned(reg1467) : $signed(reg1492)))) ?
                  $signed($unsigned(($unsigned(wire1379) ?
                      {reg1430,
                          wire1377,
                          (7'h52)} : (&forvar1507)))) : {reg1464});
              reg1518 = {(((!$signed(reg1412)) + reg1469) ?
                      $unsigned(reg1393) : $signed($signed(wire1378))),
                  $signed(reg1479)};
              reg1519 = (reg1406[(4'hc):(3'h6)] < $signed((~&(8'ha4))));
            end
          else
            begin
              reg1520 <= (&(!$unsigned($unsigned(((8'ha3) || reg1465)))));
            end
          reg1521 <= ($unsigned($unsigned(wire1381[(3'h6):(3'h6)])) ?
              {$signed($unsigned({(8'ha1),
                      reg1480}))} : reg1498[(1'h1):(1'h1)]);
          for (forvar1522 = (1'h0); (forvar1522 < (1'h1)); forvar1522 = (forvar1522 + (1'h1)))
            begin
              reg1523 = $unsigned($signed($signed(((reg1406 ?
                      reg1393 : reg1440) ?
                  (!wire1380) : reg1441[(4'hc):(1'h1)]))));
              reg1524 <= (+$unsigned(($unsigned((~|reg1415)) ?
                  (reg1493[(4'h8):(3'h7)] == $unsigned(reg1488)) : $signed((wire1377 ^ reg1498)))));
              reg1525 <= $signed((~^reg1507));
              reg1526 = forvar1499[(1'h1):(1'h1)];
              reg1527 = (8'hae);
              reg1528 <= ((+(-reg1458[(5'h17):(5'h12)])) ?
                  (-reg1385[(4'hf):(4'ha)]) : {wire1462});
              reg1529 <= $unsigned({(((reg1519 >>> reg1428) ?
                          $unsigned(reg1393) : (~|reg1481)) ?
                      $signed((^reg1513)) : reg1503)});
            end
          reg1530 = (!reg1431[(1'h1):(1'h1)]);
        end
      else
        begin
          for (forvar1511 = (1'h0); (forvar1511 < (1'h1)); forvar1511 = (forvar1511 + (1'h1)))
            begin
              reg1513 = $unsigned($unsigned(reg1516[(4'he):(4'hc)]));
              reg1517 = reg1425;
              reg1518 = reg1514;
            end
          for (forvar1519 = (1'h0); (forvar1519 < (3'h4)); forvar1519 = (forvar1519 + (1'h1)))
            begin
              reg1520 <= (reg1439[(5'h12):(3'h6)] >>> reg1467[(3'h5):(3'h4)]);
              reg1522 = (&$signed($signed(reg1480[(2'h2):(2'h2)])));
            end
          for (forvar1523 = (1'h0); (forvar1523 < (1'h1)); forvar1523 = (forvar1523 + (1'h1)))
            begin
              reg1526 = (reg1519[(5'h12):(3'h4)] ?
                  reg1503 : ($signed(reg1523) - reg1515[(4'hb):(4'h9)]));
              reg1528 <= (reg1496 ~^ $signed(($unsigned(reg1523) ?
                  {((8'haa) ? (7'h46) : reg1444), reg1452} : {{reg1504,
                          reg1432,
                          reg1483}})));
              reg1529 <= {$signed(($signed({reg1503,
                      (7'h42),
                      reg1519}) < $signed($signed(reg1509))))};
              reg1531 <= (8'hb4);
              reg1532 = $signed((({reg1523[(3'h4):(2'h2)],
                      {(8'ha5), forvar1495},
                      forvar1476} ?
                  $unsigned((reg1527 >>> reg1478)) : $signed($signed((8'ha9)))) >> (~&reg1428)));
            end
          for (forvar1533 = (1'h0); (forvar1533 < (3'h6)); forvar1533 = (forvar1533 + (1'h1)))
            begin
              reg1534 <= $unsigned(reg1482);
              reg1535 = $signed((({(reg1470 & reg1509)} ?
                  ($unsigned(wire1380) ?
                      (reg1508 != reg1507) : $unsigned(reg1469)) : $unsigned($signed(reg1406))) >= $signed((&(+reg1425)))));
              reg1536 = $unsigned({$unsigned(((reg1415 ? reg1414 : reg1515) ?
                      (reg1514 ? (8'hb4) : forvar1495) : (reg1411 ?
                          reg1472 : reg1479))),
                  reg1517[(1'h0):(1'h0)]});
              reg1537 = forvar1502[(1'h1):(1'h1)];
              reg1538 = $unsigned((+{$unsigned($unsigned(reg1444)),
                  {reg1391, $unsigned((7'h48))},
                  ((forvar1533 ? reg1490 : forvar1495) <<< {forvar1523})}));
              reg1539 = (&(8'h9e));
            end
          reg1540 = ($unsigned((reg1524 ?
                  reg1530[(5'h11):(5'h10)] : $unsigned((reg1522 ?
                      forvar1519 : (8'h9d))))) ?
              forvar1533 : reg1431);
          reg1541 = forvar1468[(4'hc):(3'h7)];
        end
      reg1542 = $unsigned(reg1528[(4'hf):(4'hd)]);
      if ((^((($signed((8'haf)) ^ (^~reg1427)) ?
              (!{forvar1488}) : ({reg1490, reg1412} >>> $signed(wire1380))) ?
          $signed($signed(reg1542)) : (|(&$signed(reg1414))))))
        begin
          reg1543 = $signed((($unsigned({reg1542}) ?
                  $unsigned($unsigned((7'h53))) : $signed(reg1425[(2'h2):(2'h2)])) ?
              ({(reg1489 > reg1530)} && forvar1495[(5'h11):(4'h8)]) : (7'h40)));
          for (forvar1544 = (1'h0); (forvar1544 < (2'h3)); forvar1544 = (forvar1544 + (1'h1)))
            begin
              reg1545 <= ($unsigned(reg1505[(3'h6):(2'h2)]) == {({$unsigned(reg1465)} || $signed((^reg1406))),
                  reg1447,
                  ($signed($unsigned((7'h53))) >= ($unsigned(reg1494) >= reg1497))});
              reg1546 <= $unsigned(reg1458[(3'h6):(3'h4)]);
              reg1547 <= $signed(reg1469[(4'hd):(4'h8)]);
              reg1548 = reg1535[(3'h7):(1'h1)];
            end
        end
      else
        begin
          if (reg1489)
            begin
              reg1544 <= $signed($signed((-((+reg1393) ?
                  (-reg1386) : reg1430[(3'h4):(1'h0)]))));
              reg1545 <= ($signed(reg1490) ?
                  reg1518 : {reg1465[(1'h0):(1'h0)]});
              reg1548 = (~|forvar1502);
              reg1549 = {$unsigned(((7'h42) ?
                      ((reg1473 ?
                          reg1439 : reg1535) > (reg1493 > reg1430)) : (+$signed(reg1445))))};
            end
          else
            begin
              reg1544 <= $signed($unsigned(($unsigned($unsigned(reg1428)) | ((^(8'h9e)) < $signed(reg1487)))));
              reg1548 = reg1492[(2'h2):(1'h1)];
              reg1550 <= (((reg1496 ?
                          {reg1534[(4'h8):(2'h3)],
                              (+reg1430),
                              $signed((7'h56))} : reg1508) ?
                      (($signed(reg1441) ^ reg1525) <<< ({(7'h4c)} ?
                          ((7'h48) ?
                              reg1493 : (8'hb3)) : reg1464[(5'h14):(2'h3)])) : reg1447) ?
                  $unsigned(reg1475[(1'h1):(1'h1)]) : $signed({{reg1465},
                      reg1544[(5'h12):(4'he)]}));
              reg1551 = $signed(((~reg1543) ?
                  ((((8'ha8) ?
                      forvar1495 : reg1385) ~^ (forvar1502 ^ (7'h48))) << (~^reg1439[(5'h15):(5'h12)])) : $unsigned(($unsigned(reg1493) ?
                      (reg1534 & reg1496) : reg1497[(2'h3):(1'h0)]))));
              reg1552 <= reg1515[(4'ha):(4'ha)];
              reg1553 <= reg1496;
            end
          reg1554 = ((-reg1515) & (~^{wire1378}));
          reg1555 = forvar1522[(4'he):(2'h2)];
          reg1556 <= ({$unsigned(({reg1490} ?
                      $unsigned(forvar1476) : (~reg1458))),
                  ($signed($signed(reg1512)) < $signed(reg1479))} ?
              $unsigned((!reg1528)) : ($unsigned(forvar1519) ?
                  ((-$unsigned(reg1471)) ?
                      $unsigned({reg1482,
                          reg1452,
                          reg1451}) : $signed(reg1531[(4'hf):(4'he)])) : {reg1411[(4'hb):(3'h6)],
                      ($unsigned(reg1516) == (+reg1498)),
                      (-(!reg1435))}));
          reg1557 = reg1487[(4'hc):(3'h6)];
          for (forvar1558 = (1'h0); (forvar1558 < (3'h5)); forvar1558 = (forvar1558 + (1'h1)))
            begin
              reg1559 <= $unsigned(forvar1476);
              reg1560 <= reg1430[(3'h4):(1'h0)];
              reg1561 <= (!$signed((reg1504[(4'he):(4'hc)] ~^ forvar1558[(2'h3):(2'h2)])));
              reg1562 = ($signed((({reg1446, reg1529, (8'hb7)} ?
                      reg1517[(2'h2):(1'h1)] : $signed(reg1526)) >>> (~^reg1487[(3'h6):(2'h3)]))) ?
                  (&((((7'h40) == (7'h45)) >>> $unsigned(reg1386)) || {(forvar1507 == reg1544),
                      $signed((8'ha7)),
                      (reg1487 * reg1502)})) : (reg1447[(4'hf):(4'hc)] <= (^(+((7'h51) ?
                      reg1504 : reg1546)))));
              reg1563 <= {(~&$unsigned(reg1496)),
                  ($unsigned(((reg1474 ^ forvar1511) ?
                      (~^reg1496) : $unsigned(forvar1522))) ^~ (~{(reg1483 ?
                          (8'hbd) : reg1456),
                      {(8'had), reg1477, reg1456},
                      $signed(reg1503)}))};
              reg1564 <= {reg1482[(2'h3):(2'h3)],
                  $unsigned((^~(reg1563[(5'h11):(1'h0)] ^ reg1454))),
                  ((reg1435[(5'h14):(2'h3)] <= reg1498) ?
                      $unsigned(((^~reg1483) ?
                          $signed(wire1380) : reg1453[(3'h4):(1'h0)])) : (((reg1519 ?
                              (7'h4b) : (7'h49)) | reg1513[(5'h11):(5'h10)]) ?
                          ({reg1515, reg1554} ?
                              reg1513[(4'he):(4'he)] : (~|reg1432)) : ($signed(reg1463) ^ reg1562[(3'h5):(2'h2)])))};
              reg1565 <= {reg1466,
                  ((&$signed((reg1483 ? reg1564 : reg1532))) ?
                      (8'hac) : {$signed($signed(reg1464)),
                          (reg1502 | (^~reg1466))}),
                  {(^$signed($unsigned(reg1504))),
                      ({reg1412[(2'h2):(1'h1)],
                          (reg1524 - reg1553),
                          ((8'hb6) ^~ reg1444)} ^~ ($unsigned(wire1379) ^~ (forvar1519 && reg1436))),
                      $unsigned(reg1385)}};
            end
        end
    end
  assign wire1566 = (&(((reg1528[(5'h1b):(5'h1a)] | $unsigned((7'h51))) + {{reg1446,
                            (8'hb5)}}) * reg1496[(5'h13):(3'h6)]));
  assign wire1567 = reg1561[(4'h8):(1'h0)];
  always
    @(posedge clk) begin
      reg1568 <= ($signed({reg1485,
          {$signed(reg1489)},
          (&reg1485[(3'h7):(3'h6)])}) * (|reg1509[(5'h18):(4'h8)]));
      for (forvar1569 = (1'h0); (forvar1569 < (1'h0)); forvar1569 = (forvar1569 + (1'h1)))
        begin
          reg1570 = reg1481;
          reg1571 = (^~(&$unsigned(reg1485[(4'h9):(4'h9)])));
          if (reg1544)
            begin
              reg1572 <= $unsigned((~reg1445[(1'h1):(1'h1)]));
              reg1573 <= reg1572[(2'h2):(1'h0)];
              reg1574 = (~$signed((($signed((7'h4a)) ?
                      $signed(reg1427) : $unsigned(reg1509)) ?
                  (reg1464 > $signed(reg1508)) : reg1485[(3'h4):(2'h3)])));
              reg1575 <= (+{reg1447[(3'h5):(1'h1)],
                  (reg1556[(2'h2):(1'h0)] | (reg1529 && reg1426))});
            end
          else
            begin
              reg1574 = (reg1573[(3'h6):(3'h5)] ?
                  {($signed((7'h48)) ?
                          ($signed((8'ha4)) ^~ reg1430[(3'h4):(3'h4)]) : ((8'ha0) || ((8'ha9) ?
                              reg1393 : reg1507))),
                      reg1451} : $unsigned($signed((&{reg1427, (7'h58)}))));
              reg1575 <= reg1521[(1'h0):(1'h0)];
              reg1576 <= ($signed((reg1510[(4'h8):(3'h5)] >>> ((reg1473 ?
                      forvar1569 : (7'h53)) + (~|reg1544)))) ?
                  $signed((((wire1377 * (8'hbf)) ?
                      wire1461 : {reg1440,
                          reg1474,
                          reg1544}) + (~(~^reg1505)))) : reg1436[(4'h9):(3'h4)]);
              reg1577 <= $signed($signed($signed($signed(reg1550))));
              reg1578 = reg1508[(5'h14):(4'hf)];
              reg1579 = (wire1378 || $unsigned((reg1428 & (reg1447 ~^ $unsigned(reg1427)))));
              reg1580 = (~|({wire1377[(4'h9):(1'h0)],
                  $signed($unsigned((7'h57))),
                  (forvar1569[(4'hd):(1'h0)] ?
                      (!reg1534) : (^~reg1458))} ^~ reg1552));
            end
          reg1581 <= $unsigned((~^($signed(reg1550[(4'h8):(3'h6)]) ?
              reg1520 : $signed((reg1483 | reg1472)))));
        end
      reg1582 <= (~&(reg1556 ?
          {{(~&(7'h4f))}} : (reg1577[(1'h1):(1'h1)] ?
              (&(-reg1496)) : ({reg1478, reg1577} ?
                  reg1560[(5'h17):(4'hc)] : $unsigned(reg1467)))));
    end
  assign wire1583 = $signed(reg1561[(4'hc):(4'ha)]);
  assign wire1584 = (reg1568[(3'h5):(2'h2)] || $signed($unsigned((!(reg1452 ?
                        (8'h9d) : reg1479)))));
  assign wire1585 = reg1561[(5'h11):(4'ha)];
  always
    @(posedge clk) begin
      if ($unsigned($signed(reg1458[(5'h10):(2'h3)])))
        begin
          for (forvar1586 = (1'h0); (forvar1586 < (3'h5)); forvar1586 = (forvar1586 + (1'h1)))
            begin
              reg1587 = $signed({(~^{(reg1508 * reg1493)}),
                  $signed(((reg1415 ? reg1556 : wire1381) ?
                      reg1563 : (forvar1586 ? reg1534 : forvar1586))),
                  $unsigned($signed($unsigned((7'h40))))});
              reg1588 <= reg1546[(4'h9):(4'h9)];
              reg1589 <= reg1411[(5'h12):(5'h10)];
              reg1590 <= $unsigned($signed((reg1445[(5'h11):(4'hd)] ?
                  wire1461 : ((reg1445 ?
                      reg1386 : reg1510) + $unsigned((7'h51))))));
              reg1591 <= (({($unsigned(reg1552) ?
                              $unsigned(wire1584) : (~&(8'hbf))),
                          $unsigned((~^reg1393)),
                          ((reg1544 & (7'h45)) - (reg1544 * (8'ha4)))} ?
                      (-($unsigned(reg1510) ?
                          $unsigned(wire1422) : (reg1441 * forvar1586))) : reg1431[(5'h13):(3'h4)]) ?
                  (^(forvar1586 * reg1406[(3'h4):(2'h2)])) : reg1573);
            end
          if (reg1500)
            begin
              reg1592 <= ({($signed($signed(reg1544)) == $signed(reg1478)),
                      $signed($unsigned((^~reg1582)))} ?
                  (reg1500[(2'h3):(2'h2)] < $unsigned(((-reg1465) >> ((8'hb4) & reg1552)))) : ($signed($unsigned(reg1391)) ?
                      {$unsigned($signed((7'h47)))} : $signed(wire1381[(1'h0):(1'h0)])));
              reg1593 <= reg1502;
            end
          else
            begin
              reg1594 = {$signed(reg1545)};
              reg1595 <= (-reg1465);
              reg1596 = reg1559[(2'h2):(1'h0)];
              reg1597 = $unsigned((reg1406 ?
                  (($unsigned(reg1428) ?
                      reg1577[(1'h1):(1'h0)] : (reg1414 ?
                          reg1556 : reg1577)) ^ wire1422) : reg1414[(3'h6):(2'h2)]));
              reg1598 <= reg1591[(3'h4):(3'h4)];
              reg1599 <= ({reg1428, reg1576} ?
                  (|($unsigned($signed(reg1489)) ?
                      (reg1563 ? $signed((8'hb1)) : (8'ha3)) : {{reg1415,
                              reg1385,
                              reg1597}})) : $unsigned((-((wire1380 & reg1452) | (7'h53)))));
              reg1600 <= ($unsigned($unsigned(((reg1414 != wire1583) ?
                  (-reg1446) : $unsigned(reg1531)))) <= (|{reg1426[(1'h0):(1'h0)],
                  (reg1453 - $signed(reg1412))}));
            end
          reg1601 <= reg1415;
          for (forvar1602 = (1'h0); (forvar1602 < (3'h4)); forvar1602 = (forvar1602 + (1'h1)))
            begin
              reg1603 = $unsigned(((reg1520[(2'h2):(1'h1)] * $unsigned((reg1415 ?
                  reg1489 : wire1377))) > {(|reg1425),
                  $signed(reg1483),
                  reg1504}));
              reg1604 <= (&reg1510[(2'h3):(2'h2)]);
              reg1605 = $unsigned(reg1474[(4'hd):(4'ha)]);
              reg1606 <= $unsigned(($signed(($signed(reg1385) ?
                      $signed(wire1585) : reg1601[(1'h1):(1'h0)])) ?
                  reg1451[(2'h3):(1'h0)] : (($signed(reg1431) >= $signed(reg1529)) ?
                      $unsigned((reg1452 ? reg1568 : reg1426)) : (reg1594 ?
                          (7'h56) : {reg1596}))));
              reg1607 <= ($unsigned(($unsigned({reg1596,
                  (8'hbd),
                  reg1512}) >= (|wire1567))) >> (((reg1456 ?
                  (~reg1465) : (|reg1415)) && $signed($unsigned((7'h4a)))) ^~ $unsigned(reg1546[(2'h3):(2'h2)])));
              reg1608 <= $signed(reg1588);
            end
          if ((~^(~&$unsigned(({reg1464} ?
              (reg1564 ? reg1452 : reg1600) : (&wire1422))))))
            begin
              reg1609 = reg1415;
              reg1610 = $signed($unsigned(((~(reg1559 ^~ reg1572)) || ((reg1604 && wire1583) ?
                  (~reg1507) : $signed((8'hbc))))));
              reg1611 <= $signed((~|($signed($signed(reg1606)) ?
                  (&{reg1436, (8'hb9), reg1552}) : (7'h54))));
              reg1612 = ((|$unsigned($unsigned(reg1467[(3'h4):(1'h0)]))) ?
                  ((((reg1446 | reg1599) != ((8'h9e) ?
                      reg1439 : (8'hbf))) & reg1391) >> $signed({$unsigned(reg1473),
                      $signed(reg1386)})) : $signed({$unsigned((reg1412 || reg1582))}));
              reg1613 <= $signed(wire1461);
              reg1614 <= $signed($signed($unsigned(reg1590[(5'h19):(4'he)])));
            end
          else
            begin
              reg1611 <= (-reg1464[(5'h12):(1'h0)]);
              reg1612 = (({((!reg1397) ?
                          reg1391[(4'h8):(4'h8)] : $unsigned((7'h49))),
                      $unsigned($signed(reg1589)),
                      {reg1510}} ?
                  (~reg1600) : $signed(reg1525[(4'ha):(4'h8)])) >>> {$unsigned(reg1481),
                  (&(reg1572[(2'h3):(1'h1)] + $unsigned(reg1593))),
                  reg1425[(3'h4):(3'h4)]});
              reg1613 <= (~|{{($signed(reg1435) ?
                          (reg1592 ? reg1524 : reg1406) : (~|reg1458)),
                      reg1546[(2'h2):(1'h0)],
                      reg1453[(5'h16):(5'h11)]}});
              reg1614 <= (&$signed(forvar1586[(4'hc):(3'h5)]));
              reg1615 = $unsigned(reg1487);
              reg1616 = $signed(reg1561[(3'h7):(2'h2)]);
              reg1617 <= reg1439[(3'h5):(1'h1)];
            end
          for (forvar1618 = (1'h0); (forvar1618 < (3'h6)); forvar1618 = (forvar1618 + (1'h1)))
            begin
              reg1619 <= $signed($unsigned(((^reg1489) ?
                  (reg1439[(5'h12):(4'h8)] ?
                      $signed(reg1444) : (reg1465 ?
                          reg1508 : reg1487)) : (~reg1604[(3'h6):(2'h3)]))));
            end
          reg1620 = {{$signed((&(reg1458 ? reg1600 : reg1599))),
                  $unsigned($signed($signed((7'h4d))))},
              (~$signed(({forvar1586, reg1572} ?
                  reg1444 : ((8'ha9) + wire1566)))),
              $unsigned((((~|reg1520) ?
                      (reg1609 >= wire1566) : (reg1453 ? (8'hb8) : reg1491)) ?
                  $signed(reg1610[(3'h6):(2'h3)]) : $unsigned(reg1447)))};
        end
      else
        begin
          for (forvar1586 = (1'h0); (forvar1586 < (2'h2)); forvar1586 = (forvar1586 + (1'h1)))
            begin
              reg1587 = $signed($signed($unsigned(reg1504)));
              reg1594 = (reg1588[(1'h1):(1'h0)] && {(8'hba)});
              reg1595 <= reg1445[(4'hb):(3'h5)];
              reg1596 = (reg1594 ? reg1550[(4'hc):(3'h4)] : reg1430);
            end
          reg1597 = reg1573[(3'h4):(1'h0)];
          reg1598 <= (($unsigned(reg1614[(1'h0):(1'h0)]) << (^~(8'hac))) + $unsigned(({(reg1598 ?
                  reg1617 : reg1591),
              $unsigned(reg1534),
              (reg1415 >>> reg1501)} | forvar1602)));
          if ($signed(reg1552))
            begin
              reg1599 <= ($signed((reg1510[(4'hc):(3'h7)] ~^ (((8'ha5) ?
                  wire1380 : reg1587) | reg1521))) | $signed((reg1507[(5'h17):(4'hb)] >> (+((8'hbc) < reg1414)))));
              reg1600 <= wire1378;
            end
          else
            begin
              reg1599 <= reg1463[(4'he):(4'ha)];
              reg1602 = {$unsigned(reg1614[(2'h2):(1'h1)]),
                  (reg1521[(1'h1):(1'h1)] ?
                      {reg1559,
                          wire1381[(3'h6):(3'h4)],
                          $unsigned({reg1431})} : $unsigned(reg1458))};
              reg1603 = ((&{reg1425}) >> $unsigned((({reg1591} ?
                  reg1581 : $unsigned(reg1441)) ^~ (8'h9f))));
              reg1605 = (($signed(reg1608[(5'h12):(4'h9)]) ?
                  $unsigned(($unsigned(reg1592) > (reg1553 ?
                      (8'hb3) : reg1603))) : ($signed(reg1588) + reg1603)) >= $unsigned(reg1534[(4'hc):(2'h3)]));
              reg1609 = {reg1568,
                  forvar1602[(4'h8):(4'h8)],
                  (((8'ha0) ?
                      (^{reg1559}) : ((!reg1473) ?
                          (reg1464 >>> reg1485) : $signed(reg1386))) >= $unsigned(($unsigned(reg1525) | reg1616)))};
            end
          reg1610 = $signed((|(reg1609[(4'ha):(1'h1)] >>> ($signed(reg1531) != (!reg1573)))));
          reg1611 <= reg1591;
          reg1613 <= $signed($unsigned((~|reg1561[(4'h9):(4'h9)])));
        end
      reg1621 = reg1559[(4'h8):(3'h4)];
      if (reg1587[(1'h1):(1'h0)])
        begin
          for (forvar1622 = (1'h0); (forvar1622 < (1'h0)); forvar1622 = (forvar1622 + (1'h1)))
            begin
              reg1623 <= (reg1576[(4'h8):(4'h8)] ?
                  (reg1436 ? wire1566 : reg1485) : reg1512);
              reg1624 <= $unsigned((^$signed($signed((forvar1586 + reg1605)))));
              reg1625 <= $unsigned($signed(($unsigned((reg1609 ?
                  reg1561 : reg1613)) != $signed((7'h4e)))));
            end
          if (($unsigned($signed($unsigned($unsigned((8'hb0))))) ?
              $signed({forvar1622}) : (~(~^$signed((~&reg1573))))))
            begin
              reg1626 <= $signed($unsigned(reg1621));
              reg1627 = $signed((~reg1613[(4'hc):(1'h1)]));
              reg1628 = $unsigned((+reg1521));
              reg1629 = $unsigned($signed((~^reg1600)));
            end
          else
            begin
              reg1627 = (^reg1516[(5'h17):(5'h16)]);
              reg1628 = {(^~$signed(($signed(reg1478) < $unsigned(wire1584)))),
                  (7'h42),
                  (^{$unsigned(((8'ha3) ^~ reg1565))})};
              reg1630 <= (reg1411[(5'h11):(4'hb)] || reg1415[(5'h1e):(5'h14)]);
              reg1631 <= ((reg1491[(3'h4):(2'h2)] ?
                  {$signed((~reg1601)),
                      ((&wire1461) + (~^reg1630)),
                      (+(+reg1629))} : $signed(reg1456)) >>> reg1486);
              reg1632 = reg1616;
              reg1633 <= ($signed(reg1613) ?
                  (~|reg1425) : (reg1564 ?
                      ({(^reg1628),
                              reg1577[(1'h0):(1'h0)],
                              ((8'hba) ? reg1440 : reg1520)} ?
                          reg1556 : {(reg1508 ?
                                  reg1589 : reg1500)}) : {(~(reg1531 - reg1388))}));
              reg1634 = reg1452[(2'h2):(1'h1)];
            end
          reg1635 = $signed($signed(reg1606[(4'hd):(4'hb)]));
          for (forvar1636 = (1'h0); (forvar1636 < (3'h4)); forvar1636 = (forvar1636 + (1'h1)))
            begin
              reg1637 <= $signed((8'ha6));
            end
          for (forvar1638 = (1'h0); (forvar1638 < (2'h3)); forvar1638 = (forvar1638 + (1'h1)))
            begin
              reg1639 <= ($signed((8'hbd)) >> reg1435);
              reg1640 = ((reg1473[(3'h4):(1'h0)] > (-$signed(reg1504))) ?
                  $signed((forvar1636 & (!$unsigned(reg1391)))) : ({(8'h9d),
                      $signed((!wire1380))} == (|(&$unsigned((8'hb5))))));
              reg1641 <= $unsigned(reg1593);
              reg1642 <= $signed(reg1564[(2'h2):(1'h0)]);
            end
          reg1643 <= (wire1378[(3'h4):(2'h2)] >> {(($unsigned((8'ha5)) != (reg1568 ?
                  (8'hb1) : (8'ha1))) - (&reg1444[(5'h12):(4'ha)])),
              {(|{reg1454}),
                  ({(7'h4d), reg1564} ? (reg1573 >>> reg1564) : wire1378),
                  reg1546[(2'h2):(1'h0)]},
              ($unsigned($unsigned(reg1576)) << reg1639)});
        end
      else
        begin
          reg1622 <= {$signed(((reg1577 >= (~&(7'h56))) ?
                  reg1588 : $signed((reg1528 >>> reg1639)))),
              $signed((wire1567[(4'h9):(3'h4)] <= (^~reg1444)))};
          reg1627 = $signed(({($signed(reg1613) ?
                  (reg1528 >> reg1528) : $signed((7'h40)))} ~^ $unsigned($signed((~&wire1462)))));
          reg1630 <= reg1593[(1'h0):(1'h0)];
          if ((^$unsigned($signed($signed(reg1529)))))
            begin
              reg1632 = $unsigned($unsigned(({(!reg1454),
                  (reg1485 ? reg1575 : reg1629)} << (+((8'had) ?
                  reg1515 : reg1613)))));
              reg1633 <= $signed((~^((reg1439[(5'h11):(2'h3)] ?
                  (~|reg1561) : (reg1615 * wire1461)) < $unsigned(reg1613[(5'h17):(4'h9)]))));
              reg1634 = (reg1598[(3'h7):(1'h0)] <<< (~&$signed((~^(&reg1577)))));
            end
          else
            begin
              reg1632 = (reg1487[(4'hd):(3'h5)] ?
                  ((reg1593 ?
                      (wire1379 ?
                          forvar1618[(2'h2):(1'h0)] : reg1531) : reg1594[(4'ha):(3'h4)]) <<< (~&reg1547[(3'h4):(1'h0)])) : $signed((((reg1486 ?
                          reg1556 : reg1415) && reg1486) ?
                      reg1626[(4'hc):(1'h0)] : ({reg1613, reg1493, reg1588} ?
                          reg1454 : (~&reg1611)))));
              reg1634 = reg1611[(5'h12):(5'h12)];
            end
          reg1635 = $signed($unsigned(($signed($signed((7'h4f))) != wire1584[(3'h5):(2'h3)])));
        end
      reg1644 <= reg1504[(2'h2):(2'h2)];
      reg1645 <= reg1575;
      reg1646 = reg1605;
    end
  assign wire1647 = (-$unsigned(reg1493[(3'h6):(2'h3)]));
  assign wire1648 = (((((reg1617 + (8'had)) || $unsigned(reg1565)) >> $signed(reg1451[(5'h11):(4'ha)])) ?
                        (!reg1505) : (~&($unsigned(reg1534) ?
                            reg1479[(5'h12):(4'hb)] : reg1524))) << (^$signed((^{(7'h4c),
                        reg1385,
                        reg1553}))));
  always
    @(posedge clk) begin
      reg1649 = ((({(reg1529 ? reg1431 : reg1613),
              (reg1510 ? (7'h57) : reg1445)} ?
          reg1436[(4'h8):(1'h0)] : ($unsigned(reg1600) + $unsigned(wire1584))) != $unsigned((~^(7'h58)))) ~^ {($signed(reg1515) ?
              $signed($signed(reg1501)) : $signed((reg1633 ?
                  reg1624 : reg1478)))});
      if (((+$signed($unsigned(reg1446))) ?
          (((8'ha4) ?
                  $signed((reg1582 || reg1426)) : $unsigned((wire1585 << (7'h40)))) ?
              reg1520[(1'h1):(1'h0)] : $signed($unsigned($unsigned(reg1456)))) : (($unsigned((8'hb0)) * $unsigned(wire1584[(1'h1):(1'h0)])) ?
              reg1598[(2'h2):(1'h1)] : (+((reg1453 ? reg1576 : (8'hb7)) ?
                  (wire1422 != reg1414) : reg1573[(2'h3):(1'h0)])))))
        begin
          reg1650 <= $unsigned(reg1625);
          if (reg1485[(4'hc):(2'h2)])
            begin
              reg1651 = (7'h4a);
              reg1652 <= $signed({((reg1439 ?
                          (reg1465 + reg1486) : (reg1486 ? reg1452 : reg1623)) ?
                      $signed((8'ha9)) : (~&$unsigned(reg1637))),
                  (^~(-((7'h4c) & (8'hba)))),
                  {(reg1393 > wire1584[(3'h4):(3'h4)]),
                      $unsigned((reg1501 ? reg1624 : reg1483))}});
              reg1653 = (^((&(reg1391 >= reg1644[(4'hc):(3'h6)])) << (^~$signed($unsigned(reg1652)))));
              reg1654 = (7'h49);
              reg1655 = reg1644;
              reg1656 = $signed(reg1491[(4'he):(3'h6)]);
              reg1657 = ($signed({reg1478[(3'h6):(3'h4)]}) ?
                  ((~^$signed($signed(reg1501))) ?
                      reg1655 : reg1508[(2'h2):(1'h0)]) : $signed((7'h41)));
            end
          else
            begin
              reg1652 <= (+(8'hb6));
              reg1658 <= reg1426;
              reg1659 = $signed({reg1608,
                  ((^~reg1445[(4'he):(1'h0)]) * $signed($signed(reg1576))),
                  reg1432});
              reg1660 <= reg1630;
              reg1661 <= reg1441[(4'hc):(4'h9)];
              reg1662 <= $signed((((8'hb7) ?
                  reg1524 : ($unsigned(wire1648) * reg1453[(5'h15):(4'hf)])) != $signed((~^$signed(wire1461)))));
              reg1663 <= reg1425;
            end
          reg1664 = $signed(reg1496);
        end
      else
        begin
          reg1650 <= ($signed(reg1614) ?
              (reg1599 ?
                  $unsigned($unsigned({reg1565})) : {((wire1648 ?
                          reg1653 : reg1444) >>> ((8'hae) ^~ wire1584)),
                      reg1651[(2'h2):(2'h2)],
                      reg1426[(5'h13):(4'hf)]}) : reg1553[(4'hb):(4'h8)]);
        end
    end
  always
    @(posedge clk) begin
      reg1665 = $unsigned((~|((~^reg1397[(3'h5):(2'h2)]) >= $unsigned(reg1427))));
      reg1666 = (!reg1483[(2'h2):(1'h0)]);
      reg1667 = (|$signed(($unsigned($signed(reg1521)) | reg1391)));
    end
  assign wire1668 = reg1590;
  assign wire1669 = $unsigned($unsigned($signed(reg1630)));
  always
    @(posedge clk) begin
      if ((~&(($signed($signed(reg1525)) && ($signed(wire1648) * (reg1467 ?
          reg1606 : reg1441))) != (|$signed($signed(reg1560))))))
        begin
          reg1670 <= {$unsigned(reg1534), (-(~reg1619[(4'h8):(3'h6)]))};
          reg1671 <= reg1556;
        end
      else
        begin
          if ({(&{(~&(reg1631 ? (8'hbe) : reg1473)),
                  {reg1414, $signed(reg1661), $unsigned(reg1595)}}),
              reg1520[(2'h2):(1'h1)]})
            begin
              reg1670 <= $signed((wire1566 ?
                  $signed(wire1668[(2'h3):(1'h1)]) : (!$signed($unsigned(reg1500)))));
              reg1671 <= wire1668[(1'h1):(1'h0)];
              reg1672 = ($signed((reg1427 ?
                      reg1568[(5'h13):(4'hc)] : (~$signed(reg1397)))) ?
                  $unsigned(reg1452[(2'h3):(2'h2)]) : $unsigned(((~(~reg1573)) ?
                      ((+reg1604) && $signed(wire1462)) : $signed((&reg1592)))));
              reg1673 <= (reg1560[(4'hc):(1'h1)] ?
                  ($signed((reg1456[(3'h4):(2'h3)] ?
                          $signed(reg1544) : reg1606)) ?
                      $unsigned({(~^reg1510),
                          reg1412,
                          $signed(reg1504)}) : ($signed((reg1652 >>> (8'hb6))) >> (wire1583 > reg1393))) : (reg1593[(3'h7):(2'h2)] ?
                      reg1576 : ({(~&reg1661)} ~^ $unsigned((^~reg1454)))));
              reg1674 = ($unsigned($signed($unsigned((reg1561 <= reg1658)))) ?
                  reg1509[(3'h5):(2'h3)] : {($unsigned(((8'hb1) | reg1432)) ?
                          (~|(reg1525 ^ reg1626)) : reg1444[(4'hb):(2'h2)]),
                      $signed((reg1588 && (wire1585 ? reg1547 : reg1606)))});
            end
          else
            begin
              reg1670 <= $signed((-$unsigned($signed((reg1486 ?
                  reg1607 : reg1510)))));
            end
          reg1675 = reg1491[(3'h7):(3'h4)];
          reg1676 = $unsigned(reg1393);
          if ($signed(reg1591[(1'h1):(1'h0)]))
            begin
              reg1677 = reg1575;
              reg1678 <= (($unsigned((!(reg1650 + reg1545))) ?
                      ({wire1583[(3'h6):(3'h5)],
                          (^~reg1388)} <<< $signed(reg1563[(1'h1):(1'h1)])) : reg1673) ?
                  $unsigned(reg1637) : $signed(reg1599));
              reg1679 = reg1645;
              reg1680 = (reg1456[(3'h4):(1'h1)] << reg1677);
              reg1681 <= wire1583;
              reg1682 <= ((($signed(reg1622[(3'h4):(1'h0)]) ?
                      ($unsigned(reg1590) ?
                          {reg1496} : reg1681) : $unsigned($signed(reg1504))) | (reg1604 - ((reg1550 || reg1510) ?
                      (reg1545 + reg1674) : (reg1486 && wire1462)))) ?
                  $unsigned($signed({$signed(reg1608)})) : ((wire1378[(1'h1):(1'h0)] ?
                      (reg1614[(2'h3):(2'h2)] ?
                          (reg1534 ?
                              reg1639 : reg1613) : reg1528[(4'h9):(2'h2)]) : ({reg1622,
                              reg1411} ?
                          $signed((7'h49)) : (reg1660 ^ (7'h44)))) < ($signed((reg1521 ?
                          (8'hbf) : reg1452)) ?
                      (-(~^reg1520)) : $signed(reg1556[(2'h2):(1'h1)]))));
              reg1683 <= $unsigned(reg1516[(5'h1e):(2'h2)]);
            end
          else
            begin
              reg1678 <= ($signed((+(((7'h46) ? reg1546 : reg1670) ?
                      (reg1559 && (8'ha7)) : reg1452[(2'h2):(1'h1)]))) ?
                  (~&(reg1552[(4'hd):(1'h1)] ?
                      reg1675[(1'h0):(1'h0)] : ((reg1581 >>> reg1561) | reg1486[(2'h2):(1'h0)]))) : {(((wire1462 + (7'h43)) ?
                              (|reg1458) : $unsigned(reg1502)) ?
                          $signed(reg1673) : ((&(8'hb3)) ~^ $signed(reg1441))),
                      ($unsigned($unsigned(reg1463)) ?
                          (&(~reg1575)) : (~&reg1607[(2'h3):(2'h2)])),
                      (7'h55)});
              reg1681 <= $unsigned(({{$signed(reg1556),
                          (wire1460 ? reg1544 : reg1568),
                          reg1670},
                      reg1588,
                      reg1415} ?
                  ($unsigned($unsigned(reg1658)) ?
                      (7'h42) : reg1406) : $signed(reg1485)));
              reg1684 = reg1674[(3'h6):(3'h4)];
              reg1685 <= reg1600;
            end
          if ((~&(~(&$unsigned($unsigned(wire1379))))))
            begin
              reg1686 = (($signed(($unsigned(reg1464) ?
                  (^~reg1572) : $signed((8'ha4)))) <<< reg1479) - reg1525);
              reg1687 <= $unsigned(({reg1491} << $signed(reg1512)));
              reg1688 <= (&(($signed(((8'ha1) ? reg1582 : reg1601)) ?
                  $signed(reg1644) : (&((8'h9d) ?
                      reg1451 : wire1669))) & ((-$signed(reg1473)) ?
                  $unsigned($signed(reg1593)) : $unsigned((reg1440 == reg1560)))));
              reg1689 <= reg1593[(2'h3):(2'h3)];
              reg1690 <= (8'ha8);
            end
          else
            begin
              reg1686 = {reg1474,
                  (reg1472[(1'h1):(1'h1)] <= (($signed(reg1599) ?
                          (reg1467 <= reg1534) : (reg1456 ^~ (8'ha3))) ?
                      reg1601[(5'h17):(4'hf)] : {(reg1670 ~^ (7'h48)),
                          (reg1662 ? reg1561 : reg1412)}))};
              reg1687 <= reg1446;
              reg1691 = $unsigned(reg1451);
            end
        end
      if (reg1683[(5'h10):(4'hc)])
        begin
          for (forvar1692 = (1'h0); (forvar1692 < (3'h6)); forvar1692 = (forvar1692 + (1'h1)))
            begin
              reg1693 = (((^~(reg1684[(4'h8):(3'h6)] >= (reg1642 ?
                      reg1677 : reg1411))) != reg1591) ?
                  reg1470 : (reg1689 ? wire1584 : (reg1623 << (~reg1675))));
              reg1694 = ($signed({reg1529,
                  ((~|(8'hba)) ?
                      reg1508[(4'ha):(3'h4)] : reg1516[(5'h1e):(5'h16)])}) + (-$signed($unsigned(reg1577))));
              reg1695 <= ((-$unsigned(($unsigned((8'ha7)) <= reg1568[(4'h9):(2'h3)]))) >> (-reg1600[(1'h1):(1'h1)]));
              reg1696 = reg1613[(3'h6):(3'h5)];
              reg1697 <= reg1504[(5'h17):(4'hc)];
              reg1698 <= reg1505[(3'h5):(2'h2)];
            end
          reg1699 = reg1661[(2'h3):(1'h0)];
          reg1700 <= ((~^(reg1682 >= (-(~reg1445)))) ?
              (^reg1619) : $signed((&$unsigned(reg1440[(3'h5):(3'h4)]))));
          for (forvar1701 = (1'h0); (forvar1701 < (2'h3)); forvar1701 = (forvar1701 + (1'h1)))
            begin
              reg1702 <= $unsigned(($unsigned(reg1385[(5'h10):(4'hb)]) > (~^$unsigned((7'h58)))));
              reg1703 = (8'ha4);
              reg1704 <= (!(($signed($unsigned((8'hbc))) ^~ {{reg1486},
                  (reg1684 >> reg1553),
                  (-reg1489)}) > $signed(reg1472)));
              reg1705 <= (8'ha6);
            end
        end
      else
        begin
          reg1692 = reg1604;
          for (forvar1693 = (1'h0); (forvar1693 < (3'h4)); forvar1693 = (forvar1693 + (1'h1)))
            begin
              reg1694 = reg1444[(5'h12):(4'h9)];
            end
          reg1696 = $signed((reg1550[(5'h10):(4'hb)] < (reg1556[(2'h3):(1'h1)] - $signed(((8'hac) ?
              reg1630 : (8'hab))))));
          reg1699 = (({((reg1565 ? reg1588 : reg1700) < $signed(reg1512))} ?
              {$signed((-reg1388)),
                  ((reg1590 >= (8'hab)) < (reg1489 ^~ reg1700))} : reg1575) || (reg1650[(1'h0):(1'h0)] ?
              (($unsigned(wire1668) & $unsigned(reg1531)) >>> $signed((reg1550 >> reg1592))) : $unsigned(((~|reg1547) ~^ $signed(reg1691)))));
        end
      for (forvar1706 = (1'h0); (forvar1706 < (1'h0)); forvar1706 = (forvar1706 + (1'h1)))
        begin
          for (forvar1707 = (1'h0); (forvar1707 < (1'h0)); forvar1707 = (forvar1707 + (1'h1)))
            begin
              reg1708 <= reg1393[(4'ha):(3'h7)];
              reg1709 <= $unsigned({reg1505,
                  {reg1705},
                  {{(wire1583 ? reg1593 : (8'haf))}, reg1465}});
              reg1710 <= reg1576[(1'h0):(1'h0)];
              reg1711 <= $signed(reg1385);
              reg1712 <= $unsigned(reg1671);
              reg1713 <= (-(&(((reg1453 ? reg1695 : reg1525) | (reg1619 ?
                      reg1572 : reg1547)) ?
                  $unsigned($unsigned((8'hba))) : reg1572[(1'h0):(1'h0)])));
              reg1714 <= reg1690[(3'h7):(3'h5)];
            end
          reg1715 <= {($unsigned(reg1507) ? reg1391 : (!reg1693))};
          reg1716 <= $unsigned((|$unsigned({{reg1516}})));
          if (reg1516[(3'h4):(3'h4)])
            begin
              reg1717 <= reg1593;
            end
          else
            begin
              reg1718 = reg1463;
            end
          reg1719 <= $unsigned($unsigned($signed($signed({reg1716,
              wire1647}))));
        end
      reg1720 <= (reg1663[(2'h2):(2'h2)] | (~((^(+(7'h4b))) ?
          (8'ha7) : reg1625[(3'h5):(3'h5)])));
      reg1721 <= $unsigned(wire1462[(1'h0):(1'h0)]);
      if ((~^(reg1697 ?
          reg1465[(1'h0):(1'h0)] : (reg1454 && ($signed((7'h4e)) ?
              $signed(reg1721) : $unsigned(reg1670))))))
        begin
          reg1722 = (&((&$unsigned((8'hb3))) | $signed({reg1619[(4'ha):(4'ha)],
              wire1422,
              (reg1626 || reg1479)})));
        end
      else
        begin
          reg1722 = (reg1699 > $signed({$signed((reg1568 >> reg1631)),
              $signed($signed(reg1430)),
              $signed((reg1703 ? reg1577 : reg1556))}));
          reg1723 = (&($signed((-(reg1710 - reg1676))) ?
              reg1662 : reg1658[(3'h6):(3'h6)]));
          for (forvar1724 = (1'h0); (forvar1724 < (3'h4)); forvar1724 = (forvar1724 + (1'h1)))
            begin
              reg1725 = reg1451;
              reg1726 <= reg1593;
            end
          for (forvar1727 = (1'h0); (forvar1727 < (1'h0)); forvar1727 = (forvar1727 + (1'h1)))
            begin
              reg1728 = $signed(reg1528[(5'h15):(4'hd)]);
              reg1729 = reg1670;
              reg1730 <= ((reg1690 <<< {{(reg1728 >> wire1462)},
                      (~reg1630[(4'hc):(4'h8)])}) ?
                  (7'h48) : reg1711);
              reg1731 = ((-{((reg1509 ? reg1720 : reg1445) * (~&reg1685)),
                      reg1606[(5'h11):(2'h3)]}) ?
                  (~^(~&(&$unsigned(reg1411)))) : reg1631[(5'h10):(3'h7)]);
              reg1732 <= reg1514;
            end
          reg1733 <= (~^(reg1624 ?
              ((reg1592[(1'h1):(1'h0)] || reg1481) ?
                  ($unsigned(forvar1701) ?
                      reg1718[(3'h7):(3'h7)] : $unsigned((7'h43))) : {((7'h48) + reg1658)}) : forvar1692));
          reg1734 <= $unsigned((!reg1565));
          for (forvar1735 = (1'h0); (forvar1735 < (3'h4)); forvar1735 = (forvar1735 + (1'h1)))
            begin
              reg1736 = reg1695;
              reg1737 = reg1430;
              reg1738 = (~reg1679);
              reg1739 <= (^~reg1391[(2'h2):(1'h1)]);
            end
        end
      reg1740 <= {(!$unsigned(reg1604)), (8'hb1)};
    end
  always
    @(posedge clk) begin
      for (forvar1741 = (1'h0); (forvar1741 < (2'h3)); forvar1741 = (forvar1741 + (1'h1)))
        begin
          reg1742 <= $unsigned($signed($signed(reg1708)));
          if (($unsigned(reg1524[(1'h1):(1'h0)]) <<< ((!$signed(reg1713[(3'h7):(2'h2)])) ?
              ((~&(reg1690 ?
                  reg1671 : reg1688)) - reg1606[(4'he):(4'h8)]) : reg1524[(3'h6):(2'h2)])))
            begin
              reg1743 <= reg1508[(4'hd):(1'h1)];
            end
          else
            begin
              reg1743 <= $unsigned(reg1582);
              reg1744 <= wire1381[(2'h3):(1'h0)];
              reg1745 = reg1637;
              reg1746 <= reg1700;
              reg1747 <= {reg1439[(4'he):(2'h3)]};
              reg1748 <= $signed(reg1463);
              reg1749 = (reg1623 ?
                  {(reg1712[(1'h1):(1'h1)] ?
                          ($signed(reg1458) == (reg1622 ?
                              reg1702 : (8'hb6))) : {(+reg1619)}),
                      $unsigned(reg1435[(4'ha):(2'h3)])} : ($unsigned(($signed(reg1688) <= reg1385[(3'h6):(2'h3)])) << (((reg1451 ?
                              reg1726 : reg1732) ?
                          (reg1550 ?
                              (8'hb6) : reg1681) : reg1595[(2'h2):(2'h2)]) ?
                      (reg1529[(4'hb):(3'h5)] << $unsigned(reg1414)) : (|(reg1573 ?
                          (7'h4e) : reg1577)))));
            end
          for (forvar1750 = (1'h0); (forvar1750 < (3'h4)); forvar1750 = (forvar1750 + (1'h1)))
            begin
              reg1751 = $signed(reg1545[(4'hc):(3'h7)]);
              reg1752 <= (!($unsigned(((reg1451 ? reg1515 : reg1644) ?
                  ((7'h53) ? wire1460 : reg1559) : (8'haa))) != reg1439));
            end
          for (forvar1753 = (1'h0); (forvar1753 < (2'h3)); forvar1753 = (forvar1753 + (1'h1)))
            begin
              reg1754 = reg1633[(4'hc):(3'h7)];
              reg1755 <= reg1563[(5'h10):(3'h5)];
            end
          reg1756 = ((({reg1512[(3'h5):(3'h4)], reg1556, $unsigned(reg1516)} ?
                  $unsigned($signed((7'h4e))) : $unsigned($unsigned(reg1430))) ?
              reg1716[(1'h1):(1'h0)] : (7'h44)) <= ((^((reg1748 ?
                  reg1520 : reg1734) ?
              (~^reg1531) : reg1702)) ^ (&reg1743)));
          reg1757 = reg1588;
          reg1758 <= ($unsigned({reg1745[(2'h3):(1'h0)],
              reg1650,
              $unsigned($signed(reg1622))}) & ($signed((reg1472[(1'h1):(1'h0)] & reg1493)) ?
              (reg1726 ?
                  reg1391[(4'ha):(3'h6)] : ({reg1550} ?
                      (forvar1753 * reg1415) : $unsigned(reg1642))) : reg1704[(4'ha):(3'h7)]));
        end
      reg1759 <= $signed($unsigned($unsigned(reg1708)));
    end
  assign wire1760 = (~&reg1397[(4'ha):(3'h6)]);
  assign wire1761 = ((|$unsigned($unsigned(reg1601[(2'h2):(1'h1)]))) ?
                        (((reg1568 > {reg1719, reg1582, reg1397}) != (reg1531 ?
                                reg1447[(5'h13):(4'hb)] : ((7'h4e) ?
                                    wire1462 : reg1576))) ?
                            reg1573 : reg1486) : wire1461[(5'h11):(4'he)]);
  assign wire1762 = reg1502;
  assign wire1763 = $unsigned(wire1761);
  assign wire1764 = reg1688[(3'h4):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar1765 = (1'h0); (forvar1765 < (3'h6)); forvar1765 = (forvar1765 + (1'h1)))
        begin
          reg1766 <= reg1673;
          reg1767 = (7'h4e);
          reg1768 = reg1447[(1'h1):(1'h1)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1059
#(parameter param1324 = (((+{((8'hb9) ? (7'h48) : (8'haf)), (^(8'ha7)), {(8'hb3)}}) ? ({((8'hb2) ? (8'ha9) : (8'ha8)), ((7'h41) ? (8'ha0) : (7'h41))} != (~^((8'hb5) ? (8'h9f) : (8'ha4)))) : ({((8'hba) ? (7'h57) : (8'h9e))} <<< (((8'hb7) <<< (7'h52)) <<< ((8'hab) ? (7'h47) : (8'ha9))))) ? ({(!(|(8'hba))), (7'h45), ((^(8'hbc)) & {(7'h52), (7'h57)})} << (7'h42)) : (!({((8'ha0) > (7'h47)), (~&(7'h4c)), ((8'ha7) ? (8'ha4) : (8'hb0))} ? (+(!(8'hae))) : (~|{(7'h4e), (7'h56)})))), 
parameter param1325 = (param1324 ~^ ((((^~param1324) | {(8'haf), param1324, param1324}) ? ((~^param1324) & (-param1324)) : (param1324 ? (^~param1324) : {(7'h46), param1324, (7'h4e)})) != (~^(~(~|param1324))))), 
parameter param1326 = (param1325 << (((+{param1324, (8'hbc), param1325}) > param1324) ? param1324 : ((~^(param1325 ? (7'h53) : param1324)) ? {{param1324, param1325, param1325}} : (-{param1324, param1324, param1325})))))
(y, clk, wire1064, wire1063, wire1062, wire1061, wire1060);
  output wire [(32'h1124):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire1064;
  input wire signed [(3'h7):(1'h0)] wire1063;
  input wire signed [(5'h12):(1'h0)] wire1062;
  input wire signed [(5'h15):(1'h0)] wire1061;
  input wire signed [(4'he):(1'h0)] wire1060;
  wire [(5'h19):(1'h0)] wire1217;
  wire [(4'he):(1'h0)] wire1216;
  wire signed [(5'h15):(1'h0)] wire1215;
  wire [(5'h15):(1'h0)] wire1195;
  wire signed [(2'h2):(1'h0)] wire1094;
  wire signed [(5'h11):(1'h0)] wire1065;
  reg [(2'h2):(1'h0)] reg1323 = (1'h0);
  reg [(5'h16):(1'h0)] reg1319 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1318 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1317 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1315 = (1'h0);
  reg [(4'he):(1'h0)] reg1314 = (1'h0);
  reg [(4'hb):(1'h0)] reg1313 = (1'h0);
  reg [(4'h9):(1'h0)] reg1308 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1307 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1304 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1301 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1300 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1298 = (1'h0);
  reg [(5'h12):(1'h0)] reg1294 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1293 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1291 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1289 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1285 = (1'h0);
  reg [(5'h19):(1'h0)] reg1282 = (1'h0);
  reg [(4'h9):(1'h0)] reg1278 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1272 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1268 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1267 = (1'h0);
  reg [(5'h13):(1'h0)] reg1265 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1262 = (1'h0);
  reg [(4'h9):(1'h0)] reg1261 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1259 = (1'h0);
  reg [(5'h13):(1'h0)] reg1257 = (1'h0);
  reg [(5'h12):(1'h0)] reg1256 = (1'h0);
  reg [(4'h8):(1'h0)] reg1254 = (1'h0);
  reg [(5'h14):(1'h0)] reg1250 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1248 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1247 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1246 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1241 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1239 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1238 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1237 = (1'h0);
  reg [(5'h12):(1'h0)] reg1235 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1233 = (1'h0);
  reg [(2'h3):(1'h0)] reg1231 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1229 = (1'h0);
  reg [(3'h6):(1'h0)] reg1228 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1226 = (1'h0);
  reg [(5'h19):(1'h0)] reg1221 = (1'h0);
  reg [(3'h5):(1'h0)] reg1213 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1210 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1209 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1207 = (1'h0);
  reg [(4'h9):(1'h0)] reg1206 = (1'h0);
  reg [(4'hf):(1'h0)] reg1204 = (1'h0);
  reg [(5'h15):(1'h0)] reg1202 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1200 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1199 = (1'h0);
  reg [(3'h7):(1'h0)] reg1198 = (1'h0);
  reg [(2'h3):(1'h0)] reg1192 = (1'h0);
  reg [(3'h5):(1'h0)] reg1191 = (1'h0);
  reg [(5'h12):(1'h0)] reg1187 = (1'h0);
  reg [(5'h18):(1'h0)] reg1186 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1185 = (1'h0);
  reg [(5'h11):(1'h0)] reg1183 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1178 = (1'h0);
  reg [(5'h18):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1174 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1169 = (1'h0);
  reg [(5'h19):(1'h0)] reg1167 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1163 = (1'h0);
  reg [(4'ha):(1'h0)] reg1162 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1161 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1158 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1155 = (1'h0);
  reg [(4'he):(1'h0)] reg1153 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1151 = (1'h0);
  reg [(3'h6):(1'h0)] reg1150 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1149 = (1'h0);
  reg [(5'h15):(1'h0)] reg1148 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1144 = (1'h0);
  reg [(4'hb):(1'h0)] reg1143 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1142 = (1'h0);
  reg [(4'hc):(1'h0)] reg1138 = (1'h0);
  reg [(5'h11):(1'h0)] reg1137 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1136 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1135 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1133 = (1'h0);
  reg [(5'h11):(1'h0)] reg1131 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1130 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1129 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1126 = (1'h0);
  reg [(5'h13):(1'h0)] reg1124 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1120 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1119 = (1'h0);
  reg [(5'h15):(1'h0)] reg1118 = (1'h0);
  reg [(4'hd):(1'h0)] reg1116 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1115 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1113 = (1'h0);
  reg [(2'h2):(1'h0)] reg1112 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1108 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1104 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1103 = (1'h0);
  reg [(3'h7):(1'h0)] reg1102 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1101 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1096 = (1'h0);
  reg [(4'hf):(1'h0)] reg1093 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1091 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1088 = (1'h0);
  reg [(3'h5):(1'h0)] reg1087 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1085 = (1'h0);
  reg [(4'hd):(1'h0)] reg1084 = (1'h0);
  reg [(5'h18):(1'h0)] reg1082 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1080 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1073 = (1'h0);
  reg [(4'h9):(1'h0)] reg1072 = (1'h0);
  reg [(4'hf):(1'h0)] reg1069 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1068 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1067 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1322 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1321 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1320 = (1'h0);
  reg [(5'h18):(1'h0)] reg1316 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1312 = (1'h0);
  reg [(5'h17):(1'h0)] reg1311 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1310 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1309 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1306 = (1'h0);
  reg [(4'hf):(1'h0)] reg1305 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1303 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1302 = (1'h0);
  reg [(3'h5):(1'h0)] reg1299 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1297 = (1'h0);
  reg [(4'hf):(1'h0)] reg1296 = (1'h0);
  reg [(3'h6):(1'h0)] reg1295 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1292 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1290 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1288 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1287 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1286 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1284 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1283 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1281 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1280 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1279 = (1'h0);
  reg [(3'h4):(1'h0)] reg1277 = (1'h0);
  reg [(5'h15):(1'h0)] reg1276 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1275 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1274 = (1'h0);
  reg [(5'h16):(1'h0)] reg1273 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1271 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1270 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1269 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1266 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1264 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1263 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1260 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1258 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1255 = (1'h0);
  reg [(4'h9):(1'h0)] reg1253 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1252 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1251 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1249 = (1'h0);
  reg [(5'h17):(1'h0)] reg1245 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1244 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1243 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1242 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1240 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1236 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1234 = (1'h0);
  reg [(5'h15):(1'h0)] reg1232 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1230 = (1'h0);
  reg [(3'h6):(1'h0)] reg1227 = (1'h0);
  reg [(4'hc):(1'h0)] reg1225 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1224 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1223 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1222 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1220 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1219 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1218 = (1'h0);
  reg [(4'he):(1'h0)] reg1214 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1212 = (1'h0);
  reg [(2'h2):(1'h0)] reg1211 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1208 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1205 = (1'h0);
  reg [(4'he):(1'h0)] reg1203 = (1'h0);
  reg [(5'h19):(1'h0)] reg1201 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1197 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1196 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1194 = (1'h0);
  reg [(5'h14):(1'h0)] reg1193 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1190 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1189 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1188 = (1'h0);
  reg [(4'hc):(1'h0)] reg1184 = (1'h0);
  reg [(4'h8):(1'h0)] reg1182 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1181 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1180 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1179 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1177 = (1'h0);
  reg [(5'h17):(1'h0)] reg1175 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1173 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1172 = (1'h0);
  reg [(4'hf):(1'h0)] reg1171 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1170 = (1'h0);
  reg [(4'hd):(1'h0)] reg1168 = (1'h0);
  reg [(2'h2):(1'h0)] reg1164 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1160 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1166 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1165 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1164 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1160 = (1'h0);
  reg [(2'h3):(1'h0)] reg1159 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1157 = (1'h0);
  reg [(3'h5):(1'h0)] reg1156 = (1'h0);
  reg [(3'h5):(1'h0)] reg1154 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1152 = (1'h0);
  reg [(5'h12):(1'h0)] reg1147 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1146 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1145 = (1'h0);
  reg [(3'h7):(1'h0)] reg1141 = (1'h0);
  reg [(3'h4):(1'h0)] reg1140 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1139 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1134 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar1131 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1132 = (1'h0);
  reg [(4'h9):(1'h0)] reg1128 = (1'h0);
  reg [(5'h14):(1'h0)] reg1127 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1125 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1123 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1122 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1121 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1117 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1114 = (1'h0);
  reg [(3'h5):(1'h0)] reg1107 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1099 = (1'h0);
  reg [(5'h16):(1'h0)] reg1111 = (1'h0);
  reg [(4'hd):(1'h0)] reg1110 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1109 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1107 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1106 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1105 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1100 = (1'h0);
  reg [(5'h18):(1'h0)] reg1099 = (1'h0);
  reg [(3'h4):(1'h0)] reg1098 = (1'h0);
  reg [(5'h14):(1'h0)] reg1097 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1095 = (1'h0);
  reg [(5'h18):(1'h0)] reg1092 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1090 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1089 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1086 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1083 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1081 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1079 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1078 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1077 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1076 = (1'h0);
  reg [(5'h16):(1'h0)] reg1075 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1074 = (1'h0);
  reg [(5'h15):(1'h0)] reg1071 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1070 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1066 = (1'h0);
  assign y = {wire1217,
                 wire1216,
                 wire1215,
                 wire1195,
                 wire1094,
                 wire1065,
                 reg1323,
                 reg1319,
                 reg1318,
                 reg1317,
                 reg1315,
                 reg1314,
                 reg1313,
                 reg1308,
                 reg1307,
                 reg1304,
                 reg1301,
                 reg1300,
                 reg1298,
                 reg1294,
                 reg1293,
                 reg1291,
                 reg1289,
                 reg1285,
                 reg1282,
                 reg1278,
                 reg1272,
                 reg1268,
                 reg1267,
                 reg1265,
                 reg1262,
                 reg1261,
                 reg1259,
                 reg1257,
                 reg1256,
                 reg1254,
                 reg1250,
                 reg1248,
                 reg1247,
                 reg1246,
                 reg1241,
                 reg1239,
                 reg1238,
                 reg1237,
                 reg1235,
                 reg1233,
                 reg1231,
                 reg1229,
                 reg1228,
                 reg1226,
                 reg1221,
                 reg1213,
                 reg1210,
                 reg1209,
                 reg1207,
                 reg1206,
                 reg1204,
                 reg1202,
                 reg1200,
                 reg1199,
                 reg1198,
                 reg1192,
                 reg1191,
                 reg1187,
                 reg1186,
                 reg1185,
                 reg1183,
                 reg1178,
                 reg1176,
                 reg1174,
                 reg1169,
                 reg1167,
                 reg1163,
                 reg1162,
                 reg1161,
                 reg1158,
                 reg1155,
                 reg1153,
                 reg1151,
                 reg1150,
                 reg1149,
                 reg1148,
                 reg1144,
                 reg1143,
                 reg1142,
                 reg1138,
                 reg1137,
                 reg1136,
                 reg1135,
                 reg1133,
                 reg1131,
                 reg1130,
                 reg1129,
                 reg1126,
                 reg1124,
                 reg1120,
                 reg1119,
                 reg1118,
                 reg1116,
                 reg1115,
                 reg1113,
                 reg1112,
                 reg1108,
                 reg1104,
                 reg1103,
                 reg1102,
                 reg1101,
                 reg1096,
                 reg1093,
                 reg1091,
                 reg1088,
                 reg1087,
                 reg1085,
                 reg1084,
                 reg1082,
                 reg1080,
                 reg1073,
                 reg1072,
                 reg1069,
                 reg1068,
                 reg1067,
                 reg1322,
                 reg1321,
                 reg1320,
                 reg1316,
                 reg1312,
                 reg1311,
                 reg1310,
                 reg1309,
                 forvar1306,
                 reg1305,
                 reg1303,
                 reg1302,
                 reg1299,
                 reg1297,
                 reg1296,
                 reg1295,
                 reg1292,
                 reg1290,
                 forvar1288,
                 forvar1287,
                 reg1286,
                 forvar1284,
                 reg1283,
                 forvar1281,
                 reg1280,
                 reg1279,
                 reg1277,
                 reg1276,
                 reg1275,
                 reg1274,
                 reg1273,
                 reg1271,
                 reg1270,
                 reg1269,
                 forvar1266,
                 forvar1264,
                 reg1263,
                 reg1260,
                 forvar1258,
                 reg1255,
                 reg1253,
                 reg1252,
                 reg1251,
                 reg1249,
                 reg1245,
                 reg1244,
                 reg1243,
                 reg1242,
                 reg1240,
                 reg1236,
                 reg1234,
                 reg1232,
                 reg1230,
                 reg1227,
                 reg1225,
                 forvar1224,
                 forvar1223,
                 reg1222,
                 reg1220,
                 forvar1219,
                 forvar1218,
                 reg1214,
                 forvar1212,
                 reg1211,
                 reg1208,
                 reg1205,
                 reg1203,
                 reg1201,
                 forvar1197,
                 forvar1196,
                 reg1194,
                 reg1193,
                 forvar1190,
                 reg1189,
                 reg1188,
                 reg1184,
                 reg1182,
                 forvar1181,
                 reg1180,
                 reg1179,
                 reg1177,
                 reg1175,
                 forvar1173,
                 reg1172,
                 reg1171,
                 reg1170,
                 reg1168,
                 reg1164,
                 reg1160,
                 reg1166,
                 reg1165,
                 forvar1164,
                 forvar1160,
                 reg1159,
                 reg1157,
                 reg1156,
                 reg1154,
                 reg1152,
                 reg1147,
                 reg1146,
                 reg1145,
                 reg1141,
                 reg1140,
                 reg1139,
                 reg1134,
                 forvar1131,
                 reg1132,
                 reg1128,
                 reg1127,
                 reg1125,
                 forvar1123,
                 reg1122,
                 reg1121,
                 forvar1117,
                 forvar1114,
                 reg1107,
                 forvar1099,
                 reg1111,
                 reg1110,
                 reg1109,
                 forvar1107,
                 reg1106,
                 reg1105,
                 reg1100,
                 reg1099,
                 reg1098,
                 reg1097,
                 forvar1095,
                 reg1092,
                 reg1090,
                 reg1089,
                 reg1086,
                 reg1083,
                 reg1081,
                 reg1079,
                 forvar1078,
                 forvar1077,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1071,
                 reg1070,
                 forvar1066,
                 (1'h0)};
  assign wire1065 = (&(^~(|(^~(wire1060 & wire1063)))));
  always
    @(posedge clk) begin
      for (forvar1066 = (1'h0); (forvar1066 < (3'h5)); forvar1066 = (forvar1066 + (1'h1)))
        begin
          reg1067 <= (~|wire1063[(3'h4):(3'h4)]);
          reg1068 <= (~|{($signed((wire1062 && forvar1066)) != $unsigned($signed((7'h41))))});
          reg1069 <= (+$unsigned(wire1062[(2'h2):(2'h2)]));
          reg1070 = (7'h41);
          if (forvar1066[(3'h6):(3'h6)])
            begin
              reg1071 = wire1063[(2'h2):(1'h0)];
              reg1072 <= reg1069;
              reg1073 <= wire1060;
              reg1074 = ((reg1073 ?
                  $unsigned($unsigned((reg1069 | wire1060))) : (7'h52)) * (^~reg1073[(4'h8):(3'h7)]));
            end
          else
            begin
              reg1072 <= ((^wire1065[(2'h3):(1'h1)]) ?
                  $unsigned(wire1063) : (~&{((wire1060 > wire1065) ?
                          $signed((8'hbb)) : (forvar1066 >> wire1061)),
                      $signed(reg1070[(5'h1a):(4'hb)])}));
            end
          reg1075 = (+{$unsigned(((reg1074 ?
                  reg1068 : forvar1066) && reg1067[(3'h7):(3'h5)])),
              $signed($signed((7'h45)))});
          reg1076 = reg1074;
        end
      for (forvar1077 = (1'h0); (forvar1077 < (3'h5)); forvar1077 = (forvar1077 + (1'h1)))
        begin
          for (forvar1078 = (1'h0); (forvar1078 < (3'h6)); forvar1078 = (forvar1078 + (1'h1)))
            begin
              reg1079 = $unsigned(((wire1065[(3'h4):(2'h3)] ?
                      (wire1064[(2'h3):(2'h2)] ?
                          (^~wire1065) : $unsigned(forvar1078)) : (8'h9c)) ?
                  (($signed(reg1067) ?
                      $unsigned(reg1073) : (-wire1064)) >>> {reg1073[(5'h10):(4'hb)],
                      forvar1066}) : {({reg1073, forvar1078} + (|reg1068)),
                      (&forvar1078[(2'h2):(2'h2)]),
                      (~((7'h48) ~^ (8'hba)))}));
              reg1080 <= wire1064;
              reg1081 = reg1068[(2'h2):(1'h0)];
              reg1082 <= ((((reg1067 > (reg1081 ?
                      wire1062 : reg1067)) ~^ ({forvar1066} != $signed(wire1064))) == reg1079[(4'hc):(2'h2)]) ?
                  reg1072[(2'h2):(2'h2)] : (forvar1078 ?
                      $signed(wire1061) : reg1072[(2'h2):(1'h1)]));
              reg1083 = $signed($unsigned((reg1072 ^ ($signed(reg1074) - reg1072))));
            end
          if ((8'h9e))
            begin
              reg1084 <= {wire1062, (~|reg1076)};
              reg1085 <= $unsigned($signed(reg1082[(5'h13):(5'h13)]));
            end
          else
            begin
              reg1086 = (wire1062 < {$unsigned(wire1061),
                  $unsigned($signed(((8'hb5) - (8'hb1))))});
              reg1087 <= (^~$signed(reg1080[(2'h2):(2'h2)]));
              reg1088 <= $unsigned(reg1083);
              reg1089 = reg1072;
              reg1090 = $unsigned(((7'h4f) >= {reg1073,
                  ((|reg1075) ? {reg1075} : {forvar1077})}));
              reg1091 <= ((~|(+reg1067)) ?
                  (!(+$unsigned((|wire1063)))) : reg1074);
              reg1092 = {($signed($signed(reg1073)) ?
                      {($unsigned(reg1074) << $unsigned(reg1075)),
                          {$unsigned(wire1062)},
                          ((8'ha9) ?
                              reg1069[(3'h4):(1'h1)] : $unsigned(reg1069))} : reg1073)};
            end
          reg1093 <= reg1088[(3'h4):(2'h3)];
        end
    end
  assign wire1094 = reg1072[(3'h6):(2'h3)];
  always
    @(posedge clk) begin
      for (forvar1095 = (1'h0); (forvar1095 < (2'h3)); forvar1095 = (forvar1095 + (1'h1)))
        begin
          reg1096 <= wire1060;
          reg1097 = $unsigned($signed((-(^~{(8'hbf), reg1085, reg1087}))));
          reg1098 = ({(8'hbe)} ?
              ($signed(reg1082[(4'h8):(3'h7)]) ?
                  $signed(wire1060) : {(reg1067[(4'hf):(3'h7)] >= (reg1082 ?
                          forvar1095 : reg1087)),
                      ((reg1069 & reg1067) < (forvar1095 ~^ reg1096)),
                      $signed((reg1067 < wire1060))}) : wire1060[(1'h1):(1'h0)]);
        end
      if ({wire1060[(3'h6):(2'h3)],
          $unsigned((reg1085[(2'h2):(1'h1)] >> reg1082[(1'h1):(1'h1)]))})
        begin
          if ($signed((-reg1067)))
            begin
              reg1099 = wire1094[(1'h1):(1'h1)];
              reg1100 = reg1096;
              reg1101 <= (reg1088 | (7'h44));
              reg1102 <= $unsigned(reg1098);
              reg1103 <= (~|($unsigned($unsigned($unsigned(wire1064))) ?
                  ((reg1082 & $unsigned(reg1102)) == ({(7'h56), wire1063} ?
                      $unsigned(reg1091) : reg1084)) : {(wire1094 ?
                          $unsigned(reg1099) : wire1063[(3'h5):(2'h3)]),
                      forvar1095[(3'h6):(3'h6)]}));
              reg1104 <= ($unsigned((({(8'h9e)} < (~|reg1082)) > (~(reg1098 ?
                      reg1098 : reg1084)))) ?
                  $unsigned($signed($signed(((7'h40) > (7'h46))))) : ($signed(((reg1100 <= wire1060) * $signed((7'h4b)))) + ($signed($signed(reg1103)) * $signed($signed((7'h50))))));
            end
          else
            begin
              reg1099 = ((^(7'h4a)) >>> (reg1073[(4'h8):(3'h6)] ^~ ($unsigned({reg1069}) ^~ reg1072[(2'h2):(1'h0)])));
              reg1101 <= $unsigned($signed(($signed(reg1085) <= ((forvar1095 ~^ reg1101) <<< $signed(wire1065)))));
              reg1102 <= (8'hb7);
              reg1103 <= (reg1073 ?
                  ({(8'hb5)} << (reg1099[(5'h13):(3'h6)] ?
                      $unsigned((wire1061 == reg1098)) : $unsigned($unsigned(reg1098)))) : {(((reg1067 << reg1103) ?
                              forvar1095[(4'hf):(2'h2)] : wire1094[(1'h1):(1'h1)]) ?
                          {{reg1080}, reg1067} : {$signed(reg1073),
                              $signed(reg1082),
                              (7'h4d)})});
              reg1105 = (~&reg1093[(3'h5):(2'h3)]);
              reg1106 = {(reg1099[(1'h1):(1'h1)] ?
                      $signed((7'h4b)) : ($unsigned($unsigned(reg1072)) && reg1104))};
            end
          for (forvar1107 = (1'h0); (forvar1107 < (3'h5)); forvar1107 = (forvar1107 + (1'h1)))
            begin
              reg1108 <= $signed((reg1093[(4'hf):(3'h5)] ?
                  (&$signed((reg1098 >>> reg1068))) : (8'hbb)));
              reg1109 = (((forvar1107 ?
                  ((8'ha4) < ((8'hbf) ~^ reg1101)) : (!forvar1107[(1'h1):(1'h1)])) > $signed(($signed((7'h50)) | (|reg1102)))) >>> (wire1094 != (~|(+$signed(reg1100)))));
              reg1110 = (reg1069 ?
                  (^~(~((reg1093 ? reg1098 : forvar1095) ?
                      (reg1099 ?
                          (8'ha0) : (8'hbd)) : wire1094))) : $signed(reg1096));
              reg1111 = (($signed({(reg1084 ? reg1097 : reg1104),
                      reg1087[(1'h0):(1'h0)]}) ?
                  $signed($unsigned((reg1087 ?
                      reg1096 : reg1105))) : wire1064) == wire1060);
            end
        end
      else
        begin
          for (forvar1099 = (1'h0); (forvar1099 < (3'h4)); forvar1099 = (forvar1099 + (1'h1)))
            begin
              reg1100 = reg1068[(2'h3):(1'h1)];
              reg1105 = (^~reg1096[(4'hb):(3'h6)]);
              reg1106 = $signed($signed({(reg1108 ^~ $signed(reg1111)),
                  ({reg1110} ^ (reg1109 ? wire1094 : wire1065))}));
              reg1107 = reg1088;
              reg1109 = reg1096[(4'hf):(4'hb)];
            end
          if ((7'h50))
            begin
              reg1110 = (((&reg1072[(3'h5):(1'h0)]) ?
                  $unsigned($signed(reg1098)) : {(~|$unsigned(reg1088)),
                      (~&reg1098),
                      {$unsigned(wire1060)}}) >= {(~$signed($unsigned(reg1073))),
                  (((reg1073 | wire1065) ?
                      forvar1095 : reg1100[(2'h3):(1'h1)]) || (~|(wire1061 ?
                      (7'h43) : reg1103)))});
              reg1111 = ((~reg1108) ?
                  (reg1068 ?
                      ($signed(reg1087) ?
                          (~|$unsigned(reg1106)) : $unsigned((forvar1099 < reg1110))) : (reg1082 << (wire1061[(5'h10):(3'h7)] ?
                          (wire1094 ?
                              reg1103 : reg1085) : (!reg1103)))) : wire1094);
              reg1112 <= ($unsigned((!$unsigned({wire1063}))) & (((7'h52) ?
                      (-reg1103) : (~^$signed(reg1073))) ?
                  {{$signed(reg1082), $signed(reg1084)},
                      reg1108,
                      reg1093} : {{(reg1072 ? reg1084 : reg1067),
                          $unsigned(reg1072),
                          reg1067},
                      $unsigned(reg1111),
                      (8'had)}));
            end
          else
            begin
              reg1112 <= (reg1069 ?
                  (~|$unsigned(($unsigned(reg1088) ?
                      (reg1088 ?
                          reg1096 : wire1061) : forvar1107[(2'h2):(1'h0)]))) : (({(^reg1096),
                          $signed(reg1112)} || reg1108[(3'h7):(3'h5)]) ?
                      reg1108[(3'h5):(3'h5)] : (reg1100 ?
                          (!$unsigned((8'hb8))) : forvar1107)));
              reg1113 <= reg1109;
            end
          for (forvar1114 = (1'h0); (forvar1114 < (1'h0)); forvar1114 = (forvar1114 + (1'h1)))
            begin
              reg1115 <= $unsigned($signed((~reg1097[(3'h6):(1'h0)])));
              reg1116 <= wire1061;
            end
          for (forvar1117 = (1'h0); (forvar1117 < (3'h5)); forvar1117 = (forvar1117 + (1'h1)))
            begin
              reg1118 <= ($unsigned($unsigned((reg1068[(2'h3):(2'h2)] - $signed(forvar1095)))) >>> $signed($signed((+{reg1087,
                  reg1091,
                  reg1085}))));
            end
          if (reg1100)
            begin
              reg1119 <= wire1060[(4'hb):(4'h8)];
              reg1120 <= $unsigned($signed((reg1087[(2'h2):(1'h0)] ^ (+((8'ha3) ~^ reg1082)))));
            end
          else
            begin
              reg1121 = ($signed($signed((|$unsigned(forvar1117)))) ?
                  $unsigned($signed((-{reg1072}))) : (wire1062[(2'h2):(2'h2)] ^ {(reg1111[(5'h10):(4'hb)] ~^ (|(8'hb8))),
                      $unsigned($unsigned(reg1096))}));
              reg1122 = (((wire1060[(4'h8):(4'h8)] <= (+(~&forvar1117))) >>> $signed(((forvar1114 ?
                  reg1085 : reg1118) >= $unsigned(reg1119)))) + ($unsigned($signed((reg1116 | reg1104))) ?
                  (wire1060[(4'ha):(1'h1)] ?
                      wire1061 : $unsigned((~|reg1069))) : (^($unsigned(reg1113) == (-(8'ha9))))));
            end
        end
      if (reg1108)
        begin
          for (forvar1123 = (1'h0); (forvar1123 < (1'h1)); forvar1123 = (forvar1123 + (1'h1)))
            begin
              reg1124 <= (reg1088[(2'h2):(2'h2)] ?
                  $signed($signed((7'h51))) : (($unsigned($signed(reg1099)) ?
                          $unsigned((+reg1106)) : (wire1065 && (^~(8'hbd)))) ?
                      (!($signed(reg1120) ?
                          $unsigned(reg1067) : (reg1100 > reg1106))) : (~&$unsigned(reg1116[(3'h4):(3'h4)]))));
              reg1125 = reg1105[(5'h14):(4'hc)];
            end
          if ((+{($unsigned((8'hb5)) * reg1113),
              (~&(~|(~|reg1098))),
              $unsigned((~&(reg1115 ? reg1103 : reg1113)))}))
            begin
              reg1126 <= wire1063;
              reg1127 = (((8'hae) ?
                      ($signed($unsigned(forvar1117)) == (8'ha2)) : reg1097[(3'h6):(3'h6)]) ?
                  $signed($unsigned(wire1063[(2'h2):(1'h0)])) : {{{(forvar1114 ?
                                  reg1102 : forvar1099),
                              (~|reg1106),
                              (reg1099 ? reg1096 : reg1103)},
                          {{reg1069}}},
                      (+$unsigned(reg1111)),
                      $signed({(~^reg1104)})});
              reg1128 = (forvar1123 ?
                  reg1069[(4'ha):(4'h8)] : (reg1116[(4'hc):(4'ha)] * $unsigned($signed($unsigned(reg1103)))));
              reg1129 <= {$unsigned((((reg1105 ? reg1087 : reg1069) ?
                          forvar1099[(3'h7):(2'h3)] : reg1098) ?
                      (!{forvar1099, reg1115}) : $unsigned($signed(reg1120)))),
                  $unsigned((!((reg1069 ? reg1103 : wire1060) ?
                      ((7'h57) | reg1072) : wire1094)))};
              reg1130 <= reg1127[(4'hc):(1'h1)];
              reg1131 <= ($unsigned((($unsigned(reg1128) - $unsigned((8'haa))) ^~ reg1109)) ?
                  reg1104[(1'h0):(1'h0)] : $unsigned(wire1064[(4'hf):(1'h0)]));
              reg1132 = $signed({{reg1068, reg1100[(2'h2):(1'h0)]},
                  reg1122[(2'h2):(1'h0)]});
            end
          else
            begin
              reg1126 <= $unsigned((~|reg1097[(3'h6):(1'h0)]));
              reg1129 <= reg1100[(5'h19):(3'h7)];
            end
        end
      else
        begin
          for (forvar1123 = (1'h0); (forvar1123 < (1'h0)); forvar1123 = (forvar1123 + (1'h1)))
            begin
              reg1125 = ((($signed((+reg1080)) & wire1064) ?
                  wire1064[(2'h3):(1'h0)] : ($signed(reg1093[(4'hf):(4'hb)]) >> ((wire1065 < (8'hb6)) << (+(8'h9d))))) > ($unsigned($unsigned((reg1121 * reg1125))) ~^ (|reg1115)));
              reg1126 <= ((~{((8'hbb) && {forvar1114, reg1096})}) > reg1080);
              reg1129 <= reg1103;
            end
          reg1130 <= $unsigned((((|reg1129) ?
              (~^(~wire1063)) : reg1115) < $unsigned((reg1118 ?
              wire1063 : {reg1132, (8'hbf)}))));
          for (forvar1131 = (1'h0); (forvar1131 < (3'h6)); forvar1131 = (forvar1131 + (1'h1)))
            begin
              reg1133 <= (wire1063[(2'h3):(2'h2)] <<< ((reg1120 <<< ($signed(wire1062) ?
                      (+(8'ha7)) : (reg1118 ? reg1068 : reg1119))) ?
                  reg1103 : forvar1131[(5'h14):(5'h13)]));
              reg1134 = (reg1120[(1'h0):(1'h0)] ?
                  wire1064 : ($signed((~&reg1093)) ?
                      forvar1114[(1'h1):(1'h1)] : (^~(~(reg1105 ?
                          reg1115 : forvar1131)))));
              reg1135 <= $unsigned(reg1098);
              reg1136 <= reg1112[(2'h2):(2'h2)];
              reg1137 <= (~reg1127);
            end
          if ((~^reg1122))
            begin
              reg1138 <= wire1061;
              reg1139 = reg1091[(5'h16):(5'h13)];
              reg1140 = $signed($unsigned($signed((reg1129 ?
                  $unsigned((7'h44)) : reg1088[(1'h0):(1'h0)]))));
              reg1141 = (reg1101[(5'h14):(5'h11)] ^~ (($signed({(8'hb3)}) ?
                      forvar1095[(3'h4):(1'h0)] : reg1130[(2'h2):(1'h1)]) ?
                  reg1109 : $unsigned((^~(~&forvar1114)))));
            end
          else
            begin
              reg1138 <= reg1111;
            end
          if ((~$signed(($unsigned((reg1085 | reg1085)) ~^ $unsigned((~^wire1094))))))
            begin
              reg1142 <= ($signed($signed($signed((~|(7'h40))))) ?
                  ($unsigned({reg1106[(1'h0):(1'h0)],
                      wire1063[(3'h7):(2'h2)],
                      (wire1061 <= reg1069)}) & $unsigned(($signed(reg1080) ?
                      $unsigned(reg1087) : reg1099))) : ($signed($signed((-reg1134))) && reg1080));
              reg1143 <= $signed((~&$unsigned($signed({reg1087}))));
              reg1144 <= reg1104[(3'h4):(1'h1)];
              reg1145 = $signed(((forvar1114 - wire1094) ?
                  $signed(reg1122[(3'h6):(2'h2)]) : (~&(^~(reg1106 - (8'hb6))))));
            end
          else
            begin
              reg1142 <= $signed($signed($unsigned((^$unsigned(reg1129)))));
              reg1143 <= (((reg1087 ?
                  reg1121 : ($signed((8'hb5)) ?
                      (&(7'h57)) : (forvar1095 || wire1061))) ~^ $unsigned((reg1121 - forvar1123))) | ((~(-$signed(reg1110))) >>> (8'hb1)));
              reg1145 = $unsigned(reg1119[(1'h0):(1'h0)]);
              reg1146 = $unsigned(($unsigned($unsigned(forvar1123[(2'h2):(1'h0)])) <<< $unsigned($unsigned(reg1129))));
              reg1147 = wire1061[(4'hb):(1'h0)];
              reg1148 <= (reg1146 - ({reg1091[(5'h16):(5'h10)],
                      {(reg1084 >>> reg1106)}} ?
                  $signed(reg1072) : (+($unsigned(reg1099) ?
                      (&reg1126) : (reg1093 ? reg1098 : (7'h53))))));
              reg1149 <= reg1128[(2'h3):(2'h3)];
            end
        end
      if ((8'hbc))
        begin
          reg1150 <= $signed(($signed(reg1126[(3'h6):(1'h0)]) ?
              {(^~(&reg1106)), (~|{reg1121})} : $signed(reg1147)));
          reg1151 <= $unsigned(reg1096);
          if ($signed(((reg1108 + reg1107) ?
              (($signed(reg1111) ?
                  $unsigned(reg1150) : $unsigned(forvar1107)) >> reg1131[(4'hf):(3'h6)]) : reg1140)))
            begin
              reg1152 = {(|(wire1062[(2'h2):(1'h1)] ?
                      ((forvar1107 ?
                          reg1133 : reg1127) <<< $unsigned(reg1098)) : $signed(reg1107)))};
              reg1153 <= (7'h42);
              reg1154 = forvar1107;
              reg1155 <= $unsigned((^~$signed({(~^reg1115)})));
              reg1156 = reg1135;
            end
          else
            begin
              reg1152 = (^~(+$unsigned((^~(^~reg1116)))));
              reg1154 = ((8'h9f) ?
                  ((reg1139[(2'h3):(1'h0)] >>> wire1094[(1'h0):(1'h0)]) ?
                      (+(8'hba)) : (($unsigned(wire1094) >= (reg1098 >= reg1115)) ?
                          $signed(reg1124) : ($signed((7'h41)) ?
                              (reg1102 ?
                                  (7'h50) : reg1152) : $unsigned(reg1137)))) : reg1119);
              reg1156 = $unsigned(reg1127[(5'h13):(1'h0)]);
              reg1157 = $signed($signed((reg1115[(4'h9):(3'h6)] ^~ ($unsigned(reg1141) << (^reg1072)))));
            end
          reg1158 <= (~reg1148);
          reg1159 = forvar1095[(5'h10):(4'hd)];
          for (forvar1160 = (1'h0); (forvar1160 < (1'h0)); forvar1160 = (forvar1160 + (1'h1)))
            begin
              reg1161 <= $signed($unsigned(reg1146));
              reg1162 <= $unsigned((reg1149 < (^~reg1135)));
              reg1163 <= $signed((-forvar1123[(4'hd):(4'h9)]));
            end
          for (forvar1164 = (1'h0); (forvar1164 < (3'h5)); forvar1164 = (forvar1164 + (1'h1)))
            begin
              reg1165 = (reg1158 ? $signed(reg1156) : reg1153);
              reg1166 = (8'hae);
            end
        end
      else
        begin
          if ($unsigned(reg1139[(2'h2):(1'h0)]))
            begin
              reg1152 = reg1136[(1'h1):(1'h1)];
              reg1154 = forvar1099;
              reg1155 <= {$signed($signed(reg1154[(2'h2):(2'h2)])),
                  $unsigned($signed($unsigned((forvar1164 ?
                      reg1125 : reg1093)))),
                  $signed(({{(8'hb9), (7'h57), (8'ha3)},
                      (&reg1103),
                      (reg1146 >= reg1162)} ^ wire1061))};
              reg1156 = reg1131[(2'h2):(1'h1)];
            end
          else
            begin
              reg1150 <= $unsigned(wire1062[(2'h3):(2'h3)]);
              reg1152 = ($signed(wire1060) ?
                  reg1096[(5'h18):(3'h5)] : (^reg1124[(1'h1):(1'h0)]));
              reg1154 = $signed($signed(reg1132));
            end
          if ($unsigned((!wire1060[(1'h0):(1'h0)])))
            begin
              reg1157 = $unsigned($unsigned(((reg1129 ?
                  reg1132[(3'h7):(3'h5)] : ((7'h41) ?
                      (8'ha7) : reg1158)) ^~ $unsigned($signed(reg1125)))));
              reg1158 <= $signed(reg1136);
              reg1159 = reg1140[(2'h2):(2'h2)];
              reg1160 = (((8'hbc) ?
                      (|({(8'hb6), reg1093, reg1099} ?
                          (-wire1061) : (~&reg1128))) : $unsigned(((reg1151 ?
                          reg1163 : reg1115) * $unsigned(reg1073)))) ?
                  $unsigned({wire1065[(5'h11):(4'hb)]}) : ($unsigned(($unsigned(forvar1123) >> (reg1118 ^~ forvar1117))) ?
                      $unsigned((reg1135[(5'h19):(4'hc)] ?
                          (reg1150 ?
                              reg1122 : reg1115) : reg1139[(1'h1):(1'h1)])) : reg1161[(1'h1):(1'h1)]));
              reg1161 <= $signed($unsigned($signed($unsigned($signed(reg1154)))));
              reg1164 = $unsigned(($signed((~&reg1116[(3'h4):(2'h2)])) ?
                  {$signed($signed(reg1105))} : forvar1160));
            end
          else
            begin
              reg1158 <= (+(+reg1154));
              reg1161 <= (reg1160 ?
                  $unsigned($signed(reg1120)) : $unsigned($unsigned(reg1093[(4'h8):(2'h3)])));
              reg1162 <= $signed(((reg1091[(4'hd):(4'hd)] >> (~^reg1164[(2'h2):(1'h1)])) ?
                  $signed(forvar1114[(1'h0):(1'h0)]) : $signed(reg1084[(3'h7):(2'h2)])));
              reg1164 = {$unsigned(($unsigned((~(8'hab))) ?
                      (8'haf) : (&reg1073[(5'h18):(5'h16)])))};
              reg1167 <= $unsigned(reg1146);
            end
          if ($unsigned((reg1133[(4'h9):(3'h5)] ?
              ((+{reg1159, forvar1117}) ?
                  {reg1121[(4'ha):(4'h9)],
                      (reg1132 << reg1108),
                      (reg1129 <= forvar1114)} : reg1152[(5'h11):(2'h2)]) : {(reg1130 >>> (^~(8'haa))),
                  {reg1105[(1'h1):(1'h1)]},
                  $signed(reg1098)})))
            begin
              reg1168 = reg1072[(1'h0):(1'h0)];
              reg1169 <= $unsigned(reg1138);
            end
          else
            begin
              reg1168 = (8'ha4);
              reg1170 = $unsigned($signed(({((7'h4a) ^~ reg1113),
                      (^reg1115),
                      (+reg1080)} ?
                  (8'hae) : reg1102[(1'h0):(1'h0)])));
              reg1171 = (forvar1123[(4'he):(3'h5)] & $signed(((~reg1108[(4'ha):(1'h0)]) & $unsigned((-reg1143)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg1172 = $signed((^wire1061));
      if (($signed((({wire1065, reg1161, reg1068} ?
          $signed(reg1126) : reg1150[(2'h2):(1'h1)]) < $unsigned($signed(reg1119)))) | (!wire1062)))
        begin
          for (forvar1173 = (1'h0); (forvar1173 < (3'h6)); forvar1173 = (forvar1173 + (1'h1)))
            begin
              reg1174 <= (reg1137[(2'h2):(1'h0)] << ((((wire1064 | reg1150) & $unsigned(wire1061)) ?
                  reg1151[(1'h1):(1'h1)] : $signed((reg1151 != (8'h9e)))) * $signed($signed(forvar1173[(5'h10):(3'h5)]))));
              reg1175 = $unsigned(reg1082);
            end
          if ((8'hb5))
            begin
              reg1176 <= ({($unsigned($unsigned(reg1172)) && (!(reg1113 >>> reg1133)))} || $signed(reg1155));
            end
          else
            begin
              reg1176 <= $unsigned(reg1137[(2'h3):(1'h0)]);
              reg1177 = wire1062;
              reg1178 <= reg1129;
              reg1179 = {({(reg1101[(4'hc):(2'h2)] ?
                          (8'hb2) : $signed(reg1149)),
                      (((8'hab) ?
                          reg1169 : reg1175) * reg1144)} <= reg1085[(3'h7):(3'h7)]),
                  wire1094[(1'h0):(1'h0)],
                  $signed($signed($signed(((8'hab) && reg1176))))};
            end
        end
      else
        begin
          for (forvar1173 = (1'h0); (forvar1173 < (3'h6)); forvar1173 = (forvar1173 + (1'h1)))
            begin
              reg1174 <= (^$signed(((reg1158 ?
                      (reg1119 ? (7'h40) : reg1082) : ((7'h48) << reg1093)) ?
                  (+(reg1178 ~^ (8'hbd))) : $signed((reg1113 ?
                      (7'h51) : reg1142)))));
              reg1176 <= (-reg1148[(3'h7):(3'h4)]);
              reg1177 = reg1103;
              reg1179 = $signed(reg1169);
              reg1180 = $unsigned($unsigned(reg1129));
            end
          for (forvar1181 = (1'h0); (forvar1181 < (3'h6)); forvar1181 = (forvar1181 + (1'h1)))
            begin
              reg1182 = ({(+(8'hbe)),
                      ((~&$unsigned(reg1124)) ?
                          (8'ha1) : ($signed((7'h43)) ?
                              ((7'h53) >> reg1135) : reg1178))} ?
                  $unsigned($unsigned((reg1150[(3'h4):(1'h1)] ?
                      $unsigned(reg1084) : (reg1101 ~^ reg1158)))) : reg1144[(4'hf):(4'ha)]);
              reg1183 <= (+($unsigned($signed({(8'hbc), reg1178, reg1161})) ?
                  {reg1174[(4'hf):(2'h2)]} : $unsigned((~|reg1102[(3'h5):(1'h0)]))));
              reg1184 = ((({((7'h4c) <<< reg1151),
                          (reg1169 ~^ reg1183),
                          $signed(reg1138)} ^~ (!$signed(reg1088))) ?
                      reg1178 : ((^~$signed((8'hb6))) ?
                          reg1115 : (reg1161 ?
                              (reg1169 + reg1183) : $signed(reg1120)))) ?
                  (~^$unsigned((8'h9e))) : (+$signed(((reg1118 ?
                          reg1137 : reg1149) ?
                      reg1175 : (forvar1173 ? reg1177 : wire1063)))));
              reg1185 <= (8'hb3);
              reg1186 <= reg1155[(5'h16):(5'h16)];
              reg1187 <= $signed((~^{reg1161[(5'h11):(3'h7)],
                  $unsigned($unsigned((8'hbc)))}));
              reg1188 = reg1182;
            end
          reg1189 = ((~&$signed((^~reg1150))) >> (^~reg1068[(3'h5):(2'h3)]));
          for (forvar1190 = (1'h0); (forvar1190 < (3'h6)); forvar1190 = (forvar1190 + (1'h1)))
            begin
              reg1191 <= $signed(reg1187[(1'h0):(1'h0)]);
              reg1192 <= (reg1087[(3'h4):(1'h0)] ?
                  $unsigned(reg1167[(5'h19):(5'h19)]) : ($unsigned($unsigned((reg1073 ?
                          reg1176 : forvar1173))) ?
                      reg1096[(5'h1a):(4'hd)] : reg1151));
              reg1193 = reg1174;
            end
        end
      reg1194 = $unsigned($unsigned($signed($unsigned($signed(reg1085)))));
    end
  assign wire1195 = {$signed($unsigned(((reg1167 + reg1113) * wire1065))),
                        (($unsigned(reg1155) ?
                                {{reg1118, (7'h53), (8'ha5)},
                                    reg1072,
                                    (~^wire1061)} : reg1102[(2'h2):(1'h0)]) ?
                            $signed(reg1131[(4'hb):(1'h0)]) : (&$signed(reg1191[(3'h4):(3'h4)])))};
  always
    @(posedge clk) begin
      for (forvar1196 = (1'h0); (forvar1196 < (2'h2)); forvar1196 = (forvar1196 + (1'h1)))
        begin
          for (forvar1197 = (1'h0); (forvar1197 < (1'h0)); forvar1197 = (forvar1197 + (1'h1)))
            begin
              reg1198 <= reg1104[(1'h0):(1'h0)];
              reg1199 <= reg1091;
              reg1200 <= (|($unsigned((~&(reg1116 != (8'ha4)))) ?
                  (~&(^~reg1126)) : $signed(reg1158[(1'h0):(1'h0)])));
              reg1201 = $unsigned((reg1120 != (~^((~reg1069) ?
                  reg1093[(2'h3):(2'h3)] : (reg1136 < (7'h4b))))));
              reg1202 <= ((&(!((~(8'ha5)) <= {reg1108, reg1072, reg1072}))) ?
                  reg1133[(1'h1):(1'h0)] : reg1104[(3'h5):(3'h4)]);
              reg1203 = reg1112;
              reg1204 <= (~((reg1191[(3'h4):(1'h0)] ?
                  ((&reg1102) ?
                      $signed(reg1118) : $unsigned(reg1142)) : $signed((^~(8'ha1)))) >= (&(8'haa))));
            end
          reg1205 = $signed(reg1088);
        end
      reg1206 <= $unsigned(($signed(reg1198[(3'h6):(3'h4)]) ?
          (({reg1169, reg1203, (7'h46)} ?
                  reg1202[(5'h10):(4'hb)] : $unsigned(reg1167)) ?
              $unsigned($unsigned(reg1137)) : ((~reg1103) ?
                  $signed((8'hbc)) : (wire1195 >> reg1085))) : reg1091[(3'h4):(2'h3)]));
      reg1207 <= $unsigned(reg1069);
      reg1208 = $signed((~&((~|(~^wire1094)) ?
          reg1130 : $unsigned($unsigned(reg1082)))));
      reg1209 <= reg1204[(3'h5):(2'h3)];
      reg1210 <= (-$signed(reg1126));
      if ((^~($signed($signed({reg1143, reg1108})) ^~ (7'h58))))
        begin
          reg1211 = (~wire1094[(1'h1):(1'h1)]);
          for (forvar1212 = (1'h0); (forvar1212 < (2'h2)); forvar1212 = (forvar1212 + (1'h1)))
            begin
              reg1213 <= reg1136;
              reg1214 = ($unsigned($signed($signed((7'h48)))) ?
                  reg1199 : ($unsigned(({reg1207, reg1155} ?
                      ((8'hbe) <= reg1072) : (~&reg1131))) ^ reg1150[(2'h3):(1'h1)]));
            end
        end
      else
        begin
          reg1211 = (reg1136[(1'h1):(1'h0)] && $unsigned($signed(reg1068[(3'h7):(3'h6)])));
        end
    end
  assign wire1215 = ((~|reg1169) | reg1120[(4'ha):(3'h4)]);
  assign wire1216 = $signed($unsigned($signed($signed((~&(7'h54))))));
  assign wire1217 = reg1148[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar1218 = (1'h0); (forvar1218 < (3'h5)); forvar1218 = (forvar1218 + (1'h1)))
        begin
          for (forvar1219 = (1'h0); (forvar1219 < (3'h4)); forvar1219 = (forvar1219 + (1'h1)))
            begin
              reg1220 = reg1096[(5'h11):(4'hf)];
              reg1221 <= $signed(reg1135);
              reg1222 = (((wire1063 > reg1104) <= (reg1213 ?
                      (8'hb0) : ((reg1108 ?
                          wire1062 : reg1185) != (reg1202 << reg1084)))) ?
                  $unsigned((~|(~^{reg1144, reg1150, reg1221}))) : reg1183);
            end
        end
      for (forvar1223 = (1'h0); (forvar1223 < (1'h0)); forvar1223 = (forvar1223 + (1'h1)))
        begin
          for (forvar1224 = (1'h0); (forvar1224 < (2'h2)); forvar1224 = (forvar1224 + (1'h1)))
            begin
              reg1225 = $unsigned(reg1082);
              reg1226 <= (~reg1178[(3'h4):(2'h2)]);
              reg1227 = {$signed($signed((^$signed(reg1176))))};
              reg1228 <= (~|(~|reg1113[(2'h3):(2'h3)]));
              reg1229 <= wire1094;
            end
          reg1230 = ((~^{reg1138[(3'h6):(2'h3)]}) ?
              {reg1209[(4'ha):(4'h9)],
                  reg1207[(4'hc):(3'h5)],
                  (~$unsigned($unsigned(reg1202)))} : reg1161[(5'h16):(4'h8)]);
          reg1231 <= ($signed($signed({$unsigned(reg1101),
                  (reg1149 ^~ wire1063)})) ?
              $unsigned(((+$signed(wire1061)) == reg1186[(5'h11):(3'h5)])) : (7'h58));
          reg1232 = $signed(({(reg1225[(1'h1):(1'h0)] ^ $unsigned((7'h46))),
              $unsigned($unsigned(reg1191)),
              {(|reg1221), reg1204[(2'h2):(2'h2)]}} >>> ($unsigned((reg1163 ?
                  reg1210 : (7'h40))) ?
              ((~^wire1062) ?
                  $signed((8'hbf)) : $unsigned(wire1062)) : reg1082[(1'h0):(1'h0)])));
          reg1233 <= (reg1120[(1'h0):(1'h0)] ?
              (7'h51) : reg1131[(4'hd):(4'h8)]);
          reg1234 = reg1073[(5'h1a):(3'h7)];
        end
      if (reg1135[(2'h3):(2'h2)])
        begin
          if (reg1191[(2'h2):(1'h1)])
            begin
              reg1235 <= (^~$unsigned($unsigned((reg1230[(1'h0):(1'h0)] ^ $unsigned(reg1209)))));
              reg1236 = reg1199;
              reg1237 <= reg1080[(5'h10):(4'he)];
              reg1238 <= $signed(((|reg1131) ? $unsigned(reg1082) : reg1119));
              reg1239 <= (reg1084[(4'hd):(1'h1)] ?
                  ($signed(({reg1185} ?
                      {(7'h4c)} : (~reg1131))) && reg1174) : (~|{$unsigned($unsigned(reg1153)),
                      reg1200[(4'ha):(1'h0)],
                      ((reg1142 ? reg1234 : reg1144) ?
                          {reg1226, reg1237, reg1213} : {reg1202,
                              reg1155,
                              reg1238})}));
              reg1240 = ($signed(reg1151[(2'h3):(2'h2)]) == $unsigned($signed($signed($unsigned(reg1210)))));
              reg1241 <= reg1239;
            end
          else
            begin
              reg1236 = (~reg1131);
              reg1237 <= ((~|reg1167[(4'h9):(3'h6)]) != {(wire1062[(4'h9):(3'h7)] && reg1080),
                  $signed({wire1063, reg1232[(2'h3):(2'h2)]}),
                  $signed($unsigned((&reg1209)))});
              reg1238 <= (((^~$signed(reg1158[(5'h15):(5'h10)])) ^~ $signed(reg1101[(4'ha):(3'h7)])) * (reg1102 && $signed(($unsigned((7'h54)) ?
                  $signed(reg1135) : (reg1176 || wire1216)))));
              reg1240 = {($signed((reg1113 ?
                      (reg1136 ? reg1176 : reg1176) : (~reg1129))) == reg1187)};
              reg1242 = wire1062[(4'hc):(1'h0)];
            end
          if (($unsigned($signed((reg1183[(5'h10):(3'h6)] ?
                  (reg1192 ? reg1227 : reg1191) : (~&reg1206)))) ?
              $signed((~|$signed((^~reg1239)))) : (($signed($unsigned(reg1103)) ?
                  reg1206[(2'h2):(2'h2)] : ((reg1234 ? reg1088 : wire1215) ?
                      $unsigned(reg1135) : reg1129[(5'h12):(4'ha)])) > reg1151[(2'h2):(2'h2)])))
            begin
              reg1243 = wire1065[(4'hb):(1'h0)];
              reg1244 = wire1060;
              reg1245 = (&(reg1232[(4'hc):(4'h8)] ?
                  $unsigned($unsigned((-reg1151))) : (($signed(forvar1223) < $signed(reg1227)) ?
                      ((!reg1088) ?
                          $unsigned(reg1136) : reg1235[(3'h5):(3'h5)]) : ((reg1186 | (8'ha8)) * (^reg1232)))));
              reg1246 <= {(forvar1219 ?
                      (!(~^(wire1094 > (8'ha6)))) : (!$unsigned((7'h46)))),
                  (reg1093 || ($unsigned((reg1220 <= (8'hb4))) ?
                      ($unsigned(reg1087) ?
                          $signed(reg1067) : ((7'h48) + reg1150)) : {{reg1069,
                              reg1080},
                          reg1133}))};
              reg1247 <= reg1240;
              reg1248 <= wire1195[(3'h4):(1'h0)];
            end
          else
            begin
              reg1243 = reg1135;
              reg1246 <= ($signed(($signed((forvar1224 ?
                  reg1238 : reg1198)) << $unsigned({reg1246}))) > $signed(reg1112));
            end
        end
      else
        begin
          if ($unsigned((~({(forvar1223 <= reg1248), reg1153[(1'h0):(1'h0)]} ?
              reg1200[(4'hd):(1'h1)] : reg1135))))
            begin
              reg1235 <= reg1192[(1'h1):(1'h1)];
              reg1236 = ($unsigned(($signed($signed(reg1210)) ?
                  (8'ha4) : reg1234)) <= ((~&$unsigned(reg1221)) || reg1247));
              reg1240 = reg1115;
              reg1241 <= {reg1229[(4'he):(2'h2)]};
            end
          else
            begin
              reg1236 = reg1088;
              reg1240 = (8'ha5);
              reg1241 <= $signed((&reg1158[(2'h3):(1'h0)]));
              reg1242 = (reg1243 ?
                  (reg1187 ?
                      (~reg1246[(4'h9):(3'h6)]) : {reg1148,
                          (~&((7'h4f) ? reg1143 : reg1206))}) : wire1065);
              reg1243 = wire1062;
              reg1246 <= (~|$signed(reg1227));
              reg1249 = ((8'ha0) == reg1183[(3'h7):(3'h5)]);
            end
          if ((&{$signed(((reg1233 ? reg1102 : reg1240) ?
                  (~^reg1118) : wire1062[(4'hc):(4'ha)])),
              $unsigned($signed($unsigned((7'h44))))}))
            begin
              reg1250 <= ((($unsigned(((7'h41) ?
                          wire1216 : reg1161)) && (~(~|reg1091))) ?
                      (|reg1233) : $unsigned($unsigned((reg1116 ?
                          (7'h40) : reg1206)))) ?
                  $unsigned((reg1126[(4'h8):(2'h2)] >>> (reg1206 >> (wire1217 ?
                      reg1149 : reg1150)))) : wire1216[(3'h6):(1'h1)]);
              reg1251 = (7'h4c);
              reg1252 = ((7'h44) | (^$signed(reg1207)));
              reg1253 = (8'hb8);
              reg1254 <= $unsigned((reg1068 ?
                  (!((reg1085 >> reg1236) ^ reg1202)) : (~|$unsigned($unsigned(reg1116)))));
              reg1255 = {reg1144,
                  (((8'ha3) ?
                      {{reg1116}} : (reg1207[(3'h6):(1'h0)] >>> {reg1198,
                          wire1065})) >> reg1103[(4'hd):(4'h9)]),
                  reg1230};
              reg1256 <= (($unsigned(reg1242[(3'h6):(3'h5)]) ^ ((!reg1178) ?
                  (!$signed(wire1065)) : (((8'hb1) ? reg1124 : reg1252) ?
                      $unsigned((7'h45)) : (reg1118 ?
                          reg1119 : reg1101)))) << (!$signed(wire1217)));
            end
          else
            begin
              reg1251 = (~&(reg1112[(1'h1):(1'h0)] ?
                  (7'h49) : $signed(($unsigned(wire1065) ?
                      reg1167 : $signed(reg1238)))));
              reg1254 <= ($unsigned(reg1167) ?
                  {$signed(((!(7'h45)) ?
                          (reg1115 ?
                              reg1178 : reg1234) : (reg1120 != (7'h45))))} : $unsigned($unsigned(reg1162[(4'h8):(3'h6)])));
              reg1256 <= reg1246[(1'h1):(1'h0)];
              reg1257 <= $unsigned((((~&$signed(reg1239)) ?
                      $unsigned((reg1133 ?
                          (8'ha0) : reg1149)) : (~&$unsigned(wire1094))) ?
                  wire1094[(2'h2):(1'h1)] : reg1088));
            end
          for (forvar1258 = (1'h0); (forvar1258 < (3'h4)); forvar1258 = (forvar1258 + (1'h1)))
            begin
              reg1259 <= ((^~(reg1118 - (^~reg1129))) ?
                  {(-$unsigned(reg1169[(1'h1):(1'h0)])),
                      (($unsigned((8'hb1)) <= reg1226) ?
                          {(+reg1158),
                              (wire1065 != (8'hb8))} : wire1094)} : ((8'hac) ?
                      $unsigned(($signed(reg1096) ?
                          $signed(reg1243) : reg1073[(3'h5):(3'h4)])) : ((^$unsigned(reg1200)) && $signed(reg1225[(2'h2):(1'h1)]))));
              reg1260 = wire1215[(2'h2):(1'h1)];
              reg1261 <= $unsigned(reg1229[(5'h1b):(3'h4)]);
              reg1262 <= ($signed($unsigned(reg1131[(4'hf):(4'hd)])) ?
                  $signed(reg1072) : $signed($signed($unsigned({reg1256}))));
            end
          reg1263 = $signed(reg1115[(1'h1):(1'h0)]);
        end
      for (forvar1264 = (1'h0); (forvar1264 < (1'h0)); forvar1264 = (forvar1264 + (1'h1)))
        begin
          reg1265 <= (reg1263 ^~ reg1237[(2'h2):(2'h2)]);
          for (forvar1266 = (1'h0); (forvar1266 < (1'h1)); forvar1266 = (forvar1266 + (1'h1)))
            begin
              reg1267 <= (~&(reg1235 ?
                  $unsigned({(reg1248 < reg1226),
                      reg1209}) : ($unsigned($unsigned(reg1245)) ?
                      (8'ha7) : {(reg1200 ? reg1253 : reg1096),
                          $unsigned(reg1227)})));
              reg1268 <= $unsigned((reg1252[(4'hf):(2'h2)] >> (reg1253[(3'h5):(1'h1)] ^ ((reg1229 ?
                  reg1120 : reg1148) & $signed(reg1260)))));
              reg1269 = $unsigned(reg1256[(4'hc):(3'h5)]);
              reg1270 = ({reg1235[(4'hd):(3'h5)],
                      $signed(((forvar1223 >> wire1062) <= reg1144)),
                      $unsigned(((|reg1232) ? reg1112 : (reg1080 ^ reg1149)))} ?
                  (~^$signed($unsigned((reg1228 ?
                      (7'h43) : reg1072)))) : reg1222[(3'h5):(2'h2)]);
              reg1271 = $signed(((&reg1232[(5'h11):(4'h8)]) ?
                  ($unsigned((reg1202 ?
                      reg1254 : reg1198)) > ((reg1148 < reg1227) == $unsigned(reg1150))) : ($unsigned(reg1256) && (|{forvar1224,
                      (8'hbb),
                      reg1247}))));
              reg1272 <= (~^$signed((^$unsigned((forvar1264 << reg1142)))));
            end
          if ($signed(reg1242[(3'h4):(1'h0)]))
            begin
              reg1273 = reg1103[(5'h11):(4'he)];
            end
          else
            begin
              reg1273 = reg1103;
              reg1274 = $signed((7'h58));
            end
          if ((~^$unsigned(($unsigned($signed(reg1254)) ?
              wire1217[(5'h12):(3'h4)] : $signed(reg1227[(1'h0):(1'h0)])))))
            begin
              reg1275 = {{$unsigned((reg1256 ^ ((7'h58) ^ wire1062)))},
                  reg1250[(5'h12):(4'h8)]};
              reg1276 = ($unsigned((((reg1088 ? reg1137 : forvar1223) ?
                      $signed(reg1115) : (reg1265 ? (7'h46) : forvar1266)) ?
                  $signed(reg1247[(1'h0):(1'h0)]) : {(!reg1080),
                      $unsigned(reg1244)})) ^~ (reg1124[(5'h11):(4'hf)] && (((reg1262 ?
                          reg1112 : wire1063) ?
                      (reg1198 ? wire1215 : reg1229) : reg1237) ?
                  reg1131 : ((reg1096 != reg1186) ?
                      (reg1187 ? (7'h4c) : reg1183) : {reg1091,
                          reg1230,
                          reg1080}))));
              reg1277 = (8'ha0);
            end
          else
            begin
              reg1275 = (~((reg1091 ?
                  (^~$unsigned((8'hb2))) : $unsigned({reg1254,
                      reg1239,
                      reg1248})) >= (&reg1101[(2'h3):(1'h1)])));
              reg1276 = ((8'h9f) << $unsigned(reg1238));
              reg1277 = ($unsigned(((|(~(8'hb9))) || reg1235)) ?
                  $signed((~|$unsigned(reg1240))) : reg1131[(3'h4):(3'h4)]);
              reg1278 <= $signed(((7'h48) != {({reg1236, (8'haa), reg1229} ?
                      $signed(reg1163) : (~forvar1266))}));
              reg1279 = reg1233;
            end
          reg1280 = $unsigned(reg1267[(3'h5):(1'h0)]);
        end
      for (forvar1281 = (1'h0); (forvar1281 < (2'h3)); forvar1281 = (forvar1281 + (1'h1)))
        begin
          reg1282 <= {$unsigned((|reg1135[(4'hb):(3'h4)]))};
          reg1283 = ($unsigned((reg1068[(2'h2):(1'h1)] ^~ $signed($unsigned(reg1257)))) ?
              (8'ha9) : (reg1226 ~^ $unsigned((~&(reg1210 ?
                  reg1142 : reg1067)))));
        end
      for (forvar1284 = (1'h0); (forvar1284 < (3'h6)); forvar1284 = (forvar1284 + (1'h1)))
        begin
          reg1285 <= ((({reg1245, $signed((7'h43)), reg1153[(4'hc):(1'h0)]} ?
                      ($signed(reg1101) ?
                          (reg1263 ~^ reg1130) : reg1155[(4'hc):(2'h3)]) : {(reg1221 + (8'haa)),
                          {reg1209}}) ?
                  wire1065[(4'h8):(3'h6)] : ((reg1144 ?
                      reg1278 : reg1082[(1'h0):(1'h0)]) >>> ($signed((8'ha5)) ^ reg1231[(2'h3):(1'h0)]))) ?
              $signed({(reg1280[(3'h5):(1'h0)] ?
                      $unsigned(reg1278) : $unsigned(reg1202)),
                  (-reg1246[(5'h16):(2'h3)]),
                  (^~(reg1080 < reg1137))}) : reg1220[(2'h2):(1'h1)]);
          reg1286 = $signed($signed(reg1261));
        end
      for (forvar1287 = (1'h0); (forvar1287 < (3'h6)); forvar1287 = (forvar1287 + (1'h1)))
        begin
          for (forvar1288 = (1'h0); (forvar1288 < (3'h4)); forvar1288 = (forvar1288 + (1'h1)))
            begin
              reg1289 <= $unsigned(reg1251[(4'h8):(1'h1)]);
              reg1290 = ((forvar1223 - (^~($signed(reg1247) ^ (reg1254 ?
                  (8'ha4) : reg1256)))) >>> (~&(reg1251[(4'h9):(3'h5)] ?
                  $unsigned($signed(reg1236)) : $signed(forvar1281[(3'h4):(1'h0)]))));
              reg1291 <= (&reg1277);
              reg1292 = ((reg1233[(5'h1f):(3'h5)] ?
                      reg1155 : (~reg1232[(4'hf):(4'ha)])) ?
                  (reg1200[(4'hb):(1'h1)] ?
                      reg1192[(2'h3):(2'h2)] : $signed($unsigned(((7'h46) ?
                          wire1094 : reg1158)))) : (reg1087 ?
                      (8'hb6) : $unsigned(((~&forvar1219) ?
                          $signed(reg1091) : (reg1269 ? wire1216 : reg1254)))));
              reg1293 <= ((&(8'hb8)) ? reg1278[(4'h8):(4'h8)] : wire1060);
            end
          reg1294 <= wire1217;
          reg1295 = ((~&((7'h58) ?
              (7'h45) : $unsigned((^~reg1292)))) >= ((reg1084[(2'h3):(1'h1)] << (7'h45)) ?
              ($signed((7'h50)) ?
                  $unsigned((7'h57)) : (~&$unsigned((8'h9d)))) : ($unsigned($unsigned(reg1268)) ?
                  reg1174[(4'hd):(2'h2)] : $signed((reg1237 ^~ reg1191)))));
          if (reg1163)
            begin
              reg1296 = $unsigned($unsigned(reg1155));
              reg1297 = ($unsigned($unsigned(((reg1259 << reg1230) ?
                      {reg1198, reg1246, reg1268} : forvar1266))) ?
                  (($signed($signed((7'h54))) == (~^$unsigned(reg1144))) >= {((~^reg1271) ?
                          ((8'h9e) + reg1244) : (^~forvar1223))}) : (7'h40));
              reg1298 <= $unsigned($unsigned({reg1243[(1'h1):(1'h1)]}));
              reg1299 = reg1271;
              reg1300 <= (($unsigned(reg1142[(5'h14):(4'hd)]) >>> {forvar1258[(4'h8):(3'h7)]}) ?
                  $signed(($unsigned(reg1285[(4'h8):(1'h1)]) == reg1262)) : forvar1281[(2'h2):(1'h0)]);
              reg1301 <= (reg1250 ?
                  ($signed(reg1126[(3'h7):(3'h5)]) ?
                      (((!reg1163) ~^ {reg1169,
                          reg1115,
                          reg1084}) >> (~$signed(reg1176))) : (((&reg1249) <<< {reg1072,
                          reg1142,
                          reg1153}) >> ((reg1209 >= reg1119) ?
                          $signed(reg1137) : $unsigned(reg1240)))) : {{($unsigned(reg1282) != (&reg1191)),
                          (!(reg1103 ? reg1178 : reg1085)),
                          (!(~|reg1296))},
                      reg1245});
            end
          else
            begin
              reg1296 = (-(&$unsigned(($unsigned(forvar1258) + reg1286))));
              reg1298 <= {$unsigned({reg1130, $unsigned($unsigned(reg1235))})};
              reg1299 = {{(8'hba),
                      ({$unsigned(reg1277),
                          (-reg1249),
                          $unsigned(reg1280)} ~^ reg1178[(3'h5):(1'h0)]),
                      reg1243[(4'h8):(1'h1)]},
                  reg1103[(4'hc):(2'h2)]};
              reg1302 = (((reg1274[(2'h2):(1'h0)] * (~reg1093[(4'hf):(4'hb)])) ^ $unsigned((~|(reg1174 ?
                      (7'h41) : wire1062)))) ?
                  (~&(($signed(reg1245) ?
                      (^reg1254) : reg1252[(4'hb):(3'h7)]) | $signed(reg1279))) : reg1253[(3'h4):(2'h2)]);
              reg1303 = $signed(wire1215[(4'hc):(4'hb)]);
              reg1304 <= $unsigned($signed((reg1269 ?
                  ((reg1178 * reg1120) - reg1091[(5'h16):(4'he)]) : $unsigned((+(7'h56))))));
              reg1305 = reg1239;
            end
          for (forvar1306 = (1'h0); (forvar1306 < (1'h1)); forvar1306 = (forvar1306 + (1'h1)))
            begin
              reg1307 <= $unsigned($signed(reg1102[(3'h4):(1'h0)]));
              reg1308 <= $signed(reg1187[(3'h4):(2'h2)]);
              reg1309 = reg1210;
              reg1310 = $signed($unsigned(reg1282[(4'ha):(2'h3)]));
              reg1311 = ($signed((8'h9f)) <<< $unsigned((-$signed({reg1213}))));
              reg1312 = ($unsigned($unsigned($signed(reg1267))) == (~^$unsigned((~^(reg1297 ?
                  (8'ha0) : forvar1306)))));
              reg1313 <= reg1103;
            end
          reg1314 <= $unsigned(((-$unsigned((8'hb6))) ?
              ((7'h43) ^~ (((8'ha9) ? reg1233 : reg1277) ?
                  $signed(reg1085) : reg1151[(2'h3):(2'h3)])) : reg1233));
          if (reg1108)
            begin
              reg1315 <= reg1163[(1'h0):(1'h0)];
              reg1316 = (reg1202[(3'h5):(2'h3)] && (~({$signed((7'h53))} ?
                  reg1292 : (8'hbb))));
              reg1317 <= reg1135[(5'h12):(4'hf)];
              reg1318 <= reg1183;
              reg1319 <= $unsigned(((~|(^$signed(wire1062))) & $unsigned(reg1233)));
            end
          else
            begin
              reg1315 <= reg1213;
              reg1316 = ((reg1279[(4'he):(3'h6)] <= reg1120) ?
                  $unsigned((~|(^(reg1186 ? reg1236 : (7'h40))))) : (7'h53));
              reg1317 <= {$signed(wire1216[(4'hc):(4'hb)]),
                  $unsigned($unsigned((7'h4b)))};
              reg1320 = ($unsigned({({reg1143, (7'h49)} ?
                          $unsigned((8'ha3)) : reg1112),
                      {reg1096},
                      $signed(((8'ha1) ? reg1299 : (7'h48)))}) ?
                  (-(($unsigned(reg1199) & (~reg1253)) >>> (7'h56))) : (7'h46));
              reg1321 = reg1191;
              reg1322 = reg1200[(3'h6):(2'h2)];
              reg1323 <= $unsigned(($unsigned(reg1322) || ($unsigned((8'hae)) >> reg1294[(2'h2):(1'h1)])));
            end
        end
    end
endmodule