(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h43c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire0;
  input wire [(5'h17):(1'h0)] wire1;
  input wire signed [(5'h16):(1'h0)] wire2;
  input wire signed [(4'he):(1'h0)] wire3;
  input wire signed [(5'h16):(1'h0)] wire4;
  wire signed [(5'h11):(1'h0)] wire765;
  wire [(4'h8):(1'h0)] wire764;
  wire [(4'ha):(1'h0)] wire763;
  wire [(3'h4):(1'h0)] wire762;
  wire signed [(3'h5):(1'h0)] wire761;
  wire [(4'h8):(1'h0)] wire760;
  wire [(3'h4):(1'h0)] wire759;
  wire signed [(3'h7):(1'h0)] wire749;
  reg [(5'h16):(1'h0)] reg5 = (1'h0);
  reg [(4'h8):(1'h0)] reg6 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7 = (1'h0);
  reg [(4'ha):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar11 = (1'h0);
  reg [(5'h13):(1'h0)] reg12 = (1'h0);
  reg [(5'h16):(1'h0)] reg13 = (1'h0);
  reg [(5'h15):(1'h0)] reg14 = (1'h0);
  reg signed [(4'he):(1'h0)] reg15 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg16 = (1'h0);
  reg [(5'h13):(1'h0)] reg17 = (1'h0);
  reg [(5'h16):(1'h0)] reg18 = (1'h0);
  reg [(5'h16):(1'h0)] reg19 = (1'h0);
  reg [(5'h11):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg21 = (1'h0);
  reg [(4'hb):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg23 = (1'h0);
  reg [(5'h10):(1'h0)] reg24 = (1'h0);
  reg [(5'h14):(1'h0)] forvar25 = (1'h0);
  reg [(5'h13):(1'h0)] reg26 = (1'h0);
  reg [(3'h6):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg28 = (1'h0);
  reg [(5'h13):(1'h0)] reg29 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg30 = (1'h0);
  reg [(5'h11):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg32 = (1'h0);
  reg [(4'hf):(1'h0)] reg33 = (1'h0);
  reg [(5'h14):(1'h0)] reg34 = (1'h0);
  reg [(4'hc):(1'h0)] reg35 = (1'h0);
  reg [(5'h14):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg37 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg38 = (1'h0);
  reg [(2'h3):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg40 = (1'h0);
  reg [(3'h7):(1'h0)] forvar41 = (1'h0);
  reg signed [(4'he):(1'h0)] reg42 = (1'h0);
  reg [(4'hd):(1'h0)] reg43 = (1'h0);
  reg [(4'ha):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg45 = (1'h0);
  reg [(4'ha):(1'h0)] reg46 = (1'h0);
  reg [(5'h10):(1'h0)] reg47 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg48 = (1'h0);
  reg [(5'h14):(1'h0)] reg49 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg50 = (1'h0);
  reg [(3'h4):(1'h0)] reg51 = (1'h0);
  reg [(5'h10):(1'h0)] reg52 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar53 = (1'h0);
  reg [(4'ha):(1'h0)] reg54 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg55 = (1'h0);
  reg [(5'h11):(1'h0)] reg56 = (1'h0);
  reg [(5'h16):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar58 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg59 = (1'h0);
  reg [(5'h15):(1'h0)] reg60 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire61;
  wire [(5'h16):(1'h0)] wire62;
  wire [(3'h4):(1'h0)] wire747;
  reg [(4'hf):(1'h0)] forvar751 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar752 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg753 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg754 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar755 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg756 = (1'h0);
  wire [(5'h13):(1'h0)] wire757;
  assign y = {wire765,
                 wire764,
                 wire763,
                 wire762,
                 wire761,
                 wire760,
                 wire759,
                 wire749,
                 reg5,
                 reg6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 forvar11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 forvar25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 reg34,
                 reg35,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 forvar41,
                 reg42,
                 reg43,
                 reg41,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 reg52,
                 forvar53,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 forvar58,
                 reg59,
                 reg60,
                 wire61,
                 wire62,
                 wire747,
                 forvar751,
                 forvar752,
                 reg753,
                 reg754,
                 forvar755,
                 reg756,
                 wire757,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg5 <= wire1[(2'h3):(1'h0)];
      if ($signed((8'hbf)))
        begin
          if ("NeWoApT26DBhlr9dG")
            begin
              reg6 <= (wire4 << wire0[(4'he):(4'hb)]);
            end
          else
            begin
              reg6 = wire4[(4'h9):(3'h5)];
              reg7 <= (^($unsigned(reg5[(1'h0):(1'h0)]) ^ ($unsigned((+wire3)) > ((wire1 ?
                      wire1 : wire4) ?
                  $signed(wire2) : {wire1, reg5}))));
              reg8 <= reg7[(3'h7):(2'h3)];
              reg9 <= $unsigned("wzpa37o4VcwHadxDfJ4");
              reg10 <= "qNFOMe20FkRnvcSAnL";
            end
          for (forvar11 = (1'h0); (forvar11 < (1'h1)); forvar11 = (forvar11 + (1'h1)))
            begin
              reg12 <= (+$unsigned($signed(((reg10 && forvar11) ^ reg10[(4'h8):(1'h0)]))));
              reg13 = $signed(((($unsigned(reg5) - (reg6 <= wire1)) ?
                      (|$signed(reg12)) : reg9) ?
                  reg9[(1'h0):(1'h0)] : (-$signed(((8'ha1) != (7'h42))))));
              reg14 <= ((reg8 ?
                  "1xQz9JZuARWEVMPl" : (|$signed((reg12 ?
                      wire3 : (8'hb3))))) << $signed(reg10[(3'h6):(1'h0)]));
              reg15 = ($signed("YvOQfXtbHKI") ?
                  $signed(reg5[(5'h11):(3'h5)]) : {($signed($unsigned(wire1)) * reg10),
                      ({"vDABJm", $signed(reg10)} ? (8'hb1) : reg9)});
            end
          if ({$signed("EbmCpy2KUBa")})
            begin
              reg16 <= (-wire4[(2'h2):(1'h0)]);
              reg17 = $signed("L2gGcD0WSqEzhqRfz4pT");
              reg18 <= wire3;
              reg19 <= $signed((~&wire0[(4'h8):(3'h4)]));
              reg20 <= (reg19 != ("1RdTZ0BWsdqZ" ? reg7 : (&wire0)));
            end
          else
            begin
              reg16 <= $unsigned((7'h47));
              reg17 <= "Mh0uFwMOM0ErB1PaHO";
              reg18 <= (((&reg9[(4'h8):(3'h6)]) >> reg10[(4'ha):(3'h4)]) ?
                  "briRCi30afpFSNQ" : reg18[(2'h2):(1'h1)]);
              reg19 <= (~&reg14[(4'h9):(1'h1)]);
            end
        end
      else
        begin
          reg6 <= "xTFOmfa0DFDPZCUSg";
        end
      if ((8'ha9))
        begin
          if ($signed(reg5))
            begin
              reg21 <= (((~&(wire3[(3'h5):(1'h1)] ? reg14 : $signed(reg9))) ?
                      (8'hb8) : ({((8'hb6) >> reg12),
                          (reg17 || reg5)} >> $unsigned((reg10 >>> forvar11)))) ?
                  reg7[(4'h9):(2'h3)] : ((|{wire0}) & (reg19[(4'h8):(4'h8)] ^~ $signed($unsigned(reg20)))));
            end
          else
            begin
              reg21 <= $signed((($signed((reg21 ? reg9 : wire4)) ?
                  reg14[(4'he):(4'hb)] : $signed(reg5)) << ($signed("HluKg090P9VfDOuHchG") <= "3urxp3rX1v6qq6Bme")));
              reg22 <= (("I219qMfPZ7mH6XvGVml3Ng" && reg15) ?
                  ($unsigned(((wire3 <= wire2) == (forvar11 ?
                          reg21 : (7'h47)))) ?
                      $signed("zKCEM0NSdoczw") : ("sAyhqd0xQ6TEv" ^~ $unsigned("hwTfxaubnNG2TZGUpOJD"))) : reg12);
              reg23 <= (-(reg8 ?
                  reg17[(3'h7):(2'h2)] : $unsigned("RuZxzbo2fD0BBQ")));
            end
        end
      else
        begin
          if (reg16[(1'h1):(1'h1)])
            begin
              reg21 <= {(8'hba)};
              reg22 <= $unsigned(($signed(($signed(reg19) <<< "chU37MoRzSgNddqMnW")) < $signed($unsigned(reg19))));
            end
          else
            begin
              reg21 <= $signed(((("" ? $unsigned(reg21) : wire0) ?
                      (forvar11 ? {reg18} : {(7'h47)}) : {(-(8'ha0)),
                          $unsigned(wire4)}) ?
                  reg18[(3'h5):(2'h3)] : (8'hb0)));
              reg22 <= (|$unsigned(({reg13[(3'h7):(3'h5)]} == ({reg10, reg17} ?
                  $signed(reg8) : (~|reg13)))));
              reg23 = "GxNX3g";
            end
          if ($signed(wire3))
            begin
              reg24 <= ({"ArTtvSEP"} | ((reg16[(1'h0):(1'h0)] ?
                  ((reg15 <<< reg14) <= (reg20 - reg18)) : ($unsigned((8'hb9)) == (reg15 != reg14))) > ((|"uUfutFgtyt3olUA492") ?
                  $unsigned(wire4[(2'h3):(1'h0)]) : $unsigned($signed((8'hab))))));
            end
          else
            begin
              reg24 <= (8'ha5);
            end
          for (forvar25 = (1'h0); (forvar25 < (2'h2)); forvar25 = (forvar25 + (1'h1)))
            begin
              reg26 <= "4PxYXBsLYKQck4M9";
              reg27 <= reg23;
              reg28 <= wire4[(4'h9):(1'h1)];
              reg29 <= $unsigned($signed("Cz"));
              reg30 <= forvar25[(1'h0):(1'h0)];
            end
          if (reg19[(2'h3):(2'h3)])
            begin
              reg31 = {reg8[(3'h7):(3'h4)], $signed((8'hae))};
              reg32 <= $signed(reg7);
              reg33 <= "SatqnOC";
              reg34 <= {($unsigned((reg6 ?
                      $signed((8'hb1)) : (reg32 ?
                          wire2 : reg27))) < reg29[(4'hd):(1'h0)])};
            end
          else
            begin
              reg31 = "k0";
              reg32 <= ("eGxSO" || (8'hac));
              reg33 = (forvar25[(5'h11):(3'h7)] ?
                  ("t5yIF8t1bghcYApBa" * "MT1nSeYl9l3") : ("t" ?
                      (^(-"NRU7rCGbAwdMoif")) : ($unsigned($signed(wire2)) ~^ (reg10 || (reg15 ?
                          reg12 : reg28)))));
              reg34 <= "";
              reg35 <= reg20[(4'hc):(2'h3)];
            end
          if (reg13)
            begin
              reg36 <= (&$unsigned((~&(~reg35))));
              reg37 <= reg9;
              reg38 <= $signed(reg19);
              reg39 <= reg17[(3'h7):(3'h5)];
              reg40 <= {(forvar11[(1'h1):(1'h1)] ?
                      "0nQUAGPskcTFIAVQfDi" : ($unsigned(reg10) ?
                          $unsigned(((7'h43) ?
                              reg22 : wire3)) : reg37[(2'h2):(1'h1)]))};
            end
          else
            begin
              reg36 <= $unsigned((($signed(reg27) ?
                  "yM4dowpwylARMQu0QUJk" : reg26) * reg33[(4'h9):(3'h4)]));
              reg37 <= ("Ay5mtOs30KIPuW" - $signed($unsigned("EppPVZEvB")));
              reg38 <= ("UMNM6H" ? reg13 : "M8rxAXE6QcLZPRhAUUXf");
            end
        end
      if ($unsigned($signed((((reg14 ? reg40 : wire2) ?
              ((7'h48) == reg31) : $unsigned((7'h42))) ?
          ((reg18 && reg8) - (reg9 ?
              (8'h9e) : reg20)) : (((8'hb6) + (7'h45)) | (forvar11 & reg8))))))
        begin
          for (forvar41 = (1'h0); (forvar41 < (1'h0)); forvar41 = (forvar41 + (1'h1)))
            begin
              reg42 <= ({reg23} ?
                  $unsigned(({$signed((8'haf)), $unsigned(reg27)} ?
                      "kCzqVbp17" : (reg13[(1'h0):(1'h0)] ^~ (wire0 ?
                          reg9 : reg7)))) : (reg9 ?
                      ({(reg29 ^~ reg38)} ?
                          reg33 : (~|(~^forvar11))) : (({(8'ha2)} > (^reg36)) ^ $unsigned({reg9}))));
              reg43 <= "W4C5Uil2u";
            end
        end
      else
        begin
          if ((~$unsigned("CDh3xMa5T")))
            begin
              reg41 <= $unsigned(($signed(reg15) ?
                  $signed(($unsigned((8'hb2)) ?
                      $unsigned(reg20) : {reg43,
                          reg27})) : ($unsigned(reg9[(3'h6):(3'h5)]) && $signed(reg29))));
              reg42 = $signed($signed($unsigned(((reg29 && reg39) ?
                  "J" : reg27[(2'h3):(1'h0)]))));
              reg43 <= (|reg19[(5'h12):(3'h7)]);
            end
          else
            begin
              reg41 <= (~((^reg13) ?
                  ("qggMvSFTugU8YJb" - $signed($unsigned(reg19))) : (8'ha5)));
              reg42 <= $unsigned($unsigned($unsigned((forvar25[(4'ha):(1'h0)] ^ {wire0}))));
              reg43 <= reg26[(4'h8):(3'h5)];
              reg44 <= reg27[(1'h0):(1'h0)];
            end
          reg45 <= (+$signed((reg17 ?
              ((reg13 ^~ reg6) ? (reg42 ? (8'ha2) : reg7) : reg24) : reg27)));
          reg46 <= "NohUYfWDf7fo0IvGNVLT";
          if (reg15[(1'h1):(1'h0)])
            begin
              reg47 <= "IxFQBdSU6lwSvu";
              reg48 <= $unsigned($unsigned((8'hae)));
              reg49 <= "";
              reg50 <= reg45;
              reg51 <= ({reg44[(4'hd):(2'h2)],
                  {"haOgHlFOEshaTscqOY"}} << $unsigned($unsigned("Z")));
            end
          else
            begin
              reg47 = (~reg12[(4'ha):(1'h0)]);
            end
          reg52 <= reg23;
        end
      if ($signed((reg21[(4'hd):(3'h5)] * (((reg15 >>> reg29) ?
              $signed(reg15) : (wire0 ? reg44 : reg43)) ?
          ((&reg23) && $unsigned(reg6)) : $unsigned($signed(reg45))))))
        begin
          for (forvar53 = (1'h0); (forvar53 < (1'h0)); forvar53 = (forvar53 + (1'h1)))
            begin
              reg54 <= wire0;
            end
        end
      else
        begin
          for (forvar53 = (1'h0); (forvar53 < (1'h0)); forvar53 = (forvar53 + (1'h1)))
            begin
              reg54 <= "70LuflJiO4y3d";
              reg55 <= "7sd0o4ymcgkhbcuRAeG";
              reg56 <= reg6[(3'h5):(2'h2)];
              reg57 <= (^~$signed($unsigned("UOiX15D021156Ftp8m")));
            end
          for (forvar58 = (1'h0); (forvar58 < (3'h4)); forvar58 = (forvar58 + (1'h1)))
            begin
              reg59 <= ((reg13[(4'hf):(3'h4)] ?
                  ((|(reg34 || reg14)) ?
                      (reg28[(4'hf):(2'h2)] ?
                          "apn9WnAiADOa5CDkTMBb" : $signed((8'ha3))) : {$signed(reg32),
                          $signed(reg22)}) : reg40[(1'h0):(1'h0)]) & reg50);
              reg60 <= reg18;
            end
        end
    end
  assign wire61 = reg18;
  assign wire62 = ((8'h9c) ? "gU" : $unsigned(reg28));
  module63 modinst748 (.wire64(wire4), .wire67(reg15), .wire68(reg29), .y(wire747), .clk(clk), .wire66(reg40), .wire65(reg49));
  module63 modinst750 (wire749, clk, reg17, reg49, forvar25, reg36, wire2);
  always
    @(posedge clk) begin
      for (forvar751 = (1'h0); (forvar751 < (1'h1)); forvar751 = (forvar751 + (1'h1)))
        begin
          for (forvar752 = (1'h0); (forvar752 < (2'h3)); forvar752 = (forvar752 + (1'h1)))
            begin
              reg753 = reg20[(2'h2):(1'h1)];
            end
          reg754 = {$signed(reg26)};
          for (forvar755 = (1'h0); (forvar755 < (2'h3)); forvar755 = (forvar755 + (1'h1)))
            begin
              reg756 <= (forvar11[(3'h5):(3'h5)] ?
                  (reg7 ?
                      (("7sFn4mZY0evHSA91nkdCF" ?
                              $unsigned((8'hb5)) : (reg35 >= wire62)) ?
                          $signed("R6Wwmys1JmQKeN42K0tds") : {(reg13 ^ (8'hbc)),
                              (reg42 ?
                                  forvar58 : reg5)}) : (forvar755 * $signed({reg55}))) : ($signed($signed(reg56)) ?
                      (~|reg26) : (8'hb8)));
            end
        end
    end
  module374 modinst758 (.wire378(reg21), .clk(clk), .wire379(reg36), .wire376(reg753), .wire375(reg20), .wire377(reg35), .y(wire757));
  assign wire759 = reg23[(4'hb):(4'h9)];
  assign wire760 = (8'hb1);
  assign wire761 = wire61[(5'h13):(3'h7)];
  assign wire762 = forvar751[(4'hb):(4'h9)];
  assign wire763 = "GT0Ad5rV9lAxCnnRZF0qr";
  assign wire764 = {$signed((|{(wire62 ? reg40 : (8'ha2))}))};
  assign wire765 = $signed($signed($signed(wire760)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module63
#( parameter param746 = (~&((~|({(8'ha6)} << ((7'h41) ? (8'hbc) : (7'h48)))) <<< ((+(|(8'ha0))) >> {((7'h42) && (7'h45))}))) )
(y, clk, wire68, wire67, wire66, wire65, wire64);
  output wire [(32'h35a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire68;
  input wire [(4'he):(1'h0)] wire67;
  input wire [(5'h10):(1'h0)] wire66;
  input wire [(5'h14):(1'h0)] wire65;
  input wire signed [(5'h16):(1'h0)] wire64;
  reg signed [(4'h8):(1'h0)] reg737 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg745 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg744 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg743 = (1'h0);
  reg [(4'h9):(1'h0)] forvar742 = (1'h0);
  reg [(4'he):(1'h0)] reg741 = (1'h0);
  reg [(4'ha):(1'h0)] reg740 = (1'h0);
  reg [(4'h9):(1'h0)] reg739 = (1'h0);
  reg [(4'hf):(1'h0)] reg738 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar737 = (1'h0);
  reg [(5'h15):(1'h0)] reg736 = (1'h0);
  reg [(5'h12):(1'h0)] reg735 = (1'h0);
  reg [(5'h15):(1'h0)] reg734 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg733 = (1'h0);
  reg [(2'h3):(1'h0)] reg732 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar731 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg730 = (1'h0);
  reg [(5'h14):(1'h0)] forvar729 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg728 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg727 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg726 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg725 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg724 = (1'h0);
  reg [(4'h8):(1'h0)] reg723 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg722 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar721 = (1'h0);
  reg [(3'h4):(1'h0)] reg720 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg719 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire718;
  wire signed [(3'h5):(1'h0)] wire717;
  wire [(5'h13):(1'h0)] wire715;
  wire signed [(5'h17):(1'h0)] wire674;
  wire [(4'hd):(1'h0)] wire676;
  wire [(4'hb):(1'h0)] wire677;
  reg [(5'h13):(1'h0)] forvar678 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg679 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg680 = (1'h0);
  reg [(5'h13):(1'h0)] reg681 = (1'h0);
  reg [(4'h9):(1'h0)] reg682 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg683 = (1'h0);
  reg [(4'hb):(1'h0)] reg684 = (1'h0);
  reg [(5'h13):(1'h0)] reg685 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg687 = (1'h0);
  reg [(4'hc):(1'h0)] reg688 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar689 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar690 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg691 = (1'h0);
  reg [(3'h7):(1'h0)] reg692 = (1'h0);
  reg [(4'he):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg694 = (1'h0);
  reg [(3'h6):(1'h0)] reg695 = (1'h0);
  reg [(2'h3):(1'h0)] forvar696 = (1'h0);
  reg [(5'h13):(1'h0)] reg697 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg698 = (1'h0);
  reg [(5'h16):(1'h0)] reg699 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg700 = (1'h0);
  reg signed [(4'he):(1'h0)] reg701 = (1'h0);
  reg [(2'h3):(1'h0)] forvar702 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg703 = (1'h0);
  reg [(5'h16):(1'h0)] reg704 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg705 = (1'h0);
  reg [(4'hb):(1'h0)] reg706 = (1'h0);
  wire [(5'h16):(1'h0)] wire707;
  wire signed [(4'hb):(1'h0)] wire708;
  wire [(5'h11):(1'h0)] wire709;
  wire [(5'h16):(1'h0)] wire710;
  wire [(4'hb):(1'h0)] wire711;
  wire [(4'hf):(1'h0)] wire713;
  assign y = {reg737,
                 reg745,
                 reg744,
                 reg743,
                 forvar742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 forvar737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 forvar731,
                 reg730,
                 forvar729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 reg723,
                 reg722,
                 forvar721,
                 reg720,
                 reg719,
                 wire718,
                 wire717,
                 wire715,
                 wire674,
                 wire676,
                 wire677,
                 forvar678,
                 reg679,
                 reg680,
                 reg681,
                 reg682,
                 reg683,
                 reg684,
                 reg685,
                 reg686,
                 reg687,
                 reg688,
                 forvar689,
                 forvar690,
                 reg691,
                 reg692,
                 reg693,
                 reg694,
                 reg695,
                 forvar696,
                 reg697,
                 reg698,
                 reg699,
                 reg700,
                 reg701,
                 forvar702,
                 reg703,
                 reg704,
                 reg705,
                 reg706,
                 wire707,
                 wire708,
                 wire709,
                 wire710,
                 wire711,
                 wire713,
                 (1'h0)};
  module69 modinst675 (wire674, clk, wire64, wire65, wire68, wire67, wire66);
  assign wire676 = $unsigned("53X0JbfCs");
  assign wire677 = "ktYFoWx6f4TyN08Xv";
  always
    @(posedge clk) begin
      for (forvar678 = (1'h0); (forvar678 < (1'h1)); forvar678 = (forvar678 + (1'h1)))
        begin
          if (wire67[(4'he):(1'h1)])
            begin
              reg679 = $unsigned(("Qt9xw1cQ20HK2wte" ^~ $unsigned((7'h46))));
              reg680 = wire66;
            end
          else
            begin
              reg679 <= {"JR1g4D1KvX5xQTyDzk", wire66};
              reg680 <= reg679[(4'hb):(4'h8)];
              reg681 <= {{""}, $signed((wire674 > reg679))};
              reg682 = forvar678[(2'h3):(2'h3)];
            end
          reg683 <= ((~&reg679[(3'h7):(3'h5)]) ?
              {($unsigned((~|reg679)) == $unsigned(wire65[(5'h13):(2'h2)])),
                  $unsigned("rhgZguKtuRNMtv60JWQ91")} : reg682[(3'h6):(2'h2)]);
          if ((wire677[(3'h7):(1'h1)] | $signed((forvar678[(5'h10):(4'hf)] ~^ {((7'h47) > reg681),
              $unsigned(wire66)}))))
            begin
              reg684 <= {("iPmyLcStYEGmT5mu7r0s" ?
                      (&$signed("Ua4ug9v8VrcZT")) : (-wire67[(1'h0):(1'h0)]))};
              reg685 <= reg682;
              reg686 <= ($unsigned($unsigned(((-reg679) >>> (~^wire676)))) || ({(~^{wire64,
                          (8'hb7)})} ?
                  (wire67[(1'h1):(1'h0)] <= {wire674[(5'h12):(4'hc)]}) : wire65[(1'h0):(1'h0)]));
              reg687 <= ($signed({{$signed(reg680)}}) ?
                  $signed($signed(reg685[(3'h4):(2'h3)])) : "tprnQCSRIPWTbJda");
              reg688 <= ($signed(wire68[(4'he):(2'h3)]) ?
                  {(^($signed(reg679) >= (reg684 < wire677))),
                      reg681[(2'h2):(1'h0)]} : reg687);
            end
          else
            begin
              reg684 <= ($unsigned(("TKZkpiAENOz" ?
                      ((reg682 && forvar678) & wire68[(4'hf):(4'h9)]) : ((reg679 ?
                          reg683 : reg680) >> reg681[(4'h8):(2'h3)]))) ?
                  $unsigned($signed({wire64})) : reg685);
            end
        end
      for (forvar689 = (1'h0); (forvar689 < (3'h4)); forvar689 = (forvar689 + (1'h1)))
        begin
          for (forvar690 = (1'h0); (forvar690 < (2'h3)); forvar690 = (forvar690 + (1'h1)))
            begin
              reg691 <= (8'ha3);
              reg692 <= "nozNyFK6DBVifEz";
              reg693 = ((reg687[(5'h15):(5'h13)] <= "ikgAmLER") >= $signed(reg680));
              reg694 = $unsigned($signed(reg685));
              reg695 <= $signed($signed({wire66[(1'h1):(1'h0)]}));
            end
          for (forvar696 = (1'h0); (forvar696 < (1'h1)); forvar696 = (forvar696 + (1'h1)))
            begin
              reg697 <= forvar678[(5'h11):(2'h2)];
              reg698 <= wire66;
              reg699 <= $signed("9rhoZ7yyRrKPCwRypYD");
              reg700 <= "o4gwYQ4OoAc1ipXJ4";
              reg701 <= $signed(wire64);
            end
          for (forvar702 = (1'h0); (forvar702 < (2'h3)); forvar702 = (forvar702 + (1'h1)))
            begin
              reg703 <= (&$unsigned(($signed(reg692[(3'h4):(1'h1)]) ?
                  $signed("RCBmXLqC9fa95ebMR2urpZ") : reg700[(1'h0):(1'h0)])));
              reg704 <= (~^$signed($unsigned(((reg697 ?
                  reg703 : (8'hb8)) <<< $unsigned((8'hbf))))));
              reg705 <= reg687[(4'he):(4'ha)];
              reg706 <= ((8'hbc) && ($signed({$signed(reg686)}) ?
                  $unsigned(((reg681 | forvar696) ?
                      $signed(wire677) : wire65)) : (^reg687)));
            end
        end
    end
  assign wire707 = (($signed((~(reg700 ~^ forvar689))) ?
                       $unsigned(({(7'h43), reg695} ?
                           (reg698 ?
                               reg706 : reg679) : (8'hb0))) : $signed($signed("idgogdKiaC7f7KsvtvDa4"))) >> ((&$unsigned((reg692 ?
                       (8'ha2) : reg681))) & (wire67 + ((reg695 - reg705) & (forvar678 - (7'h41))))));
  assign wire708 = (((~|"LuWOWTrwV") ?
                       ("u5RAYJAy4xbFMvbo9R" ?
                           forvar702 : (reg705 ?
                               (!reg701) : (forvar690 ?
                                   reg704 : (8'ha1)))) : wire707[(2'h3):(1'h0)]) * ((reg679[(2'h3):(1'h0)] <= forvar696) ?
                       "gsEyN5GWXCMzmw" : {$signed(forvar696[(2'h3):(2'h3)]),
                           reg694}));
  assign wire709 = $signed({(8'hb7)});
  assign wire710 = $signed(((((wire707 ? wire67 : reg698) ?
                       reg705[(5'h10):(4'hd)] : {wire67}) && reg699[(3'h6):(2'h2)]) >>> $unsigned($unsigned($signed((8'hbb))))));
  module326 modinst712 (wire711, clk, wire68, reg682, reg699, reg681);
  module609 modinst714 (.wire611(reg684), .wire613(reg679), .wire614(reg688), .y(wire713), .wire612(wire676), .clk(clk), .wire610(reg685));
  module95 modinst716 (.wire98(reg699), .y(wire715), .wire99(wire710), .clk(clk), .wire96(reg706), .wire97(reg698));
  assign wire717 = (&{(8'hb3), $signed(wire67)});
  assign wire718 = {$signed(forvar696)};
  always
    @(posedge clk) begin
      reg719 <= forvar678;
      reg720 <= $unsigned(wire707[(4'hb):(3'h6)]);
      for (forvar721 = (1'h0); (forvar721 < (2'h3)); forvar721 = (forvar721 + (1'h1)))
        begin
          if (reg684)
            begin
              reg722 <= (8'hb2);
              reg723 <= (("teqQivWMCDEfI" ?
                      reg682 : (reg683 ?
                          ({wire708} <<< (forvar689 | wire676)) : reg684[(4'ha):(1'h0)])) ?
                  reg680 : "0JVllAGGAsMK3WMlDO");
              reg724 <= $unsigned((~&("lt7ubxk7XxrBIHD9GeaMz2" ?
                  (reg692[(1'h1):(1'h0)] ?
                      $signed(wire66) : $signed(reg720)) : {reg720[(2'h3):(2'h2)]})));
              reg725 <= forvar690;
              reg726 <= wire713[(1'h0):(1'h0)];
            end
          else
            begin
              reg722 <= ((("Jdz7" ?
                      (reg698 ^~ (forvar696 ?
                          reg699 : (8'hab))) : ((reg699 <<< (8'hac)) <= $unsigned((8'hb6)))) * reg722[(1'h1):(1'h1)]) ?
                  "mXpJ5HRZhcwUT7KVkgcS9A" : ((&("75szgI" ?
                          (reg680 && (8'hbf)) : {(8'h9f)})) ?
                      "qsbw8uHD1NoPCKM1qDBzx" : ($unsigned((reg724 ?
                          wire65 : wire68)) <<< ((wire707 ^ (8'hac)) <= (reg700 | forvar690)))));
            end
          if ({reg699[(2'h3):(2'h3)],
              (wire708[(1'h1):(1'h0)] + $signed((~&(reg681 ?
                  (7'h43) : reg724))))})
            begin
              reg727 <= ("dLv" >= ("pAGdt" || ""));
              reg728 <= $unsigned(($unsigned((~reg683)) ?
                  $signed(reg699[(4'hc):(4'h9)]) : $unsigned($signed($unsigned(reg687)))));
            end
          else
            begin
              reg727 = ($signed($signed(reg706)) | (-$unsigned($unsigned($unsigned(reg726)))));
            end
          for (forvar729 = (1'h0); (forvar729 < (2'h3)); forvar729 = (forvar729 + (1'h1)))
            begin
              reg730 <= (~|"YUaP32frrI3YN");
            end
          for (forvar731 = (1'h0); (forvar731 < (3'h4)); forvar731 = (forvar731 + (1'h1)))
            begin
              reg732 <= reg688[(3'h4):(1'h1)];
              reg733 <= (!$signed($signed(wire715)));
              reg734 <= (-$signed((reg686[(2'h3):(2'h2)] ?
                  wire713 : wire68[(1'h0):(1'h0)])));
              reg735 <= {"76kLdykOf2UA2E5",
                  $unsigned($signed((reg727[(2'h3):(1'h0)] ?
                      $signed(reg704) : "5")))};
            end
          reg736 <= {$unsigned(wire709[(3'h4):(2'h3)])};
        end
      if (reg726)
        begin
          for (forvar737 = (1'h0); (forvar737 < (3'h4)); forvar737 = (forvar737 + (1'h1)))
            begin
              reg738 <= (8'hbd);
              reg739 <= reg684;
              reg740 = "oe";
              reg741 <= reg704;
            end
          for (forvar742 = (1'h0); (forvar742 < (1'h0)); forvar742 = (forvar742 + (1'h1)))
            begin
              reg743 <= {(~^($unsigned((|reg693)) - {$signed(reg726)}))};
              reg744 <= forvar696[(1'h1):(1'h0)];
              reg745 <= wire710;
            end
        end
      else
        begin
          reg737 <= (~|($signed(reg695) | $unsigned(((!reg720) && $signed(forvar702)))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module69  (y, clk, wire70, wire71, wire72, wire73, wire74);
  output wire [(32'h1b1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h16):(1'h0)] wire70;
  input wire signed [(5'h14):(1'h0)] wire71;
  input wire signed [(5'h13):(1'h0)] wire72;
  input wire signed [(2'h2):(1'h0)] wire73;
  input wire [(4'hc):(1'h0)] wire74;
  wire [(4'he):(1'h0)] wire673;
  wire signed [(4'hf):(1'h0)] wire672;
  wire [(3'h7):(1'h0)] wire671;
  wire signed [(3'h6):(1'h0)] wire670;
  wire [(4'hb):(1'h0)] wire669;
  wire [(3'h5):(1'h0)] wire668;
  wire [(5'h12):(1'h0)] wire667;
  wire signed [(5'h16):(1'h0)] wire659;
  wire [(4'h9):(1'h0)] wire657;
  wire [(5'h13):(1'h0)] wire325;
  wire signed [(5'h11):(1'h0)] wire324;
  wire signed [(4'hf):(1'h0)] wire75;
  reg [(5'h16):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar77 = (1'h0);
  reg [(5'h15):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar79 = (1'h0);
  reg [(5'h10):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg81 = (1'h0);
  reg [(4'ha):(1'h0)] reg82 = (1'h0);
  reg [(4'hd):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar84 = (1'h0);
  reg [(5'h13):(1'h0)] reg85 = (1'h0);
  reg [(5'h12):(1'h0)] reg86 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg87 = (1'h0);
  wire [(5'h10):(1'h0)] wire322;
  wire [(4'he):(1'h0)] wire661;
  wire signed [(4'h9):(1'h0)] wire662;
  wire [(5'h16):(1'h0)] wire664;
  wire signed [(4'ha):(1'h0)] wire665;
  assign y = {wire673,
                 wire672,
                 wire671,
                 wire670,
                 wire669,
                 wire668,
                 wire667,
                 wire659,
                 wire657,
                 wire325,
                 wire324,
                 wire75,
                 reg76,
                 forvar77,
                 reg78,
                 forvar79,
                 reg80,
                 reg81,
                 reg82,
                 reg83,
                 forvar84,
                 reg85,
                 reg86,
                 reg87,
                 wire322,
                 wire661,
                 wire662,
                 wire664,
                 wire665,
                 (1'h0)};
  assign wire75 = $signed(wire73[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg76 <= "e4xBtHIZQYGDJ";
      for (forvar77 = (1'h0); (forvar77 < (1'h1)); forvar77 = (forvar77 + (1'h1)))
        begin
          reg78 <= $unsigned("5uR40pMTVhT5R");
        end
      for (forvar79 = (1'h0); (forvar79 < (1'h0)); forvar79 = (forvar79 + (1'h1)))
        begin
          if ((($signed("LTlPz") ?
              ("CVwrDUgqnDzGYvAvlrWv" ?
                  "2hnFm" : "Z84z7wBal6OFhiNExi") : $unsigned(reg78)) & ({$signed({wire71,
                      (8'ha6)}),
                  ({wire70} == reg76[(3'h4):(3'h4)])} ?
              $signed(wire71) : $signed(wire74))))
            begin
              reg80 <= wire73[(2'h2):(1'h0)];
              reg81 <= (7'h43);
              reg82 <= (~^$signed($signed((forvar77[(3'h6):(3'h6)] && (8'ha9)))));
              reg83 <= "bOlB3v0Lk09D3f";
            end
          else
            begin
              reg80 <= $unsigned({$unsigned(reg80[(1'h1):(1'h0)]),
                  ((wire70[(2'h2):(1'h0)] ?
                      {wire74, reg83} : reg76[(2'h3):(1'h1)]) || (|{forvar77,
                      wire75}))});
            end
          for (forvar84 = (1'h0); (forvar84 < (1'h1)); forvar84 = (forvar84 + (1'h1)))
            begin
              reg85 <= reg83[(3'h4):(2'h2)];
              reg86 <= "49Nb8RK";
            end
        end
      reg87 <= ($signed("gD31Y8nbhnii9saD4HA") == $signed(($signed("9Y3rnr0ed4AWcqknL") - $unsigned(forvar77[(4'hb):(3'h5)]))));
    end
  module88 modinst323 (.wire93(reg80), .clk(clk), .wire89(wire70), .wire91(reg85), .wire92(reg81), .y(wire322), .wire90(forvar79));
  assign wire324 = reg82;
  assign wire325 = (^~$signed(reg82));
  module326 modinst658 (.wire328(wire70), .y(wire657), .wire327(reg78), .wire330(wire72), .wire329(reg76), .clk(clk));
  module609 modinst660 (wire659, clk, wire322, forvar77, reg78, wire74, reg85);
  assign wire661 = $unsigned((^~$signed({(forvar84 <<< reg85),
                       (wire71 ^~ reg80)})));
  module326 modinst663 (wire662, clk, wire72, wire659, wire70, wire325);
  assign wire664 = wire75;
  module374 modinst666 (wire665, clk, reg81, wire664, wire70, reg87, wire72);
  assign wire667 = "NqsJ3ES19ParnSxJkIB";
  assign wire668 = (+$unsigned((wire74 <= (7'h41))));
  assign wire669 = ($unsigned(("D4mRsMKY4aGr8xWrU9" | (wire71[(4'ha):(4'h9)] + $unsigned(reg85)))) == reg78[(3'h5):(2'h3)]);
  assign wire670 = reg86[(4'hd):(2'h2)];
  assign wire671 = {$signed((~&$signed($unsigned(wire661))))};
  assign wire672 = forvar84[(2'h3):(1'h0)];
  assign wire673 = ((wire72 & $signed(wire325)) ^~ wire672);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module326
#( parameter param656 = (^~({({(8'had)} ? ((8'ha5) ? (7'h41) : (8'hbe)) : (|(8'h9f))), ((^~(8'hbe)) ? ((7'h43) ~^ (8'hbd)) : (8'hb9))} ? (((-(7'h40)) | (&(8'ha2))) < (((8'hbe) ? (8'hbb) : (8'ha0)) >>> ((8'ha9) + (8'hb2)))) : (~{{(8'hae)}}))) )
(y, clk, wire327, wire328, wire329, wire330);
  output wire [(32'h2a4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire327;
  input wire [(4'h8):(1'h0)] wire328;
  input wire signed [(5'h16):(1'h0)] wire329;
  input wire signed [(5'h13):(1'h0)] wire330;
  wire signed [(2'h2):(1'h0)] wire655;
  wire [(4'hc):(1'h0)] wire654;
  wire signed [(2'h2):(1'h0)] wire653;
  wire [(4'he):(1'h0)] wire652;
  wire [(2'h2):(1'h0)] wire651;
  wire [(3'h4):(1'h0)] wire606;
  wire signed [(5'h11):(1'h0)] wire477;
  reg signed [(4'he):(1'h0)] forvar331 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg332 = (1'h0);
  reg [(4'h9):(1'h0)] reg333 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg334 = (1'h0);
  reg [(5'h12):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg337 = (1'h0);
  reg [(5'h13):(1'h0)] reg338 = (1'h0);
  reg [(5'h14):(1'h0)] reg339 = (1'h0);
  reg [(3'h4):(1'h0)] forvar340 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg341 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg344 = (1'h0);
  reg [(4'hf):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg347 = (1'h0);
  reg [(5'h14):(1'h0)] reg348 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg350 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg351 = (1'h0);
  wire [(2'h3):(1'h0)] wire352;
  wire [(4'h9):(1'h0)] wire353;
  reg signed [(4'hb):(1'h0)] forvar354 = (1'h0);
  reg [(4'he):(1'h0)] forvar355 = (1'h0);
  reg [(5'h12):(1'h0)] reg356 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg357 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire358;
  wire [(3'h5):(1'h0)] wire359;
  wire [(5'h14):(1'h0)] wire360;
  wire [(5'h10):(1'h0)] wire361;
  wire signed [(4'he):(1'h0)] wire362;
  reg signed [(5'h16):(1'h0)] reg363 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg364 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg365 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg366 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg368 = (1'h0);
  reg [(3'h5):(1'h0)] reg369 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg370 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire371;
  wire signed [(4'hf):(1'h0)] wire372;
  wire [(5'h13):(1'h0)] wire373;
  wire signed [(3'h7):(1'h0)] wire475;
  wire [(4'hb):(1'h0)] wire608;
  wire signed [(3'h5):(1'h0)] wire649;
  assign y = {wire655,
                 wire654,
                 wire653,
                 wire652,
                 wire651,
                 wire606,
                 wire477,
                 forvar331,
                 reg332,
                 reg333,
                 reg334,
                 reg335,
                 reg336,
                 reg337,
                 reg338,
                 reg339,
                 forvar340,
                 reg341,
                 reg342,
                 reg343,
                 reg344,
                 reg345,
                 reg346,
                 reg347,
                 reg348,
                 reg349,
                 reg350,
                 reg351,
                 wire352,
                 wire353,
                 forvar354,
                 forvar355,
                 reg356,
                 reg357,
                 wire358,
                 wire359,
                 wire360,
                 wire361,
                 wire362,
                 reg363,
                 reg364,
                 reg365,
                 reg366,
                 reg367,
                 reg368,
                 reg369,
                 reg370,
                 wire371,
                 wire372,
                 wire373,
                 wire475,
                 wire608,
                 wire649,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar331 = (1'h0); (forvar331 < (3'h4)); forvar331 = (forvar331 + (1'h1)))
        begin
          reg332 = $unsigned(($unsigned(wire329) != "iZPPnmie3CNI7KPMSSAM"));
          if ($signed(wire328[(4'h8):(1'h1)]))
            begin
              reg333 <= wire330[(4'hb):(2'h2)];
              reg334 <= ($unsigned($unsigned(reg333)) ?
                  (~|"QcKIJu") : ((~&forvar331[(2'h3):(1'h1)]) ?
                      wire327[(2'h3):(2'h3)] : (($unsigned(wire327) ?
                          $signed((8'ha6)) : $signed(forvar331)) <= forvar331)));
              reg335 <= ((!((-"3") & {(wire328 ? forvar331 : wire329)})) ?
                  (~|$unsigned((&"iJq"))) : (|(+reg333[(1'h1):(1'h1)])));
              reg336 <= ($unsigned((($unsigned(forvar331) <<< (~|(8'ha8))) <<< ((~wire330) >> (&wire328)))) ~^ wire330);
            end
          else
            begin
              reg333 <= (+"EQPHHESUadpKn6wKZo");
              reg334 = ("PgYKq7" <= (reg335 ?
                  (~$signed("fGsMdxuQmiWkNdFrJUs")) : forvar331));
            end
          reg337 = reg336;
        end
      reg338 <= $unsigned(reg335[(1'h0):(1'h0)]);
      if ((wire330 >= $unsigned(reg334)))
        begin
          reg339 <= wire330[(3'h4):(1'h0)];
          for (forvar340 = (1'h0); (forvar340 < (3'h4)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 <= $signed((reg333 >= "SnpNnxJhQf5iHFV"));
              reg342 <= "I4oNCL4lG00vv";
              reg343 = reg332[(4'he):(4'h8)];
              reg344 <= (reg341 == (-$signed("l")));
              reg345 <= "Ns0VYVt5RY5c2gLsP2";
            end
          if ((|(|forvar340[(2'h3):(2'h3)])))
            begin
              reg346 <= reg337[(4'hb):(2'h2)];
              reg347 <= reg332;
              reg348 <= reg345[(4'hf):(3'h5)];
              reg349 <= ((^~"MchLgVIF") ?
                  (!("" < $unsigned({reg345,
                      reg333}))) : $signed({reg339[(2'h2):(1'h0)]}));
              reg350 <= $unsigned($unsigned((^(^~{reg338}))));
            end
          else
            begin
              reg346 = $signed(forvar340);
              reg347 <= (reg343 ?
                  (7'h47) : ((|$signed("5YyMno9BXVVql84o")) ~^ reg341[(2'h3):(1'h1)]));
              reg348 <= reg341[(3'h6):(1'h0)];
              reg349 <= reg348;
              reg350 <= $signed($signed(reg335[(1'h1):(1'h1)]));
            end
        end
      else
        begin
          reg339 <= $unsigned(((~|reg344) ?
              $signed($signed((reg335 ?
                  reg332 : (8'h9d)))) : $signed($signed({reg345, reg348}))));
        end
      reg351 <= $signed({{reg334, $signed($signed(forvar340))}});
    end
  assign wire352 = {reg333};
  assign wire353 = "apzGAQIG14JR6TlxgMmO";
  always
    @(posedge clk) begin
      for (forvar354 = (1'h0); (forvar354 < (1'h1)); forvar354 = (forvar354 + (1'h1)))
        begin
          for (forvar355 = (1'h0); (forvar355 < (1'h1)); forvar355 = (forvar355 + (1'h1)))
            begin
              reg356 <= ($unsigned("K") ?
                  (8'hbb) : ($signed($unsigned(reg337[(3'h4):(1'h0)])) ?
                      {reg333[(1'h0):(1'h0)],
                          $signed((reg347 | wire352))} : (((reg350 >>> (8'hb4)) ?
                              (^reg349) : $unsigned(reg332)) ?
                          ({reg336, reg343} ?
                              "DwlxvuZofIoJOXSmM8Y8Lz" : "7DdWhmPe1fBPA") : reg336)));
            end
        end
      reg357 <= ("tUqZ3" * (~(("D6QF0" ?
          "N445yUvkldP" : (reg349 ?
              wire330 : reg335)) <= ((~|reg347) * (+reg350)))));
    end
  assign wire358 = (&wire329);
  assign wire359 = reg333;
  assign wire360 = ($signed($unsigned(({reg349, reg335} < $signed(reg336)))) ?
                       ($signed(($unsigned(reg339) ?
                               {reg348, reg334} : (wire358 ?
                                   reg343 : reg349))) ?
                           "YuGPsh3hyeSJr1t9gd" : reg342) : (8'ha3));
  assign wire361 = (($unsigned($signed(reg356[(3'h6):(3'h5)])) * (+reg357)) ?
                       $signed(({(reg351 ? wire330 : wire359)} ?
                           $signed($unsigned(reg350)) : reg333)) : reg339);
  assign wire362 = ("0H6H4VFoCKF" - {$signed($unsigned((reg349 << wire327))),
                       $signed("hIw")});
  always
    @(posedge clk) begin
      if ($unsigned($unsigned((((reg336 ? forvar354 : wire353) < {wire327,
          reg345}) | "iNUa7trQtBVGR6VkwqsbB"))))
        begin
          reg363 = ($unsigned(reg342[(4'ha):(3'h7)]) ^~ reg357);
        end
      else
        begin
          reg363 <= reg339;
          if (("WkCU0GDvCIcG4OeV" ?
              (&((&wire329) ?
                  "QCio6DvzvAqfVJvH" : (|(wire360 ?
                      reg333 : reg333)))) : $unsigned((~&"lm1ZgELiW2Igx96y4mV"))))
            begin
              reg364 <= ("9T6PFBH3eRPGl63A8" ?
                  forvar340 : $unsigned((|wire362)));
              reg365 = ((reg351 ?
                  "CnbfDsNakJ" : ($unsigned("rFkAX") >>> $signed((wire352 ?
                      (8'hb4) : (8'ha8))))) >> (-(~($unsigned(wire362) + (forvar354 ?
                  reg339 : reg351)))));
              reg366 <= "JFPm2";
            end
          else
            begin
              reg364 <= ($signed((~&reg332[(3'h6):(2'h3)])) ?
                  ("aopZk738AEa0F0xdM" <= reg344) : (reg332[(3'h6):(1'h1)] ^ forvar340[(1'h0):(1'h0)]));
              reg365 <= reg365[(2'h3):(1'h1)];
              reg366 <= (+"IRsIn");
              reg367 = "1X";
            end
          if ($signed($unsigned(reg351)))
            begin
              reg368 <= ({$signed(""), "vdrQhG0pDkpEy4qd"} ?
                  "u1Ye" : wire361[(1'h1):(1'h0)]);
              reg369 <= $unsigned(($signed("E") ?
                  {"3uxQYtJUWykGaTIuyM5qp"} : $signed(({(7'h46), reg334} ?
                      $signed(reg367) : wire361[(1'h0):(1'h0)]))));
              reg370 <= reg365;
            end
          else
            begin
              reg368 <= reg370;
            end
        end
    end
  assign wire371 = ("o" < (&"k2ovD6P"));
  assign wire372 = reg356[(4'ha):(1'h0)];
  assign wire373 = $signed(("7YWnYWld" ?
                       (~|$unsigned((reg337 ? reg356 : reg367))) : reg335));
  module374 modinst476 (wire475, clk, wire327, reg343, wire362, reg368, reg348);
  assign wire477 = reg345;
  module478 modinst607 (wire606, clk, reg337, reg338, reg346, reg334, wire361);
  assign wire608 = "M0";
  module609 modinst650 (.y(wire649), .wire614(wire359), .wire612(reg332), .wire611(reg370), .clk(clk), .wire610(reg368), .wire613(reg335));
  assign wire651 = $unsigned("9OrhSfJA8HRfN");
  assign wire652 = {((!"4eEQ3CdxZdfSiq") & (|wire359[(1'h1):(1'h0)]))};
  assign wire653 = (reg357[(4'hb):(3'h4)] + ("rLWTDSqlNlZS4PB3yW" ?
                       {"0OqcrT9O005cOG3QZ",
                           ({reg351} ?
                               (wire328 ?
                                   wire330 : wire329) : (~&reg339))} : "TOw9a8aXbU32Wy6MRM"));
  assign wire654 = reg338;
  assign wire655 = $signed(((("IR2unvfgPx5YgmInz" ^ {reg351,
                           reg366}) > ((wire328 * wire373) ~^ (~^wire359))) ?
                       reg351[(1'h0):(1'h0)] : reg344[(5'h11):(3'h6)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module88  (y, clk, wire93, wire92, wire91, wire90, wire89);
  output wire [(32'h253):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire93;
  input wire signed [(5'h10):(1'h0)] wire92;
  input wire signed [(4'hb):(1'h0)] wire91;
  input wire signed [(5'h12):(1'h0)] wire90;
  input wire signed [(5'h13):(1'h0)] wire89;
  reg signed [(3'h6):(1'h0)] reg321 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire320;
  wire signed [(5'h10):(1'h0)] wire319;
  wire [(4'h9):(1'h0)] wire318;
  wire [(4'hb):(1'h0)] wire317;
  wire signed [(4'hc):(1'h0)] wire316;
  wire [(5'h13):(1'h0)] wire314;
  wire [(5'h13):(1'h0)] wire209;
  reg [(3'h7):(1'h0)] reg208 = (1'h0);
  reg [(5'h11):(1'h0)] reg207 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg206 = (1'h0);
  reg [(4'hc):(1'h0)] reg204 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg205 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar204 = (1'h0);
  reg [(5'h12):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg201 = (1'h0);
  reg [(3'h6):(1'h0)] reg200 = (1'h0);
  reg [(4'he):(1'h0)] reg199 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar198 = (1'h0);
  wire [(5'h15):(1'h0)] wire197;
  wire [(5'h17):(1'h0)] wire196;
  reg [(2'h3):(1'h0)] reg195 = (1'h0);
  reg [(5'h10):(1'h0)] reg194 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg193 = (1'h0);
  reg [(4'he):(1'h0)] reg192 = (1'h0);
  reg [(3'h6):(1'h0)] reg191 = (1'h0);
  reg signed [(4'he):(1'h0)] reg190 = (1'h0);
  reg [(4'h9):(1'h0)] reg189 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg188 = (1'h0);
  reg [(4'hb):(1'h0)] reg181 = (1'h0);
  reg [(3'h4):(1'h0)] reg187 = (1'h0);
  reg [(3'h4):(1'h0)] reg186 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg185 = (1'h0);
  reg [(4'he):(1'h0)] reg184 = (1'h0);
  reg signed [(4'he):(1'h0)] reg183 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar181 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg180 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg178 = (1'h0);
  reg [(4'hb):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar176 = (1'h0);
  reg [(2'h2):(1'h0)] reg175 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire174;
  wire signed [(4'ha):(1'h0)] wire172;
  wire [(5'h10):(1'h0)] wire94;
  assign y = {reg321,
                 wire320,
                 wire319,
                 wire318,
                 wire317,
                 wire316,
                 wire314,
                 wire209,
                 reg208,
                 reg207,
                 reg206,
                 reg204,
                 reg198,
                 reg205,
                 forvar204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 forvar198,
                 wire197,
                 wire196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg181,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 forvar181,
                 reg180,
                 reg179,
                 reg176,
                 reg178,
                 reg177,
                 forvar176,
                 reg175,
                 wire174,
                 wire172,
                 wire94,
                 (1'h0)};
  assign wire94 = {{wire89, wire89[(4'ha):(4'ha)]}};
  module95 modinst173 (.wire99(wire92), .wire96(wire91), .wire98(wire93), .y(wire172), .wire97(wire89), .clk(clk));
  assign wire174 = (wire93 < $signed(wire90));
  always
    @(posedge clk) begin
      if (wire174)
        begin
          reg175 <= wire89;
          for (forvar176 = (1'h0); (forvar176 < (1'h0)); forvar176 = (forvar176 + (1'h1)))
            begin
              reg177 <= $signed(wire89);
              reg178 = $unsigned({((reg177[(2'h3):(2'h2)] + $unsigned(wire174)) ?
                      ((&reg177) | (^wire172)) : {wire172})});
            end
        end
      else
        begin
          reg175 <= wire90[(1'h0):(1'h0)];
          if (((+(!"uW5iXEqc")) ?
              "6UC29ptP6XN" : ($signed({{(8'ha1)}}) <<< (wire92[(4'h9):(1'h0)] ?
                  "tV16Xm8pJhbrWZ" : ((wire91 <= wire92) ? "Zo" : {wire90})))))
            begin
              reg176 <= {$unsigned($unsigned($signed($signed((7'h40)))))};
            end
          else
            begin
              reg176 <= (reg176 ?
                  (|"DRzAkIvtMqirnzg") : {{((~^wire90) ?
                              wire174[(4'hb):(1'h1)] : reg176[(4'he):(4'h8)]),
                          $unsigned($unsigned(reg178))},
                      ((wire92[(4'hb):(2'h2)] >= {wire89}) <= "crwf5599awVDGXRfbzz0N")});
              reg177 <= wire93;
            end
          reg178 <= (~"X9K6UcT8Wdyf");
          reg179 <= wire172[(3'h6):(2'h2)];
          reg180 <= (({"", (wire90[(3'h7):(3'h6)] > $unsigned((8'ha5)))} ?
                  $unsigned("8IVsZvBxuAWabi") : ("4NFGx1Tf7cOmwcEqrZs" ?
                      $signed($unsigned(wire91)) : (+(wire89 ~^ (8'ha2))))) ?
              wire91[(3'h7):(2'h2)] : "T");
        end
      if ({($unsigned({"Y5V", $unsigned(wire174)}) ?
              (~|(!wire93)) : $unsigned((wire92 ?
                  {(8'h9c), wire94} : (forvar176 ? wire90 : wire89)))),
          ((($unsigned(wire89) ^~ (forvar176 * reg180)) ?
                  $unsigned(reg177[(1'h0):(1'h0)]) : (!(reg175 ?
                      reg179 : wire172))) ?
              "yxlL3PnVXNztLWwuyttW" : (+(reg176 ?
                  ((7'h41) ? wire94 : reg177) : wire174)))})
        begin
          for (forvar181 = (1'h0); (forvar181 < (2'h3)); forvar181 = (forvar181 + (1'h1)))
            begin
              reg182 <= reg175[(1'h0):(1'h0)];
              reg183 <= (((-(8'ha9)) ?
                      $signed({(+reg177), reg177}) : reg177[(3'h6):(3'h6)]) ?
                  wire92 : wire94);
              reg184 <= "u";
              reg185 <= {reg180[(1'h1):(1'h0)]};
              reg186 <= ("kPLvXkKttNX" || {$signed((8'h9c)), (8'h9c)});
            end
          reg187 <= wire91[(2'h2):(1'h1)];
        end
      else
        begin
          if (((8'ha4) << wire172[(2'h3):(1'h0)]))
            begin
              reg181 <= ((-(~&$signed($signed(reg186)))) - wire94[(1'h1):(1'h0)]);
            end
          else
            begin
              reg181 <= $signed(("9VqRx5EFexenqYOolh" ^ $unsigned(((^forvar176) ?
                  $unsigned(reg180) : {forvar176, (8'ha4)}))));
            end
          if ("uNnyG")
            begin
              reg182 = ($unsigned((~|($unsigned(reg181) ?
                      reg180 : (reg179 < wire93)))) ?
                  ({(reg183 ^~ $unsigned(wire92)),
                      $signed($signed(wire90))} | reg184) : ((8'ha7) >> ($signed((-reg183)) << (^((8'ha9) >>> reg180)))));
              reg183 <= {reg183};
              reg184 <= "Zfsndc2IbBYQo";
            end
          else
            begin
              reg182 <= $unsigned(((reg176 - ((reg180 ?
                  reg185 : reg181) >>> wire90)) * reg175));
            end
          reg185 <= (wire172 >> $signed((wire172[(1'h0):(1'h0)] ?
              ({(8'hb3),
                  reg184} & ((8'hb2) + (8'ha4))) : forvar176[(1'h1):(1'h1)])));
          if ((+reg184[(1'h1):(1'h1)]))
            begin
              reg186 <= "L";
              reg187 <= ((((reg175 ?
                          (wire93 ? reg179 : reg180) : $signed((8'hb7))) ?
                      "wU1PHum81Yzkdx3" : "U") ?
                  ((^~{wire91, wire91}) ?
                      (~^"PeqWNdivXNt") : (reg185 ?
                          "8SHJb2oDWQGMd" : $signed(wire174))) : reg187) & forvar176);
            end
          else
            begin
              reg186 <= "fx9zQCA26LoqtNXt1czB0";
            end
        end
      if (("a" ~^ (reg187 < $signed((~&$signed(forvar181))))))
        begin
          reg188 <= "FFNzHk1kTWAOs5m86";
        end
      else
        begin
          reg188 <= forvar181[(1'h0):(1'h0)];
          if (($signed((!$unsigned($unsigned(reg186)))) << ((|"76Y1UqQLk") ?
              ((reg179 ?
                  $signed(reg176) : (wire94 & reg184)) | ($unsigned(forvar176) >>> reg183[(3'h7):(2'h2)])) : ((+forvar181[(4'hc):(3'h7)]) ?
                  reg188[(2'h3):(1'h0)] : {((8'h9d) ? forvar181 : (8'hba))}))))
            begin
              reg189 <= {{($signed((-wire91)) ^ ((~^reg186) ?
                          (reg184 ? wire93 : reg178) : (forvar176 >= wire92))),
                      (((+reg175) && (~|(8'hb8))) ?
                          {$unsigned(reg184),
                              (^~reg187)} : $signed($unsigned(reg182)))},
                  ($unsigned(((reg185 ? forvar181 : (8'hb9)) ?
                          "JkqeL" : (wire90 - (8'hbc)))) ?
                      "0" : $signed(wire93[(4'ha):(2'h3)]))};
              reg190 <= "kt68fWWUbBetgUEv";
              reg191 <= ((reg181 ?
                      (((8'ha7) ?
                          reg183[(3'h7):(3'h6)] : (~|reg175)) * $signed(reg182[(1'h1):(1'h0)])) : (reg188 ?
                          $unsigned((forvar181 + reg187)) : $unsigned(((7'h42) - wire90)))) ?
                  ($signed((~^(reg180 >> reg188))) ^~ $signed(reg185[(2'h2):(1'h0)])) : ("siEV" == (($unsigned((8'hbf)) ?
                          "uhf8rUgzfM" : $unsigned(wire172)) ?
                      forvar176 : $unsigned((reg177 == wire93)))));
              reg192 <= $unsigned($unsigned("iRZAUwbEbgDuE"));
            end
          else
            begin
              reg189 <= $signed({wire92,
                  {$signed($signed(reg190)),
                      ($signed(reg180) ? (-reg186) : wire172)}});
              reg190 <= reg176;
            end
          reg193 <= $signed({(reg180 ?
                  $unsigned("at46Q94ouLWgNcRnY1Nu") : (7'h48))});
          reg194 <= (reg188 ?
              reg180[(1'h1):(1'h0)] : ((&$unsigned($unsigned(reg184))) ?
                  reg180 : (reg176 ~^ $unsigned($unsigned((8'ha4))))));
        end
      reg195 <= $unsigned(($signed(reg194[(4'hf):(3'h4)]) ?
          reg177[(4'ha):(1'h0)] : reg188));
    end
  assign wire196 = {($signed(reg179[(1'h1):(1'h0)]) ? "3Z" : (~&wire92)),
                       $unsigned({($signed(reg181) ?
                               (&reg180) : $signed(wire92))})};
  assign wire197 = ($unsigned(forvar176) & ("E5ZvIJstbWoRv96dBIoRUK" >>> (~|reg175[(1'h1):(1'h1)])));
  always
    @(posedge clk) begin
      if ("1bA")
        begin
          for (forvar198 = (1'h0); (forvar198 < (1'h0)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 <= (reg183 >>> "c6V81Phy1H7JeX");
              reg200 <= $signed($unsigned(reg192));
              reg201 <= (forvar176[(4'h8):(3'h6)] ?
                  $unsigned("4qaPtQOsvJn") : reg195[(2'h2):(1'h0)]);
              reg202 <= (+(reg200 || reg199));
              reg203 = reg175[(1'h0):(1'h0)];
            end
          for (forvar204 = (1'h0); (forvar204 < (1'h0)); forvar204 = (forvar204 + (1'h1)))
            begin
              reg205 <= $unsigned($signed(""));
            end
        end
      else
        begin
          if ((|(+{$unsigned({(8'hb2)}),
              (reg187[(2'h2):(2'h2)] >> "NuEXXxNmQyF")})))
            begin
              reg198 <= $signed((~{((~|forvar181) << reg176),
                  reg192[(1'h1):(1'h0)]}));
              reg199 <= $unsigned(($unsigned(((forvar181 || (8'ha0)) <<< wire92[(4'hb):(2'h2)])) > ($signed($signed((8'hac))) + (reg200[(1'h1):(1'h1)] | forvar198[(3'h7):(3'h5)]))));
              reg200 = (reg188[(1'h0):(1'h0)] | (($unsigned((reg180 ?
                      (8'hae) : forvar181)) ?
                  $unsigned(reg203[(4'ha):(1'h1)]) : "txtFnLSSBMeHaJLkVa5F") >= (~{reg193})));
              reg201 <= ("gTx1" >> (!((~|{reg201, (7'h45)}) <<< ({wire93,
                  reg193} <<< (reg188 ^ reg198)))));
              reg202 <= "nIgSLfnwy4fgSVgfBZZ";
            end
          else
            begin
              reg198 <= "KNL";
              reg199 <= (&reg190);
              reg200 <= reg183[(4'hb):(4'hb)];
              reg201 <= reg194;
              reg202 <= $signed($signed($signed(reg192[(2'h2):(2'h2)])));
            end
          if ("3S")
            begin
              reg203 <= "ZcKYZFBC";
            end
          else
            begin
              reg203 <= (|(reg184 ? (~^"zs95rPLSpnomF") : (8'hbf)));
              reg204 = (~^($unsigned({(reg187 >= reg178),
                      reg205[(5'h13):(5'h13)]}) ?
                  $unsigned(forvar176[(1'h1):(1'h1)]) : (&{{reg177}})));
              reg205 <= ((wire93[(4'h8):(2'h3)] - (wire92 ?
                  $signed($unsigned(wire91)) : ((reg184 ? reg178 : reg190) ?
                      $signed(wire92) : "8NiUtOKbScoSwtdDBGZpc"))) >>> (^~(|reg191[(3'h5):(3'h4)])));
            end
        end
      reg206 <= $unsigned("c9aEuRJy");
      reg207 <= (wire197[(3'h6):(2'h3)] >>> (~(!"Blbi6pCuGzs")));
      reg208 <= "7A7aawE";
    end
  assign wire209 = reg182[(2'h3):(2'h3)];
  module210 modinst315 (wire314, clk, reg192, reg190, reg205, reg201);
  assign wire316 = (8'hb8);
  assign wire317 = reg180[(1'h1):(1'h1)];
  assign wire318 = "Iv3Cuw";
  assign wire319 = (reg176[(1'h0):(1'h0)] ? $signed($signed(reg195)) : (7'h47));
  assign wire320 = {$unsigned(reg199),
                       ($signed((~&(wire314 ?
                           reg177 : reg178))) > (^~(reg177[(3'h7):(1'h1)] < $unsigned(wire89))))};
  always
    @(posedge clk) begin
      reg321 <= reg178[(4'hf):(4'hb)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module210
#( parameter param313 = ((((~&((8'hb6) ? (8'hbb) : (8'ha4))) >>> (((8'ha0) ? (8'haf) : (8'haa)) ? (~&(8'h9e)) : ((7'h40) > (7'h41)))) ? ((!((7'h40) + (8'ha0))) && {((7'h44) ? (8'h9e) : (7'h46)), {(7'h45)}}) : ((-(|(7'h42))) ^~ (^((7'h46) != (8'hb3))))) ? ((({(8'ha7)} > {(8'ha9)}) ? (~^(8'ha7)) : (((8'h9f) <<< (8'ha9)) == ((8'hb6) & (8'hbc)))) ? (+((^(8'had)) ^ ((8'hb1) ? (8'ha7) : (8'hbc)))) : ((((8'hb3) <<< (8'hab)) ? (^(7'h43)) : ((8'hb9) ? (8'hba) : (8'hbd))) << (((8'hb2) == (8'ha9)) || ((8'hae) ~^ (7'h43))))) : (&{((~^(8'hb8)) ? ((8'hb8) || (8'ha5)) : (+(8'ha1))), ((^~(8'ha9)) ? ((7'h43) - (8'haf)) : ((8'hb9) ? (8'hba) : (8'hb4)))})) )
(y, clk, wire214, wire213, wire212, wire211);
  output wire [(32'h4c9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire214;
  input wire signed [(3'h7):(1'h0)] wire213;
  input wire signed [(4'hd):(1'h0)] wire212;
  input wire [(5'h10):(1'h0)] wire211;
  wire [(3'h5):(1'h0)] wire312;
  wire [(4'h8):(1'h0)] wire311;
  wire [(4'h9):(1'h0)] wire310;
  wire [(3'h4):(1'h0)] wire309;
  wire signed [(4'hf):(1'h0)] wire308;
  wire signed [(3'h6):(1'h0)] wire307;
  reg signed [(5'h12):(1'h0)] reg306 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar305 = (1'h0);
  reg [(4'hc):(1'h0)] reg304 = (1'h0);
  reg [(5'h16):(1'h0)] reg303 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar302 = (1'h0);
  reg [(4'h8):(1'h0)] forvar301 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg300 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg299 = (1'h0);
  wire signed [(5'h16):(1'h0)] wire298;
  wire [(3'h5):(1'h0)] wire297;
  wire [(4'ha):(1'h0)] wire296;
  wire signed [(3'h7):(1'h0)] wire295;
  wire signed [(3'h4):(1'h0)] wire294;
  wire signed [(4'he):(1'h0)] wire293;
  wire [(2'h3):(1'h0)] wire292;
  wire signed [(4'h9):(1'h0)] wire291;
  reg signed [(5'h12):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar276 = (1'h0);
  reg [(4'h8):(1'h0)] reg290 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg289 = (1'h0);
  reg [(5'h14):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar286 = (1'h0);
  reg [(5'h14):(1'h0)] reg285 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg284 = (1'h0);
  reg [(4'ha):(1'h0)] reg283 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg281 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar280 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg278 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar277 = (1'h0);
  reg [(4'h8):(1'h0)] reg276 = (1'h0);
  reg [(3'h6):(1'h0)] reg275 = (1'h0);
  reg signed [(4'he):(1'h0)] reg274 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg272 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg271 = (1'h0);
  reg [(3'h7):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg269 = (1'h0);
  reg [(4'he):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar267 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg266 = (1'h0);
  reg [(5'h12):(1'h0)] reg265 = (1'h0);
  reg [(5'h16):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar262 = (1'h0);
  reg [(3'h4):(1'h0)] reg261 = (1'h0);
  reg [(2'h2):(1'h0)] reg260 = (1'h0);
  reg [(4'hc):(1'h0)] reg259 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg258 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg256 = (1'h0);
  reg [(3'h6):(1'h0)] reg255 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg254 = (1'h0);
  reg [(4'hf):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg252 = (1'h0);
  reg [(2'h3):(1'h0)] reg251 = (1'h0);
  reg [(5'h14):(1'h0)] forvar250 = (1'h0);
  wire [(3'h7):(1'h0)] wire249;
  wire signed [(5'h15):(1'h0)] wire248;
  wire [(3'h6):(1'h0)] wire247;
  wire [(4'h8):(1'h0)] wire246;
  wire signed [(5'h14):(1'h0)] wire245;
  wire signed [(4'hb):(1'h0)] wire244;
  reg [(2'h3):(1'h0)] reg243 = (1'h0);
  reg [(3'h5):(1'h0)] reg242 = (1'h0);
  reg [(5'h11):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar240 = (1'h0);
  reg [(4'ha):(1'h0)] reg239 = (1'h0);
  reg [(5'h14):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg237 = (1'h0);
  reg [(4'h9):(1'h0)] reg236 = (1'h0);
  reg [(5'h16):(1'h0)] reg235 = (1'h0);
  reg [(4'hb):(1'h0)] forvar234 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg233 = (1'h0);
  reg [(4'ha):(1'h0)] reg232 = (1'h0);
  reg [(3'h7):(1'h0)] forvar231 = (1'h0);
  wire [(5'h15):(1'h0)] wire230;
  reg [(5'h10):(1'h0)] reg229 = (1'h0);
  reg [(4'hd):(1'h0)] reg228 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg227 = (1'h0);
  reg [(5'h12):(1'h0)] forvar226 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg224 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg223 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg222 = (1'h0);
  reg [(4'hd):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar220 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg219 = (1'h0);
  reg [(4'hb):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg217 = (1'h0);
  reg [(4'he):(1'h0)] reg216 = (1'h0);
  reg [(3'h4):(1'h0)] reg215 = (1'h0);
  assign y = {wire312,
                 wire311,
                 wire310,
                 wire309,
                 wire308,
                 wire307,
                 reg306,
                 forvar305,
                 reg304,
                 reg303,
                 forvar302,
                 forvar301,
                 reg300,
                 reg299,
                 wire298,
                 wire297,
                 wire296,
                 wire295,
                 wire294,
                 wire293,
                 wire292,
                 wire291,
                 reg277,
                 forvar276,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 forvar286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 forvar280,
                 reg279,
                 reg278,
                 forvar277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 forvar267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 forvar262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 forvar250,
                 wire249,
                 wire248,
                 wire247,
                 wire246,
                 wire245,
                 wire244,
                 reg243,
                 reg242,
                 reg241,
                 forvar240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 forvar234,
                 reg233,
                 reg232,
                 forvar231,
                 wire230,
                 reg229,
                 reg228,
                 reg227,
                 forvar226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 forvar220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire211[(4'hc):(4'hc)])
        begin
          reg215 <= "K1Xh";
          reg216 <= (wire214 ? (!"Edr") : $signed($unsigned((^(~|wire212)))));
          if ((8'haa))
            begin
              reg217 = "z7mwzNPK3tfSrmUZ8YA";
            end
          else
            begin
              reg217 = "D4VYENDCOuyMtIgLxxp";
            end
          reg218 <= "P7pLm";
        end
      else
        begin
          if ((7'h43))
            begin
              reg215 <= {$signed({wire212[(1'h1):(1'h1)],
                      $signed((~^wire213))}),
                  $unsigned(reg216[(2'h3):(2'h2)])};
              reg216 <= {$signed("b1yslI1QzsImHRIWkBy94a"),
                  $unsigned(reg216[(1'h1):(1'h1)])};
              reg217 <= $unsigned((wire212[(4'h9):(1'h1)] != $signed(((reg216 && reg215) ?
                  $signed(reg217) : $signed(wire212)))));
            end
          else
            begin
              reg215 = "t2ZuF8qvIABd9hBVO";
              reg216 <= $unsigned({wire211[(3'h6):(1'h0)],
                  reg216[(4'he):(4'hc)]});
              reg217 = "kegRu8PN3";
              reg218 <= (("BuUlg" + ((~|(+wire211)) ?
                  (^~{(8'ha9), (8'hae)}) : (((8'ha1) ? reg217 : (8'h9e)) ?
                      "2We" : "a66vK9IhMUVi4VDKdJNAt"))) - reg216);
              reg219 <= reg215;
            end
        end
      for (forvar220 = (1'h0); (forvar220 < (2'h2)); forvar220 = (forvar220 + (1'h1)))
        begin
          reg221 <= ((wire213 + wire212[(1'h0):(1'h0)]) ~^ $unsigned((~|($unsigned((8'ha7)) >> "fa6BG2MbdxWmXozdqw"))));
          if ($signed(wire214))
            begin
              reg222 <= (-({("7p6V95wHuv0H" ?
                      (reg219 ? reg218 : reg217) : (wire214 ?
                          reg221 : wire212)),
                  ((reg217 < wire211) << $signed(reg215))} ^~ "qX9TqzSFgvRsBLA"));
              reg223 <= $signed((~((|$unsigned(wire212)) >> ($signed(reg221) > $unsigned(wire212)))));
              reg224 <= "eWL";
            end
          else
            begin
              reg222 <= ((!reg222[(1'h0):(1'h0)]) ?
                  (({(~&reg219), reg219[(1'h0):(1'h0)]} >>> {(reg224 < wire212),
                          ((8'ha7) ^~ (8'hb6))}) ?
                      reg221[(4'h8):(3'h5)] : {{(wire212 >= reg218),
                              $unsigned((8'hb6))}}) : $signed((reg223[(4'h9):(3'h5)] ?
                      (reg219[(1'h0):(1'h0)] ?
                          $signed(forvar220) : "JR") : ((8'hb5) ?
                          $signed(forvar220) : forvar220))));
            end
          reg225 <= ($unsigned(forvar220[(4'h8):(1'h1)]) ? reg222 : (|wire212));
          for (forvar226 = (1'h0); (forvar226 < (3'h4)); forvar226 = (forvar226 + (1'h1)))
            begin
              reg227 <= $unsigned("y0x");
              reg228 <= "VJcHlrZCP1Jn4BynWbU";
            end
          reg229 <= $signed({(7'h45), "3G551SKYqYv4ddlnO"});
        end
    end
  assign wire230 = reg224[(4'h8):(3'h6)];
  always
    @(posedge clk) begin
      for (forvar231 = (1'h0); (forvar231 < (1'h1)); forvar231 = (forvar231 + (1'h1)))
        begin
          reg232 <= (-(!$unsigned((reg224 ?
              forvar231 : {wire213, forvar231}))));
          reg233 <= forvar226;
          for (forvar234 = (1'h0); (forvar234 < (2'h2)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 = "rafgNTYdQ1tXo";
              reg236 = (({reg225,
                      (reg233 ? $unsigned(reg228) : reg215[(2'h3):(1'h0)])} ?
                  (((forvar226 ? reg224 : reg221) ?
                      wire230[(1'h0):(1'h0)] : $signed(reg215)) * reg222[(4'h9):(3'h6)]) : $signed("fnGwWE")) || "Y");
              reg237 <= $signed($unsigned((&reg222[(4'h9):(2'h3)])));
              reg238 <= (($unsigned(reg217) ?
                  $signed($unsigned("lUQ")) : reg224) | ({("dVPmkV" ^~ $signed(reg228)),
                      $signed(reg219)} ?
                  "gH" : (8'ha2)));
              reg239 <= (~&$signed(wire213[(2'h2):(1'h0)]));
            end
          for (forvar240 = (1'h0); (forvar240 < (3'h4)); forvar240 = (forvar240 + (1'h1)))
            begin
              reg241 <= $signed((8'had));
              reg242 <= reg229[(4'ha):(1'h1)];
              reg243 <= $signed((reg223[(2'h3):(2'h3)] ?
                  ((reg219[(2'h2):(1'h1)] ?
                      $signed(reg224) : $signed(reg224)) ^~ (-(reg217 >= reg215))) : (~^"pg1VzDAmFgf")));
            end
        end
    end
  assign wire244 = (^(^$unsigned($signed({reg228, reg227}))));
  assign wire245 = $signed("oIctixa09mrvN2B7wB9iT5");
  assign wire246 = forvar234;
  assign wire247 = ((!$unsigned("")) ^ "PdISXT1rvOrKWHGtbJvK4");
  assign wire248 = "00m1IOvlyxg";
  assign wire249 = (({(!"DoPm9JV8z9G"), (8'hab)} ?
                       $signed(wire246[(3'h5):(2'h3)]) : (reg243[(1'h0):(1'h0)] ?
                           "AYeqV0MEY" : $unsigned((|wire214)))) < {"YXooEHl",
                       $unsigned($unsigned(reg215[(2'h2):(1'h0)]))});
  always
    @(posedge clk) begin
      for (forvar250 = (1'h0); (forvar250 < (1'h1)); forvar250 = (forvar250 + (1'h1)))
        begin
          reg251 <= $signed(wire213);
          reg252 <= $unsigned(({reg216[(3'h7):(3'h6)]} ?
              $signed(reg219[(2'h2):(2'h2)]) : $unsigned($signed($signed(reg232)))));
          if (reg237)
            begin
              reg253 <= (wire230[(5'h13):(3'h4)] ?
                  (~^$signed((-(reg233 ? (8'had) : reg222)))) : reg252);
              reg254 <= "WWvP";
              reg255 <= $signed($signed((~|((reg235 || reg243) ^ $unsigned((8'h9c))))));
              reg256 <= $unsigned(reg233);
              reg257 <= (forvar220 && $unsigned("yLsEu0kHnxmLRM0p94LRPa"));
            end
          else
            begin
              reg253 <= (($unsigned(forvar250) >>> (wire212[(2'h3):(1'h1)] ^ reg257)) > "7Q4d7TKPsmTR4g");
              reg254 <= ($unsigned($unsigned(reg253[(4'hb):(4'h9)])) ?
                  {{$unsigned(reg253[(4'hf):(2'h3)])}} : wire213);
              reg255 <= {forvar231[(3'h7):(3'h4)], "IOH9CL1"};
              reg256 <= reg229[(1'h0):(1'h0)];
              reg257 <= $signed("pE0okn3wL");
            end
          if ($signed("d2AerQWB8RUMbZdy0"))
            begin
              reg258 <= reg229[(2'h3):(1'h1)];
              reg259 <= reg241[(3'h6):(3'h4)];
              reg260 <= $unsigned(($unsigned("KQ86LWeq8Vi") ?
                  reg258[(3'h4):(2'h3)] : $signed("tye4XpDpbwNo")));
              reg261 <= {((&wire212[(3'h5):(1'h1)]) ?
                      ($unsigned($signed(reg260)) ?
                          {reg215[(1'h0):(1'h0)],
                              "uk27X0F"} : reg216) : (reg238 || (8'hb4))),
                  $unsigned((($unsigned(reg241) ?
                      (reg235 << reg237) : $unsigned(wire249)) + (8'hbb)))};
            end
          else
            begin
              reg258 <= ($signed($signed("mvciTpWPY9dWL")) ^ "p4twwv");
              reg259 <= forvar240;
              reg260 <= reg223;
            end
        end
      if ($signed(($signed($unsigned((wire247 ? reg218 : reg243))) ?
          "oM1dJ27EkTMAb4O6hKuYK" : reg238)))
        begin
          for (forvar262 = (1'h0); (forvar262 < (2'h3)); forvar262 = (forvar262 + (1'h1)))
            begin
              reg263 = "";
              reg264 <= ((~wire245) ?
                  "Wk" : $unsigned((wire248[(2'h3):(1'h0)] | reg224[(5'h10):(2'h3)])));
              reg265 <= "bbi6YbM93csZHV3QuB6v2";
              reg266 <= wire248[(4'hf):(4'h9)];
            end
          for (forvar267 = (1'h0); (forvar267 < (1'h1)); forvar267 = (forvar267 + (1'h1)))
            begin
              reg268 <= forvar250[(1'h1):(1'h1)];
            end
          reg269 <= (8'hb4);
          if (((8'hbc) ?
              {(!$signed($unsigned(reg251))), reg255} : ($signed(reg227) ?
                  "QtgTsttqGsxf" : reg222)))
            begin
              reg270 <= $signed((|$unsigned((+reg258))));
              reg271 <= (~|reg242[(1'h0):(1'h0)]);
              reg272 <= $unsigned("");
              reg273 <= ($unsigned(reg258) ?
                  "PGbX7TGC0JincsIKvN" : (wire244 ~^ forvar262));
            end
          else
            begin
              reg270 <= $signed(reg263[(4'hb):(3'h7)]);
              reg271 <= reg218[(3'h5):(2'h2)];
            end
        end
      else
        begin
          for (forvar262 = (1'h0); (forvar262 < (2'h3)); forvar262 = (forvar262 + (1'h1)))
            begin
              reg263 <= {{$unsigned({$unsigned(reg241)})}};
              reg264 <= "1";
              reg265 <= (reg233 ? "KQYHzIx9ZQTsInMU" : (+$unsigned(wire213)));
            end
          reg266 <= (($unsigned($unsigned($unsigned(reg268))) ?
                  $signed($signed($unsigned(forvar267))) : ("WgNB2LXmXgKCRreI80q" ?
                      reg219 : "1rY8VR9LTV5g3vZhKvPRsu")) ?
              (^$unsigned(reg258)) : $signed(reg256[(4'hd):(4'hc)]));
          for (forvar267 = (1'h0); (forvar267 < (1'h1)); forvar267 = (forvar267 + (1'h1)))
            begin
              reg268 <= {({$signed((+reg257)), "9A2k4bGP69w8gCNTRJO3"} | "wS"),
                  ((reg235[(3'h4):(1'h0)] ?
                      $signed((wire249 ?
                          forvar220 : (8'hba))) : {$unsigned(reg217)}) == {{$signed(reg263),
                          forvar240[(5'h11):(4'hd)]}})};
              reg269 <= "vH6hM7d0vVeEPP1JW";
              reg270 = $signed((("QUgt" < {(8'ha5)}) ?
                  wire230 : $signed(reg258)));
              reg271 <= "7qqiCFeyO";
              reg272 <= reg272;
            end
          reg273 <= reg235;
          reg274 <= (8'hb1);
        end
      if ("2I7V6rv3gdGAVqMPuYYq8")
        begin
          if ((((reg223 ?
                  "Wgmm3MPfh" : ((reg221 >>> (8'hbf)) < reg239[(2'h3):(2'h2)])) & ({(~|reg225),
                      $unsigned(reg242)} ?
                  reg274 : reg227)) ?
              reg233 : ((+$signed((~^reg219))) <= (~^$signed(reg241)))))
            begin
              reg275 <= reg223[(3'h7):(1'h1)];
              reg276 <= ($unsigned("Ux") ? reg233 : $unsigned((~&"Znyy12vg")));
            end
          else
            begin
              reg275 <= ((forvar262 >= $signed((~^((8'ha8) ?
                      wire211 : reg251)))) ?
                  $signed((^($signed(wire248) ?
                      "d5eoKDoO0Xibf6pQpT" : reg223))) : (reg218[(4'hb):(4'ha)] ^ ("qEVw29G6B" ^~ reg274[(2'h2):(1'h1)])));
              reg276 <= $unsigned(((((~|reg253) ~^ {reg227}) ?
                  $signed((wire230 ?
                      reg225 : (8'hbd))) : (~reg269[(3'h4):(1'h1)])) >>> $signed((-$unsigned(forvar262)))));
            end
          for (forvar277 = (1'h0); (forvar277 < (2'h2)); forvar277 = (forvar277 + (1'h1)))
            begin
              reg278 <= reg232[(2'h3):(1'h1)];
              reg279 <= reg242;
            end
          for (forvar280 = (1'h0); (forvar280 < (1'h0)); forvar280 = (forvar280 + (1'h1)))
            begin
              reg281 <= ($unsigned($signed("vi")) * (+reg261));
              reg282 <= "JHcUmX";
              reg283 <= $signed(forvar240);
              reg284 <= {(8'hb0), "UzL"};
              reg285 <= ($unsigned(reg264[(4'h9):(2'h3)]) ?
                  $unsigned((~^$unsigned((reg278 && reg223)))) : ("SyHn2ee9rm6Q2" + (reg282[(3'h6):(3'h6)] >= reg228)));
            end
          for (forvar286 = (1'h0); (forvar286 < (1'h1)); forvar286 = (forvar286 + (1'h1)))
            begin
              reg287 <= reg283[(1'h0):(1'h0)];
              reg288 <= reg227;
              reg289 <= reg261[(1'h1):(1'h1)];
              reg290 <= ($unsigned(reg225[(4'h9):(3'h5)]) ?
                  ($unsigned(((reg223 ? wire248 : forvar250) ?
                      ((8'hbe) ?
                          reg242 : forvar226) : reg253[(2'h3):(1'h1)])) <<< ($unsigned((~^reg288)) * reg268[(4'hd):(3'h7)])) : $unsigned(reg236));
            end
        end
      else
        begin
          reg275 = reg223;
          for (forvar276 = (1'h0); (forvar276 < (1'h0)); forvar276 = (forvar276 + (1'h1)))
            begin
              reg277 <= {({reg290,
                      ({wire249, reg242} ?
                          (reg269 || reg271) : {reg290})} <<< ("2gaRU8Zvx" ?
                      reg241[(4'hc):(3'h7)] : {"ETmAb1LGq9OVKyakAex"}))};
              reg278 = (($signed($unsigned((reg253 ?
                  (8'ha9) : reg227))) >= ((((7'h46) ?
                      forvar250 : reg273) || $unsigned(reg284)) ?
                  $signed("JVXA") : "WXheKJKmeSR")) <= reg277);
            end
        end
    end
  assign wire291 = {forvar280, (^~(^~((~|reg284) <= (~&reg238))))};
  assign wire292 = $unsigned($signed((((~reg242) > (reg223 | reg289)) ?
                       ((~forvar231) >> reg279[(2'h2):(2'h2)]) : {$signed(forvar250),
                           forvar240})));
  assign wire293 = ($unsigned($unsigned(wire212)) ^~ (!$unsigned($unsigned($unsigned(reg285)))));
  assign wire294 = $signed((~|$unsigned(((8'hba) ?
                       $signed(reg283) : (7'h46)))));
  assign wire295 = wire246[(3'h6):(1'h1)];
  assign wire296 = (~^{(~^(^wire295[(1'h0):(1'h0)])), reg270});
  assign wire297 = $unsigned("oJkiSGx92oDidhfbPBRP");
  assign wire298 = $unsigned($signed((~|$unsigned((reg268 ~^ (8'hbd))))));
  always
    @(posedge clk) begin
      reg299 <= (reg255[(2'h3):(1'h0)] <= ((("Cxu10TuFu6T9M49PBN" ?
              ((8'hbc) ? wire291 : reg285) : {wire245, (7'h46)}) ?
          forvar220 : ((wire295 - reg289) ?
              (reg243 ?
                  reg238 : wire296) : reg239)) > $unsigned(("JqROwEhv9gfn" || (forvar277 ~^ reg290)))));
      reg300 <= ($signed("1aLWdBvWoz4JKe") ?
          reg263 : (reg283 ?
              "CGr8oCR19q7glrei" : (^~$unsigned($signed(reg281)))));
      for (forvar301 = (1'h0); (forvar301 < (1'h1)); forvar301 = (forvar301 + (1'h1)))
        begin
          for (forvar302 = (1'h0); (forvar302 < (2'h3)); forvar302 = (forvar302 + (1'h1)))
            begin
              reg303 <= reg229;
            end
          reg304 = (((~^wire230) ?
                  (("e7NxO" ~^ {reg253}) - reg253[(1'h0):(1'h0)]) : $unsigned($signed("6SNEF"))) ?
              $signed(("7UEZRVqAnhvg" ?
                  $signed((^reg281)) : "D2QYQL3I24fDKWeq8iz")) : {(forvar301[(2'h2):(1'h0)] ?
                      (&(reg251 != reg255)) : $signed((reg225 << reg288)))});
        end
      for (forvar305 = (1'h0); (forvar305 < (2'h3)); forvar305 = (forvar305 + (1'h1)))
        begin
          reg306 <= "DCe0vJt02aB6FKN3Ix";
        end
    end
  assign wire307 = forvar286;
  assign wire308 = "5TnVBU0FzCca84TfkoAW";
  assign wire309 = ($signed((reg279[(2'h2):(2'h2)] ?
                           forvar262 : "KPFemAW5AqJarcYTU1")) ?
                       (+wire308) : "VT5CrVU5l6NP");
  assign wire310 = $signed($signed(reg269));
  assign wire311 = (|$signed($unsigned($unsigned($unsigned((8'had))))));
  assign wire312 = $signed($unsigned((reg281[(4'hc):(3'h6)] < $unsigned((reg223 ~^ forvar302)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module95
#( parameter param171 = (~^(-((^{(7'h40), (8'hb1)}) * ((|(8'had)) << ((8'hb3) != (8'hba)))))) )
(y, clk, wire99, wire98, wire97, wire96);
  output wire [(32'h3a4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire99;
  input wire signed [(4'h8):(1'h0)] wire98;
  input wire signed [(5'h10):(1'h0)] wire97;
  input wire [(4'hb):(1'h0)] wire96;
  wire [(3'h5):(1'h0)] wire170;
  wire signed [(4'hb):(1'h0)] wire169;
  wire [(4'h9):(1'h0)] wire168;
  reg [(2'h2):(1'h0)] reg167 = (1'h0);
  reg [(4'ha):(1'h0)] reg166 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg165 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar163 = (1'h0);
  reg [(4'hd):(1'h0)] reg148 = (1'h0);
  reg [(4'hb):(1'h0)] forvar146 = (1'h0);
  reg [(5'h14):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg161 = (1'h0);
  reg [(3'h7):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg159 = (1'h0);
  reg [(2'h3):(1'h0)] reg158 = (1'h0);
  reg [(5'h10):(1'h0)] reg157 = (1'h0);
  reg [(5'h17):(1'h0)] reg156 = (1'h0);
  reg [(5'h10):(1'h0)] reg155 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg154 = (1'h0);
  reg [(3'h4):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar152 = (1'h0);
  reg [(5'h15):(1'h0)] reg151 = (1'h0);
  reg [(2'h3):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg149 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar148 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg147 = (1'h0);
  reg [(3'h4):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg144 = (1'h0);
  reg [(5'h14):(1'h0)] reg143 = (1'h0);
  reg [(5'h12):(1'h0)] reg142 = (1'h0);
  reg [(5'h10):(1'h0)] forvar141 = (1'h0);
  reg [(3'h7):(1'h0)] reg140 = (1'h0);
  reg [(4'hb):(1'h0)] reg139 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar138 = (1'h0);
  wire [(4'hf):(1'h0)] wire137;
  wire [(5'h10):(1'h0)] wire136;
  wire [(5'h11):(1'h0)] wire135;
  wire signed [(4'ha):(1'h0)] wire134;
  wire [(4'h9):(1'h0)] wire133;
  wire signed [(4'hc):(1'h0)] wire132;
  wire signed [(3'h4):(1'h0)] wire131;
  reg [(4'hd):(1'h0)] reg130 = (1'h0);
  reg [(5'h16):(1'h0)] reg129 = (1'h0);
  reg [(5'h10):(1'h0)] reg128 = (1'h0);
  reg [(5'h10):(1'h0)] reg127 = (1'h0);
  reg [(4'hc):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg106 = (1'h0);
  reg [(4'h8):(1'h0)] reg125 = (1'h0);
  reg [(2'h2):(1'h0)] reg124 = (1'h0);
  reg [(5'h10):(1'h0)] reg123 = (1'h0);
  reg [(5'h15):(1'h0)] reg122 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar120 = (1'h0);
  reg [(4'h8):(1'h0)] reg119 = (1'h0);
  reg [(4'h9):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar117 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg114 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg113 = (1'h0);
  reg signed [(4'he):(1'h0)] reg112 = (1'h0);
  reg [(3'h7):(1'h0)] reg111 = (1'h0);
  reg [(5'h16):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg108 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar106 = (1'h0);
  reg [(2'h3):(1'h0)] reg105 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire104;
  wire [(5'h14):(1'h0)] wire103;
  wire [(4'ha):(1'h0)] wire102;
  wire [(5'h15):(1'h0)] wire101;
  wire [(5'h11):(1'h0)] wire100;
  assign y = {wire170,
                 wire169,
                 wire168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 forvar163,
                 reg148,
                 forvar146,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 forvar152,
                 reg151,
                 reg150,
                 reg149,
                 forvar148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 forvar141,
                 reg140,
                 reg139,
                 forvar138,
                 wire137,
                 wire136,
                 wire135,
                 wire134,
                 wire133,
                 wire132,
                 wire131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg106,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 forvar120,
                 reg119,
                 reg118,
                 forvar117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 forvar106,
                 reg105,
                 wire104,
                 wire103,
                 wire102,
                 wire101,
                 wire100,
                 (1'h0)};
  assign wire100 = $unsigned(($unsigned(((8'ha9) ?
                       (wire96 | wire97) : $signed(wire97))) >> ("Qtq51OkUP" ?
                       ("dEd0O40TNxpyQ8s" ^~ wire98[(4'h8):(3'h7)]) : ({wire99,
                           wire97} <<< $signed(wire96)))));
  assign wire101 = $signed($signed((|wire99[(1'h0):(1'h0)])));
  assign wire102 = (|({{$unsigned(wire98)}, wire101[(4'hc):(4'ha)]} ?
                       (((~|wire97) ?
                               wire101[(5'h13):(5'h12)] : $signed(wire96)) ?
                           $signed((7'h48)) : wire100) : "Ar2E665o1dAvkvQU7yhye"));
  assign wire103 = ("NwErBy" <<< ((wire98 ?
                           $unsigned((wire98 ?
                               wire98 : wire101)) : {$signed(wire101),
                               (wire99 >> wire98)}) ?
                       $unsigned(($unsigned((8'hb2)) ~^ wire97[(2'h2):(2'h2)])) : {$signed(wire101[(2'h3):(2'h3)]),
                           wire96[(4'ha):(4'h9)]}));
  assign wire104 = "";
  always
    @(posedge clk) begin
      reg105 <= wire98[(4'h8):(3'h4)];
      if ($signed("FdW9"))
        begin
          for (forvar106 = (1'h0); (forvar106 < (1'h1)); forvar106 = (forvar106 + (1'h1)))
            begin
              reg107 = "Pl6dM0oJ";
              reg108 = wire104;
              reg109 <= forvar106[(4'h9):(3'h5)];
              reg110 = {($unsigned($unsigned(wire96)) >>> wire104),
                  {wire99,
                      (reg105[(1'h0):(1'h0)] >> $unsigned("wXB8R0JVGLGl7Q0cfYO"))}};
              reg111 <= "BBIoApbaxBhqA7xDipQ";
            end
          if ($unsigned((~|($signed(reg111) ?
              (~(~^wire97)) : wire101[(5'h14):(5'h12)]))))
            begin
              reg112 = $unsigned(wire98[(4'h8):(2'h3)]);
              reg113 <= (forvar106[(4'hb):(4'hb)] ?
                  (8'haa) : ("PkOiuy9PBtMztGY" ?
                      ($unsigned((reg109 ? wire103 : wire98)) ?
                          ("6Y" >> (reg112 >= reg108)) : wire98[(2'h3):(2'h2)]) : $unsigned((~&wire102[(3'h5):(2'h3)]))));
            end
          else
            begin
              reg112 <= (reg108[(4'hb):(1'h1)] << ("GaC" ?
                  wire100[(4'hf):(4'h8)] : ($unsigned($signed(wire104)) ?
                      {(7'h42), ((8'h9e) ^~ wire99)} : ({(8'hbc)} ?
                          {reg110} : (wire99 + reg108)))));
              reg113 <= {$signed(wire103[(5'h13):(3'h7)])};
              reg114 <= forvar106[(4'hd):(3'h7)];
              reg115 <= $signed($unsigned((wire96 ? wire103 : "1Fx")));
            end
          if ((~^(-$unsigned(((~reg112) <<< $signed((8'ha8)))))))
            begin
              reg116 <= reg113[(3'h6):(2'h3)];
            end
          else
            begin
              reg116 <= ($unsigned((~&"Mcoud0IocBQuC")) < (8'ha7));
            end
          for (forvar117 = (1'h0); (forvar117 < (1'h1)); forvar117 = (forvar117 + (1'h1)))
            begin
              reg118 <= $unsigned(reg116[(1'h1):(1'h1)]);
              reg119 <= $unsigned(wire100);
            end
          for (forvar120 = (1'h0); (forvar120 < (2'h2)); forvar120 = (forvar120 + (1'h1)))
            begin
              reg121 <= wire96;
              reg122 <= (|reg108);
              reg123 <= ((^~(&wire103[(4'ha):(1'h1)])) + ((~^$signed(wire103)) || {"mwCXiTAmuL4Fl1AhldlF",
                  ((wire100 ? (7'h43) : wire103) ?
                      "mNv86QvcXkQYmgZ2k2" : (wire104 != reg114))}));
              reg124 <= "oOl";
              reg125 <= wire103;
            end
        end
      else
        begin
          reg106 <= ((reg105 <= {"xbFdg8FHCDYNssur"}) ^ (~|$signed(wire102[(4'h8):(3'h5)])));
          reg107 <= (^reg113[(3'h7):(1'h0)]);
        end
      if ((~^$unsigned({reg109[(1'h1):(1'h1)], (|"yykGPxX4IifoFt")})))
        begin
          if (reg116[(2'h2):(1'h0)])
            begin
              reg126 <= $signed({($unsigned($signed((8'h9d))) ?
                      reg107 : ((!reg118) ?
                          $unsigned(wire98) : (reg116 ? (8'hb9) : wire96)))});
              reg127 = (~reg118);
              reg128 <= "7z2v";
              reg129 <= ((~^(reg110 != $unsigned(reg114[(5'h14):(3'h6)]))) | {forvar106[(1'h0):(1'h0)],
                  reg119});
            end
          else
            begin
              reg126 <= reg109;
              reg127 <= (~^(reg123 ?
                  forvar120[(2'h3):(2'h2)] : wire97[(3'h5):(2'h2)]));
              reg128 <= "yHOy2Jh51Kmg951OOtE";
              reg129 <= ($unsigned(((reg114[(3'h7):(1'h0)] ?
                      (~^reg116) : (reg115 ? forvar117 : wire98)) ?
                  (-(-reg113)) : reg106[(3'h7):(1'h1)])) <= wire100[(4'hb):(2'h3)]);
              reg130 = (!(!$signed(reg123)));
            end
        end
      else
        begin
          if ("uq")
            begin
              reg126 <= reg125[(1'h0):(1'h0)];
            end
          else
            begin
              reg126 = (+(reg129 ?
                  (((8'hb7) < (reg123 ?
                      (8'ha2) : forvar117)) ~^ ((|wire102) >= "JngdBkDIqJPIFJKM")) : ($unsigned(((8'had) << reg105)) ?
                      "xcDq93l9OmciQcCIDW305" : $signed((forvar120 != wire104)))));
              reg127 <= {forvar106};
            end
        end
    end
  assign wire131 = {"4l"};
  assign wire132 = $signed($signed("SBTZgs0LPL8Y6TmdbH7"));
  assign wire133 = wire103[(5'h10):(4'h8)];
  assign wire134 = $unsigned({"LPvFzfzcpFaFWnhD0"});
  assign wire135 = "eUlwWYcGt6UtE";
  assign wire136 = $signed((($unsigned((+reg106)) || reg124) ?
                       ((^((8'hb1) ^ (8'h9d))) ?
                           $signed($signed((8'hbe))) : reg123) : {reg130,
                           reg123}));
  assign wire137 = $unsigned(wire99[(4'hb):(4'h9)]);
  always
    @(posedge clk) begin
      for (forvar138 = (1'h0); (forvar138 < (2'h2)); forvar138 = (forvar138 + (1'h1)))
        begin
          reg139 <= "";
          reg140 <= (($signed($signed({wire101, reg107})) ?
                  $signed({(!reg118)}) : {"lYGO9R3KXJrSbFnPy", "n2Yd"}) ?
              ($signed($unsigned(((8'hb3) ? reg119 : (8'ha8)))) ?
                  (reg121[(1'h1):(1'h1)] ?
                      (~&wire135[(3'h4):(1'h1)]) : "q1XxXl6Q") : (7'h48)) : $signed(({(-reg113)} ^ {(-reg113)})));
        end
      for (forvar141 = (1'h0); (forvar141 < (3'h4)); forvar141 = (forvar141 + (1'h1)))
        begin
          if ((8'ha5))
            begin
              reg142 <= ({($unsigned(reg129) ? "fZDBPCCrquWywaXi2" : reg113),
                      "MHwemJpbOcgPWikoJ"} ?
                  "ufmSZHart50rW" : $unsigned($signed("HIM4weno7UfPqmzM")));
              reg143 <= ($signed((reg126 ? reg142 : reg106[(2'h2):(1'h0)])) ?
                  reg112 : $signed(($unsigned((^wire131)) ?
                      (8'h9d) : reg123[(2'h3):(1'h0)])));
            end
          else
            begin
              reg142 = (reg124 ^ (+reg119));
            end
          reg144 = {(($unsigned($signed(reg122)) ^~ wire136) ?
                  ((wire96 ?
                      {reg127} : (wire136 ?
                          wire131 : (7'h46))) && ((forvar138 ~^ wire136) ?
                      $unsigned(reg125) : "o0ZMc9eyYq")) : $unsigned({reg127,
                      (reg139 * wire97)}))};
        end
    end
  always
    @(posedge clk) begin
      reg145 <= (~&"4JaUn");
      if ((reg109[(3'h4):(3'h4)] ?
          $unsigned($signed(($unsigned(wire99) ?
              reg108[(1'h0):(1'h0)] : $unsigned(wire99)))) : "hYWVrhL"))
        begin
          reg146 = (8'ha6);
          reg147 <= (8'hb5);
          for (forvar148 = (1'h0); (forvar148 < (2'h2)); forvar148 = (forvar148 + (1'h1)))
            begin
              reg149 <= $signed((-((8'hab) ~^ $signed((~reg128)))));
              reg150 <= reg125[(3'h6):(2'h2)];
              reg151 <= $signed(wire131);
            end
          for (forvar152 = (1'h0); (forvar152 < (2'h3)); forvar152 = (forvar152 + (1'h1)))
            begin
              reg153 <= $unsigned(wire97);
              reg154 <= (~|((!$unsigned({reg113, wire137})) << (|forvar138)));
              reg155 <= $unsigned($signed(reg114[(2'h3):(2'h2)]));
              reg156 = (!(~wire104[(2'h3):(1'h1)]));
              reg157 <= (|reg128);
            end
          if (reg126[(3'h7):(1'h1)])
            begin
              reg158 <= (reg156 ?
                  ($unsigned("PFza82YmMsXc8QR5GNrtN") ?
                      wire136 : reg146[(1'h1):(1'h1)]) : $unsigned($unsigned(reg112[(3'h7):(3'h5)])));
              reg159 = reg139;
              reg160 <= ({{$unsigned({(7'h43)}), {reg157}},
                      ($signed(((8'ha1) ? reg126 : (8'hac))) ?
                          "ZqSb0AD0" : "T0zcrpLn6xPPG9")} ?
                  {({$signed(reg128), reg154[(2'h3):(2'h3)]} ?
                          (7'h48) : reg147[(3'h4):(3'h4)])} : reg159[(4'hc):(4'h9)]);
              reg161 <= "pG3f";
            end
          else
            begin
              reg158 <= reg115[(3'h4):(1'h0)];
              reg159 <= (!$signed((forvar106 <= "v7P4BTeiUpa2UA1wW")));
              reg160 <= {$signed($signed({(reg143 ? wire135 : reg116)})),
                  "Via1YHwdTu"};
              reg161 <= forvar106[(4'h8):(2'h3)];
              reg162 <= $signed((7'h47));
            end
        end
      else
        begin
          for (forvar146 = (1'h0); (forvar146 < (1'h1)); forvar146 = (forvar146 + (1'h1)))
            begin
              reg147 <= (wire103[(5'h13):(2'h3)] ? {reg112} : forvar141);
            end
          if (wire99)
            begin
              reg148 = (^$unsigned({("lcTd8" && $signed(reg127)),
                  (^{reg147})}));
            end
          else
            begin
              reg148 <= (8'hbf);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar163 = (1'h0); (forvar163 < (3'h4)); forvar163 = (forvar163 + (1'h1)))
        begin
          reg164 <= wire135[(4'hc):(4'hb)];
          if ($signed(reg122[(5'h10):(5'h10)]))
            begin
              reg165 <= (("yeUFUO2l" ?
                  "BGE2HaUlCz43btBWLVk1" : reg107[(2'h3):(1'h1)]) != $unsigned((-(^~(reg115 * reg150)))));
              reg166 <= $signed($unsigned((forvar106[(4'h8):(3'h5)] ?
                  reg113[(2'h3):(2'h3)] : ((~&wire133) ?
                      $unsigned(reg113) : "VW7YO2bgxnP"))));
            end
          else
            begin
              reg165 <= "smMAovg4Fu4";
            end
        end
      reg167 = $unsigned((~|reg153));
    end
  assign wire168 = reg115;
  assign wire169 = $unsigned((reg149[(5'h11):(4'h9)] - "WvZHFHGdDn6qpIQtvZ"));
  assign wire170 = forvar106;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module609  (y, clk, wire614, wire613, wire612, wire611, wire610);
  output wire [(32'h1d7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire614;
  input wire signed [(5'h12):(1'h0)] wire613;
  input wire signed [(3'h5):(1'h0)] wire612;
  input wire [(4'hb):(1'h0)] wire611;
  input wire signed [(5'h13):(1'h0)] wire610;
  wire [(3'h5):(1'h0)] wire648;
  wire [(5'h16):(1'h0)] wire647;
  wire signed [(3'h6):(1'h0)] wire646;
  wire [(4'h8):(1'h0)] wire645;
  wire [(2'h3):(1'h0)] wire644;
  wire [(5'h17):(1'h0)] wire643;
  wire signed [(5'h17):(1'h0)] wire642;
  wire signed [(4'hd):(1'h0)] wire641;
  wire [(2'h2):(1'h0)] wire640;
  wire signed [(5'h13):(1'h0)] wire639;
  wire [(3'h7):(1'h0)] wire638;
  wire [(4'he):(1'h0)] wire637;
  reg signed [(5'h10):(1'h0)] reg636 = (1'h0);
  reg [(4'hf):(1'h0)] reg635 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar634 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg633 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg632 = (1'h0);
  reg [(5'h13):(1'h0)] reg631 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg629 = (1'h0);
  reg [(3'h4):(1'h0)] forvar622 = (1'h0);
  reg [(5'h10):(1'h0)] forvar620 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg618 = (1'h0);
  reg [(3'h4):(1'h0)] reg630 = (1'h0);
  reg [(5'h13):(1'h0)] forvar629 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg627 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg626 = (1'h0);
  reg [(5'h10):(1'h0)] reg625 = (1'h0);
  reg [(4'h8):(1'h0)] reg624 = (1'h0);
  reg [(4'he):(1'h0)] reg623 = (1'h0);
  reg [(4'h9):(1'h0)] reg622 = (1'h0);
  reg [(4'h9):(1'h0)] reg621 = (1'h0);
  reg [(4'ha):(1'h0)] reg620 = (1'h0);
  reg [(4'he):(1'h0)] reg619 = (1'h0);
  reg [(4'h8):(1'h0)] forvar618 = (1'h0);
  reg [(5'h13):(1'h0)] reg617 = (1'h0);
  wire [(5'h17):(1'h0)] wire616;
  wire [(3'h4):(1'h0)] wire615;
  assign y = {wire648,
                 wire647,
                 wire646,
                 wire645,
                 wire644,
                 wire643,
                 wire642,
                 wire641,
                 wire640,
                 wire639,
                 wire638,
                 wire637,
                 reg636,
                 reg635,
                 forvar634,
                 reg633,
                 reg632,
                 reg631,
                 reg629,
                 forvar622,
                 forvar620,
                 reg618,
                 reg630,
                 forvar629,
                 reg628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 reg619,
                 forvar618,
                 reg617,
                 wire616,
                 wire615,
                 (1'h0)};
  assign wire615 = (!wire614);
  assign wire616 = {$signed($signed(wire614[(2'h2):(1'h0)]))};
  always
    @(posedge clk) begin
      if ("6Gcv")
        begin
          reg617 <= $signed("");
          for (forvar618 = (1'h0); (forvar618 < (1'h0)); forvar618 = (forvar618 + (1'h1)))
            begin
              reg619 <= {(wire614 >= ({wire611[(2'h2):(2'h2)],
                      (reg617 ? wire610 : wire611)} * wire612[(1'h0):(1'h0)])),
                  "xEtZuPrAn"};
              reg620 <= {($unsigned((8'ha0)) ?
                      (wire612[(3'h5):(2'h2)] ?
                          ((7'h40) <<< wire611[(3'h6):(2'h2)]) : ($unsigned(wire610) > (reg617 ?
                              forvar618 : wire616))) : (wire611 * ((|forvar618) ?
                          $signed(wire612) : (~|(8'hb3)))))};
            end
          if (($signed($signed({wire615[(1'h1):(1'h1)], $signed(reg617)})) ?
              $signed($signed(("B18gqYhN9gwDKW" ?
                  wire615 : (^wire612)))) : $unsigned((~^$signed(reg619[(3'h5):(2'h2)])))))
            begin
              reg621 = wire613;
              reg622 <= $unsigned(forvar618[(1'h1):(1'h1)]);
            end
          else
            begin
              reg621 <= $signed($signed(reg617[(3'h7):(3'h5)]));
              reg622 <= (|$signed((~^reg621)));
              reg623 <= (8'hb5);
              reg624 <= ($signed("7p1KNE3NHYCD3BgDZw9xUP") < (($unsigned(reg621) && forvar618) ?
                  wire616 : reg620));
            end
          if (wire610)
            begin
              reg625 <= reg623[(1'h0):(1'h0)];
              reg626 <= ($signed(reg617) != reg625);
              reg627 <= ({reg617,
                  $unsigned($unsigned(wire614))} || "ZacvkJky5Kk1e");
              reg628 <= ("6OEwnr1wvfZbS4E" ?
                  ((+(~|$unsigned((8'hbc)))) ?
                      {(~^$unsigned(reg627))} : $unsigned(((reg623 ?
                          reg623 : reg619) >>> $signed((8'h9c))))) : $signed(wire616[(4'hb):(4'hb)]));
            end
          else
            begin
              reg625 = $signed((reg617[(2'h2):(2'h2)] >= ((-$signed(wire610)) ?
                  (&reg627) : reg619)));
              reg626 <= (~&"6N2KVC6Oxh1qJZp6");
              reg627 = wire614;
            end
          for (forvar629 = (1'h0); (forvar629 < (2'h2)); forvar629 = (forvar629 + (1'h1)))
            begin
              reg630 <= "ihFrXGfObt3Iw3KHncyq";
            end
        end
      else
        begin
          if ($signed($unsigned($signed({reg628,
              (reg623 ? (8'ha9) : (8'ha6))}))))
            begin
              reg617 <= "oGY6D7mq8lLZVfr1RGv";
              reg618 <= $signed($signed(($signed((reg626 < wire610)) ?
                  reg628 : ("L1fwUlXXpvvdED0yw9" ^ (wire612 || (8'hbb))))));
            end
          else
            begin
              reg617 <= reg624[(4'h8):(3'h6)];
              reg618 <= wire616;
              reg619 <= reg627[(4'he):(4'hc)];
            end
          for (forvar620 = (1'h0); (forvar620 < (1'h0)); forvar620 = (forvar620 + (1'h1)))
            begin
              reg621 = "Thg7aDV";
            end
          for (forvar622 = (1'h0); (forvar622 < (1'h1)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 <= $signed((~|$unsigned(forvar618)));
              reg624 <= reg626[(3'h6):(2'h2)];
            end
          if ((reg622[(3'h4):(1'h0)] ?
              ((^~$unsigned($unsigned(reg624))) ~^ {((+wire610) - (|forvar629))}) : $unsigned($unsigned($signed((wire614 ?
                  wire614 : wire615))))))
            begin
              reg625 <= (((^~wire616) ?
                  reg623[(3'h5):(2'h3)] : ($signed("FKkN2wnVC7Sz") == $signed($unsigned(reg630)))) >> "ToXkng4");
              reg626 <= $signed(wire611);
            end
          else
            begin
              reg625 <= (~|"ZnyVOCN1SqQuvM4me");
              reg626 <= "b";
              reg627 <= (forvar622[(1'h0):(1'h0)] != (&$signed((~^reg620))));
              reg628 = $signed((^~"cFGJV8nqV"));
            end
          if ({$signed({$signed(reg627[(4'h9):(2'h3)]),
                  (^reg620[(4'ha):(4'h9)])}),
              wire614[(1'h1):(1'h1)]})
            begin
              reg629 <= reg630;
              reg630 <= ((&reg619) ?
                  $unsigned((8'hba)) : ($signed($signed((~&reg621))) ?
                      reg620[(4'h8):(4'h8)] : wire613[(4'h9):(1'h1)]));
            end
          else
            begin
              reg629 <= "YS";
              reg630 <= $signed((-reg623));
              reg631 <= $signed(reg629);
              reg632 <= ((reg625 + (8'hbc)) ?
                  "uSAPQpRGH9In49D76Trrq" : $unsigned($signed($unsigned($signed(wire616)))));
              reg633 <= $signed(({wire611} ^~ {(&$signed((8'had))),
                  $signed("IdTXFBY1oL006WGJfzN")}));
            end
        end
      for (forvar634 = (1'h0); (forvar634 < (2'h2)); forvar634 = (forvar634 + (1'h1)))
        begin
          reg635 <= "i84k8gU9BVOepmJOK";
          reg636 <= {$unsigned({forvar622[(2'h3):(1'h1)],
                  ($unsigned(forvar618) >= reg627[(4'hf):(4'h8)])})};
        end
    end
  assign wire637 = forvar629;
  assign wire638 = (^$unsigned((~^((!forvar622) ?
                       (-reg619) : (reg618 > reg635)))));
  assign wire639 = {($signed(("9lffgRB" ?
                               $signed(reg631) : (reg621 == reg619))) ?
                           $signed({wire612[(2'h3):(2'h3)]}) : {wire611[(1'h1):(1'h1)],
                               reg635})};
  assign wire640 = (+(reg635[(4'h9):(3'h5)] ?
                       (wire613 ?
                           $unsigned((reg619 << reg635)) : "5BMdqt") : (-{reg622})));
  assign wire641 = ($unsigned(reg635) ?
                       $unsigned("mApoFwMto21pO") : $signed("RfeUEvZkTHBILvZHG"));
  assign wire642 = ({$signed("xMAu0Hq6wfvBtmdnW0")} ?
                       (($signed((^~reg628)) ?
                               (^~(wire641 >>> reg624)) : reg618[(4'he):(3'h4)]) ?
                           "mG" : $signed(wire639[(4'h9):(2'h3)])) : (!(($signed(reg621) <<< wire610) ?
                           ($unsigned(reg630) ?
                               reg632 : ((8'haa) ~^ (8'hba))) : {reg619,
                               "BahnkqP1xFzOYb"})));
  assign wire643 = $signed(wire610);
  assign wire644 = (reg633[(3'h5):(3'h4)] ?
                       ($unsigned($unsigned($unsigned(forvar620))) == (($signed((8'h9c)) || "BfTcIoQQv0odwSh") ?
                           (&"nfE2tcCFVMM6RRzfgrii7f") : {"S91B4wyacu7"})) : $unsigned((reg627[(4'hb):(1'h0)] | reg632[(4'hb):(1'h0)])));
  assign wire645 = wire612;
  assign wire646 = reg627;
  assign wire647 = reg622[(1'h1):(1'h0)];
  assign wire648 = wire638;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module478
#( parameter param605 = ((^((~|(+(8'ha0))) >> {((7'h41) - (8'hbb))})) ? (&((((8'had) < (8'hae)) ? {(8'ha8), (8'ha2)} : ((8'h9e) || (8'hb3))) ? ({(7'h47)} * ((8'hac) ? (7'h47) : (8'ha4))) : {((8'hb6) || (8'hb9)), ((8'hbb) ? (8'hae) : (8'h9f))})) : (({{(8'ha4), (8'h9f)}} << (^(8'hb8))) >>> (~^(~&{(8'h9c), (8'hbc)})))) )
(y, clk, wire483, wire482, wire481, wire480, wire479);
  output wire [(32'h57a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire483;
  input wire [(2'h3):(1'h0)] wire482;
  input wire [(5'h11):(1'h0)] wire481;
  input wire signed [(5'h17):(1'h0)] wire480;
  input wire [(5'h10):(1'h0)] wire479;
  wire [(4'h8):(1'h0)] wire604;
  reg signed [(4'hd):(1'h0)] reg603 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg602 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg601 = (1'h0);
  reg [(4'h8):(1'h0)] reg600 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg599 = (1'h0);
  reg [(3'h4):(1'h0)] forvar598 = (1'h0);
  reg [(3'h6):(1'h0)] reg597 = (1'h0);
  reg [(3'h6):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg595 = (1'h0);
  reg [(4'hc):(1'h0)] reg594 = (1'h0);
  reg [(3'h7):(1'h0)] reg593 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar592 = (1'h0);
  reg [(4'h9):(1'h0)] reg591 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg590 = (1'h0);
  reg signed [(4'he):(1'h0)] reg589 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg588 = (1'h0);
  reg [(5'h17):(1'h0)] reg587 = (1'h0);
  reg [(4'ha):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg585 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg584 = (1'h0);
  reg signed [(4'he):(1'h0)] reg583 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg582 = (1'h0);
  reg [(4'hc):(1'h0)] reg581 = (1'h0);
  reg [(3'h6):(1'h0)] forvar580 = (1'h0);
  reg [(3'h4):(1'h0)] forvar579 = (1'h0);
  wire [(4'h9):(1'h0)] wire578;
  reg [(5'h16):(1'h0)] reg577 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg576 = (1'h0);
  reg [(4'he):(1'h0)] reg575 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg574 = (1'h0);
  reg [(2'h2):(1'h0)] reg573 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg572 = (1'h0);
  reg [(3'h5):(1'h0)] forvar571 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar570 = (1'h0);
  reg [(2'h2):(1'h0)] reg569 = (1'h0);
  reg [(5'h17):(1'h0)] reg568 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg567 = (1'h0);
  reg [(5'h17):(1'h0)] reg566 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg565 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar563 = (1'h0);
  reg [(4'hb):(1'h0)] forvar558 = (1'h0);
  reg [(5'h13):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg562 = (1'h0);
  reg [(4'hb):(1'h0)] reg561 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg560 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg559 = (1'h0);
  reg [(2'h2):(1'h0)] reg558 = (1'h0);
  reg [(3'h6):(1'h0)] reg557 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg556 = (1'h0);
  reg [(2'h2):(1'h0)] reg555 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg554 = (1'h0);
  reg [(5'h12):(1'h0)] reg553 = (1'h0);
  reg [(4'h9):(1'h0)] forvar552 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg550 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg549 = (1'h0);
  reg [(5'h17):(1'h0)] reg548 = (1'h0);
  reg [(4'he):(1'h0)] reg547 = (1'h0);
  reg [(2'h2):(1'h0)] forvar546 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg545 = (1'h0);
  reg [(3'h6):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg543 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg542 = (1'h0);
  reg [(2'h3):(1'h0)] reg541 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg540 = (1'h0);
  reg signed [(4'he):(1'h0)] reg539 = (1'h0);
  reg [(2'h3):(1'h0)] reg534 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg538 = (1'h0);
  reg [(5'h11):(1'h0)] reg537 = (1'h0);
  reg [(4'h9):(1'h0)] reg536 = (1'h0);
  reg [(4'he):(1'h0)] reg535 = (1'h0);
  reg [(4'hc):(1'h0)] forvar534 = (1'h0);
  reg [(3'h5):(1'h0)] reg533 = (1'h0);
  reg [(3'h7):(1'h0)] reg532 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg531 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg530 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg529 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg526 = (1'h0);
  reg [(4'hd):(1'h0)] forvar525 = (1'h0);
  reg [(4'hd):(1'h0)] reg524 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg523 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar522 = (1'h0);
  reg [(2'h3):(1'h0)] reg521 = (1'h0);
  reg [(4'h8):(1'h0)] reg520 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg519 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg518 = (1'h0);
  reg signed [(4'he):(1'h0)] reg517 = (1'h0);
  reg [(5'h11):(1'h0)] forvar516 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire515;
  reg signed [(3'h6):(1'h0)] reg514 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg513 = (1'h0);
  reg [(5'h16):(1'h0)] reg512 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg511 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg510 = (1'h0);
  reg [(4'he):(1'h0)] reg509 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg508 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg507 = (1'h0);
  reg [(2'h2):(1'h0)] reg506 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg505 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg504 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire503;
  wire signed [(3'h4):(1'h0)] wire502;
  reg [(4'h8):(1'h0)] reg501 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg500 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg498 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg497 = (1'h0);
  reg [(2'h3):(1'h0)] forvar496 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire495;
  wire [(3'h4):(1'h0)] wire494;
  wire signed [(4'hb):(1'h0)] wire493;
  wire [(4'h9):(1'h0)] wire492;
  wire [(4'hb):(1'h0)] wire491;
  wire signed [(4'hf):(1'h0)] wire490;
  wire [(5'h13):(1'h0)] wire489;
  wire [(5'h16):(1'h0)] wire488;
  wire signed [(5'h12):(1'h0)] wire487;
  wire [(3'h5):(1'h0)] wire486;
  wire signed [(4'hf):(1'h0)] wire485;
  wire signed [(5'h13):(1'h0)] wire484;
  assign y = {wire604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 forvar598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 forvar592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 forvar580,
                 forvar579,
                 wire578,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 forvar571,
                 forvar570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 reg564,
                 forvar563,
                 forvar558,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 forvar552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 forvar546,
                 reg545,
                 reg544,
                 reg543,
                 reg542,
                 reg541,
                 reg540,
                 reg539,
                 reg534,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 forvar534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 forvar525,
                 reg524,
                 reg523,
                 forvar522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 forvar516,
                 wire515,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 wire503,
                 wire502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 forvar496,
                 wire495,
                 wire494,
                 wire493,
                 wire492,
                 wire491,
                 wire490,
                 wire489,
                 wire488,
                 wire487,
                 wire486,
                 wire485,
                 wire484,
                 (1'h0)};
  assign wire484 = "aAG";
  assign wire485 = (wire482[(2'h2):(2'h2)] ?
                       (+"03QioxJ2G6bcNBLSWpO4A") : wire481[(2'h3):(1'h1)]);
  assign wire486 = "7ufuSMofZep2tSsHn6UnJy";
  assign wire487 = $unsigned((-wire483[(3'h7):(3'h4)]));
  assign wire488 = $unsigned((({wire486,
                       wire481[(3'h5):(2'h3)]} | wire480[(5'h13):(4'h9)]) - "YuDgQH203kCsx91AZ7"));
  assign wire489 = $signed(wire482);
  assign wire490 = (!wire482[(2'h3):(2'h3)]);
  assign wire491 = wire490;
  assign wire492 = wire484[(4'h8):(3'h4)];
  assign wire493 = ((!$signed("tGWETJrS9qsFI")) ?
                       $unsigned("ZWd2V") : $unsigned(($signed(wire487) ?
                           $unsigned(wire480) : (|$unsigned(wire488)))));
  assign wire494 = ($unsigned($signed(wire491[(2'h3):(1'h1)])) >= ($signed($unsigned((wire493 ?
                       wire490 : (8'haf)))) ^ $unsigned("fbdk")));
  assign wire495 = ("Jrp68b" | ($unsigned(((wire487 ? wire480 : wire490) ?
                           wire479[(5'h10):(4'hd)] : (8'ha7))) ?
                       (|wire482) : (!"kXqYZcl")));
  always
    @(posedge clk) begin
      for (forvar496 = (1'h0); (forvar496 < (3'h4)); forvar496 = (forvar496 + (1'h1)))
        begin
          if ("uhSO6J5nfJKi1TIcMx")
            begin
              reg497 <= ((-(wire483 ?
                  wire493[(2'h2):(2'h2)] : {wire489[(5'h11):(3'h7)],
                      {(7'h44), wire494}})) * $signed((!$unsigned(wire488))));
              reg498 <= wire491[(2'h2):(1'h0)];
              reg499 <= (wire486[(2'h2):(2'h2)] == reg498);
              reg500 <= (^$signed($signed(wire485)));
            end
          else
            begin
              reg497 <= $unsigned(((^($signed(wire487) > (wire480 ?
                  wire491 : (8'had)))) << $unsigned(($signed((8'hab)) ?
                  $unsigned(wire480) : wire485))));
              reg498 <= wire494[(1'h1):(1'h0)];
              reg499 <= $signed("2");
            end
        end
      reg501 <= ((7'h48) ? (^~wire485) : ("KNGcQyHSb8r00B" < wire485));
    end
  assign wire502 = ((wire479 << wire479[(4'hb):(4'ha)]) == forvar496);
  assign wire503 = ({wire482, "g2Nv"} ?
                       $signed("kr2CVYtGmZLlfu9vkJh") : ((wire486 ?
                               (8'hbc) : wire481) ?
                           ((+(-wire492)) ^~ $unsigned(wire487)) : "TTNAmLLiiaS8Ty8MKl"));
  always
    @(posedge clk) begin
      reg504 <= (wire495[(1'h1):(1'h0)] ?
          {$unsigned($signed($signed((8'hb3)))),
              $signed({{(7'h44), (8'hb9)}})} : reg499[(1'h1):(1'h1)]);
      reg505 <= ("HdBZgvBIY" << $unsigned({wire495}));
      if (($unsigned($unsigned(((wire482 & wire486) + $signed((8'hac))))) ?
          $signed($signed("3TKgu5Hc5sO1")) : $signed((!$unsigned((wire491 ^ wire493))))))
        begin
          if ({(!forvar496[(1'h0):(1'h0)])})
            begin
              reg506 <= (~&reg504);
              reg507 <= (wire479 ?
                  "4DoyctTHNKDnxC0Ltp4rfY" : ({(&wire489)} >> $unsigned("sN")));
            end
          else
            begin
              reg506 <= "ukOGN7hqRqSxFCa";
              reg507 = "U5tdwlwD4qyLeJCmlLwkw";
              reg508 <= wire495[(1'h0):(1'h0)];
              reg509 = wire491[(3'h5):(3'h4)];
              reg510 <= reg499;
            end
        end
      else
        begin
          if (reg497[(1'h1):(1'h0)])
            begin
              reg506 <= $unsigned(({$unsigned(forvar496[(1'h0):(1'h0)])} ?
                  wire503 : $unsigned(wire490[(2'h2):(2'h2)])));
              reg507 <= (~|$unsigned($signed($unsigned(wire491[(3'h5):(2'h3)]))));
              reg508 <= reg500;
            end
          else
            begin
              reg506 <= $signed((-(~^"2Z2gvAMLeMkwwgY")));
              reg507 <= reg507[(2'h3):(1'h0)];
              reg508 <= $signed({((^"oPFqeEAmCTi2A6GeNPotRl") ^~ {(wire493 < wire481)})});
            end
          reg509 <= (7'h43);
          reg510 = $unsigned((-$signed(wire502)));
          if ((^~(-(+(+(reg510 ? (8'hbe) : reg507))))))
            begin
              reg511 = (8'hb2);
            end
          else
            begin
              reg511 <= (wire481[(4'hc):(4'hc)] ? {"XOlhhYq5Hg"} : wire488);
              reg512 = ((+$unsigned(reg499[(4'hd):(4'ha)])) || ("tJe4OaU6KPwe0QPRZmV" ?
                  (({wire480} <= (reg509 ? wire484 : wire480)) ?
                      (~(~&reg504)) : wire482) : (wire491 ?
                      $signed((!(8'hb9))) : ($unsigned(wire481) ?
                          (^~(7'h43)) : (wire484 ? reg508 : reg498)))));
              reg513 <= $signed("iofuM");
            end
        end
      reg514 = wire485;
    end
  assign wire515 = (&($signed($unsigned((^~reg507))) && wire484[(4'hc):(4'hc)]));
  always
    @(posedge clk) begin
      for (forvar516 = (1'h0); (forvar516 < (2'h3)); forvar516 = (forvar516 + (1'h1)))
        begin
          if (((|"72") ?
              (&(wire485[(4'hf):(1'h1)] ?
                  ((|wire482) ?
                      wire485[(4'h8):(3'h4)] : $signed(reg511)) : wire492[(2'h2):(1'h1)])) : {wire515[(4'hd):(3'h5)],
                  (7'h45)}))
            begin
              reg517 <= "ESQc1oUsJ";
              reg518 <= wire489[(4'hf):(3'h7)];
              reg519 <= (-({$signed($signed(reg497))} - (8'ha1)));
              reg520 <= (!$unsigned((+$signed(wire485[(4'hd):(4'h9)]))));
              reg521 <= (reg504 ?
                  $unsigned({"fsh"}) : (^(~&reg497[(3'h6):(3'h6)])));
            end
          else
            begin
              reg517 <= $unsigned((wire494[(2'h3):(2'h2)] * $signed((~^"GL5P"))));
              reg518 <= reg505;
              reg519 <= ({("1kB" ^ ("9MgSRFQM1MQWQRBKIAo05M" >> wire493[(1'h0):(1'h0)]))} >>> "8g4E7rxNIu0C8sfBgYY8Z");
              reg520 <= reg518[(4'h9):(3'h5)];
              reg521 <= $unsigned(($unsigned("3") ?
                  "7LFN4ua0MB986qIVtb" : $unsigned(wire481)));
            end
          for (forvar522 = (1'h0); (forvar522 < (3'h4)); forvar522 = (forvar522 + (1'h1)))
            begin
              reg523 = wire491[(4'hb):(3'h6)];
              reg524 = $signed(($unsigned((+$unsigned(wire488))) ?
                  (!($unsigned(reg517) << $signed(reg512))) : (|$signed(wire488))));
            end
          for (forvar525 = (1'h0); (forvar525 < (3'h4)); forvar525 = (forvar525 + (1'h1)))
            begin
              reg526 <= ((~&(^~(~|(|wire484)))) ?
                  forvar496[(1'h0):(1'h0)] : ((wire495[(2'h2):(1'h0)] ?
                      (~|(~&(8'hb8))) : reg506[(1'h1):(1'h0)]) || wire488));
              reg527 <= "T2UH9UaTf3Zx";
              reg528 <= (8'hb7);
              reg529 <= $signed(reg513);
            end
          if ((+reg524))
            begin
              reg530 = ((((wire487[(3'h7):(3'h7)] + ((8'haa) ?
                          (8'hba) : reg497)) ?
                      $unsigned(reg514[(2'h2):(1'h0)]) : "p3C7vOIB0FHT4iAHcteQb") + reg510[(1'h0):(1'h0)]) ?
                  {(((forvar522 ?
                          reg507 : reg523) | (reg521 >> wire481)) ~^ reg521[(2'h3):(2'h2)]),
                      {((~|reg520) ?
                              (wire488 ? forvar522 : reg511) : "GEpL36BaSrWkY"),
                          $signed(((8'ha1) ?
                              reg505 : reg514))}} : (((~&$unsigned(reg509)) ?
                          ({wire487} == reg506[(1'h1):(1'h1)]) : $unsigned((|(8'h9c)))) ?
                      $signed(((forvar522 <= reg514) ?
                          "bO8pQKanbJ" : "SeBN7IrViUp")) : reg524));
              reg531 <= "7P9be";
            end
          else
            begin
              reg530 <= {$unsigned((7'h43))};
              reg531 = {(!(reg498 ^ (~$unsigned((8'hae)))))};
              reg532 <= $unsigned((8'haf));
            end
        end
      reg533 <= "9mNAm7Ii0OZqlg2XKwL";
      if (wire479[(2'h2):(2'h2)])
        begin
          for (forvar534 = (1'h0); (forvar534 < (2'h2)); forvar534 = (forvar534 + (1'h1)))
            begin
              reg535 <= wire486;
              reg536 = reg512[(5'h10):(3'h4)];
              reg537 <= (($unsigned((8'hba)) ^~ "VsOq") && {("KOpuZERXRRRG7C" ?
                      "SwDgZED" : {reg517, (reg513 <<< (8'ha1))})});
              reg538 <= (($unsigned($unsigned($unsigned(wire491))) >> forvar496[(1'h1):(1'h1)]) ?
                  (wire494 ?
                      (8'hb5) : forvar496[(2'h3):(2'h2)]) : {(|forvar525)});
            end
        end
      else
        begin
          reg534 <= (+(wire490[(4'h8):(3'h7)] != (reg526[(2'h3):(2'h2)] ?
              ((~wire515) ^ wire493) : "LsdN7thRbe7oAseGZwF6")));
          if (({(!"kmAP7s2O5PGR")} ?
              $unsigned((reg509[(3'h6):(3'h6)] ?
                  forvar534 : (^(wire481 && wire485)))) : (~|"Z00uhtAistdua")))
            begin
              reg535 <= $unsigned(reg521[(2'h2):(2'h2)]);
              reg536 <= (~|(((^(-reg526)) ?
                  ($signed(reg498) <<< (wire486 ?
                      reg529 : wire485)) : (~&"G11T4k1GEDa09IvxGCXpA")) <= (($unsigned(wire493) ?
                      (+(8'hb4)) : {reg533, reg531}) ?
                  ((~|(7'h47)) ?
                      reg526[(2'h3):(2'h3)] : (&(7'h47))) : $signed(reg511[(1'h1):(1'h1)]))));
              reg537 <= $signed((($signed("H0NVhHGHZkV3gEwU") + wire493[(4'h8):(1'h0)]) ^ $signed((~&(wire494 != (8'hb7))))));
              reg538 <= $unsigned(wire493[(4'ha):(3'h4)]);
              reg539 <= "ZrXAf95imqE8m4QXx";
            end
          else
            begin
              reg535 <= {$signed((|{((8'ha1) - forvar516),
                      $unsigned((8'hac))}))};
            end
          reg540 <= "3r54U9eMFw7ztUgmQ";
          reg541 = $signed($signed(reg528[(3'h4):(1'h0)]));
          if ((({$signed((~|wire488)),
              $signed((reg534 + reg527))} >>> forvar516[(4'he):(4'hd)]) | ((~^$unsigned($unsigned(reg500))) != (((wire489 ?
                      (8'hbf) : reg529) ?
                  reg535 : (wire481 < wire492)) ?
              (8'haf) : wire480))))
            begin
              reg542 <= wire492[(1'h1):(1'h0)];
              reg543 <= ((reg541[(2'h3):(1'h1)] ?
                      ((((8'haa) ? wire492 : wire484) == "5ZObv1RHXUeW0JYAV") ?
                          $unsigned($signed(reg504)) : (wire494 ?
                              {reg530,
                                  reg499} : $signed(reg506))) : ($unsigned((reg533 ?
                          reg506 : reg519)) >>> "hz5T1NOghQ")) ?
                  reg511 : (^($unsigned($signed(reg506)) ?
                      wire485 : $signed(reg514))));
              reg544 = (wire480[(2'h3):(2'h2)] ?
                  {$unsigned(reg506),
                      "dJrlE4kwDVgUpScfr"} : (~($unsigned({(8'hbd), reg531}) ?
                      $unsigned({wire491, wire493}) : wire502)));
              reg545 <= ("vDn2q" & $signed((~(|{wire515, reg506}))));
            end
          else
            begin
              reg542 <= $unsigned(reg532);
              reg543 = wire482;
              reg544 <= {$signed($unsigned((|forvar496[(1'h1):(1'h0)]))),
                  (7'h43)};
            end
        end
      for (forvar546 = (1'h0); (forvar546 < (3'h4)); forvar546 = (forvar546 + (1'h1)))
        begin
          if ($unsigned(((reg509[(3'h6):(1'h0)] ?
              $unsigned(reg498) : $unsigned(((8'h9d) - reg531))) == {(reg541 ?
                  (wire484 ? reg527 : wire495) : (wire492 * wire492))})))
            begin
              reg547 <= (reg504[(4'ha):(4'h8)] ?
                  (reg540[(3'h6):(1'h0)] ?
                      (((^reg499) > (^~reg524)) ?
                          $signed((reg504 ?
                              wire484 : forvar546)) : "Url0Mp6O1cUNw29") : {reg524[(4'hd):(3'h5)],
                          (((8'hb5) & wire483) ?
                              (wire492 || reg498) : (wire486 ?
                                  reg507 : reg537))}) : $unsigned({$unsigned(wire487[(1'h1):(1'h0)]),
                      $unsigned((reg524 ? wire483 : reg513))}));
              reg548 <= reg510[(3'h6):(3'h4)];
              reg549 <= reg529;
              reg550 <= $signed(reg548[(1'h0):(1'h0)]);
            end
          else
            begin
              reg547 = (~|reg510[(2'h3):(2'h2)]);
              reg548 <= (wire494 != wire490);
              reg549 <= "MPlsG9ZMfdxu3GEZDw6q";
              reg550 <= reg499;
              reg551 = forvar516[(4'hb):(4'hb)];
            end
          for (forvar552 = (1'h0); (forvar552 < (3'h4)); forvar552 = (forvar552 + (1'h1)))
            begin
              reg553 <= $unsigned((^reg505));
              reg554 <= reg548[(4'hf):(4'hd)];
              reg555 <= (wire484[(3'h5):(2'h3)] ?
                  {(-reg527[(5'h11):(1'h1)])} : $unsigned(reg512[(2'h3):(2'h2)]));
              reg556 <= ({$signed(wire486)} ^ ($signed(reg519[(3'h4):(2'h2)]) ?
                  (-((wire483 >>> wire490) ?
                      (+reg555) : reg523)) : "QL2NtaQSasHYSr"));
              reg557 = ($unsigned($unsigned(((reg521 || reg535) ?
                      wire495[(3'h4):(3'h4)] : wire489))) ?
                  $unsigned(reg542[(2'h2):(1'h0)]) : reg555);
            end
        end
      if ((^(~|reg506)))
        begin
          reg558 <= (wire493 | $unsigned($signed(reg557)));
          if ((~(|reg556)))
            begin
              reg559 <= $signed($signed($signed(($signed(wire482) ?
                  $unsigned(reg540) : forvar516))));
              reg560 <= (reg553 ?
                  $signed($unsigned($signed((!reg534)))) : $signed({wire491[(3'h6):(3'h6)],
                      $signed($signed(reg534))}));
              reg561 <= forvar516[(2'h2):(2'h2)];
              reg562 <= reg560;
              reg563 <= (wire485 ? (8'haf) : (~^"YnRZ"));
            end
          else
            begin
              reg559 <= (wire489[(3'h6):(2'h2)] ?
                  (&(~&$unsigned((reg513 >> forvar516)))) : (reg557[(3'h6):(3'h4)] >= reg560[(5'h14):(4'h9)]));
              reg560 <= ($signed($unsigned($signed((reg560 * reg538)))) ?
                  $unsigned(wire494[(2'h3):(1'h1)]) : (~^(~$unsigned("dyNJpF8m3a7F"))));
              reg561 = "ZyzScYO";
              reg562 <= $signed((!$signed($unsigned($signed(reg514)))));
            end
        end
      else
        begin
          for (forvar558 = (1'h0); (forvar558 < (1'h0)); forvar558 = (forvar558 + (1'h1)))
            begin
              reg559 <= ("" ?
                  ((!($unsigned(reg532) ?
                      "5HX2JqERzuJmOg9" : $unsigned(reg554))) < "SXSCdrMwVVLpPhbQxiEO") : ((&$signed($unsigned((8'ha7)))) + $signed(reg528[(2'h3):(1'h1)])));
              reg560 <= $signed((8'hbb));
              reg561 <= $unsigned("d9Wh7filTlD");
            end
          if ({$unsigned($unsigned($signed(reg537))), reg497})
            begin
              reg562 = "YHVKS5ZwBx9ktqDI";
            end
          else
            begin
              reg562 <= $unsigned(($unsigned($signed(wire492)) ^ "kYrAbsZJzWkwQw"));
            end
          for (forvar563 = (1'h0); (forvar563 < (3'h4)); forvar563 = (forvar563 + (1'h1)))
            begin
              reg564 <= $signed({$signed(((|reg511) ^~ reg497))});
              reg565 <= wire503[(4'h8):(3'h7)];
              reg566 <= (reg504[(4'h9):(1'h0)] <= (^(&((reg512 ?
                      wire479 : reg547) ?
                  $signed(wire488) : (reg560 * reg563)))));
              reg567 <= ($signed($signed(({reg538} ?
                      reg555[(2'h2):(2'h2)] : (reg509 > reg550)))) ?
                  reg520[(3'h4):(2'h3)] : $unsigned("QDZGS0"));
            end
          reg568 <= ($unsigned(({reg500[(1'h1):(1'h0)], $signed(reg559)} ?
                  $signed("lSu6Vub0qS2GlU") : forvar534[(1'h1):(1'h1)])) ?
              reg557[(2'h2):(2'h2)] : "tOn34aF9UmtRsXQsHrB");
        end
    end
  always
    @(posedge clk) begin
      reg569 = $signed($unsigned("lLbvxab7CfNsURc"));
      for (forvar570 = (1'h0); (forvar570 < (1'h1)); forvar570 = (forvar570 + (1'h1)))
        begin
          for (forvar571 = (1'h0); (forvar571 < (2'h2)); forvar571 = (forvar571 + (1'h1)))
            begin
              reg572 <= reg544;
              reg573 <= ({$signed($signed({reg518, reg542}))} ?
                  (~|reg540[(4'hd):(3'h6)]) : (reg558 == {("Gt" <<< "Tq0"),
                      {(~^reg572), $unsigned(reg509)}}));
              reg574 <= reg539[(1'h0):(1'h0)];
            end
          reg575 <= $unsigned(reg519[(1'h1):(1'h0)]);
          reg576 <= {$unsigned($signed(reg548[(4'he):(3'h5)])),
              {$unsigned((7'h45))}};
        end
      reg577 <= $unsigned(wire503[(2'h2):(1'h0)]);
    end
  assign wire578 = (&"FFyoG9nihDsEPlyN");
  always
    @(posedge clk) begin
      for (forvar579 = (1'h0); (forvar579 < (1'h0)); forvar579 = (forvar579 + (1'h1)))
        begin
          for (forvar580 = (1'h0); (forvar580 < (3'h4)); forvar580 = (forvar580 + (1'h1)))
            begin
              reg581 = ((|reg530) & $unsigned(($unsigned({reg523,
                  reg532}) && reg563)));
              reg582 = ((wire482 ?
                  $unsigned((!$unsigned(wire482))) : wire480) | wire494[(1'h0):(1'h0)]);
              reg583 = (8'h9f);
            end
          if ((+(~|"KQNdkHmb")))
            begin
              reg584 <= $signed((reg551[(4'hd):(4'hb)] >= ((~|"RtyLk5IrK") * $unsigned((reg533 > reg577)))));
            end
          else
            begin
              reg584 <= (-reg547);
              reg585 <= (~|((^~"wZBaiRxre") ?
                  (reg566 ?
                      {(~&(8'ha5))} : (~^(reg527 ^~ forvar579))) : (("RNMNBY" ?
                      "iyGlUOwv0NXZ82Wc2tv" : (reg541 ?
                          (8'had) : reg550)) * ((reg562 ? reg558 : reg553) ?
                      (reg565 - reg527) : reg561))));
              reg586 <= $unsigned(((^~wire486[(3'h5):(1'h1)]) + wire490));
            end
          if (reg530)
            begin
              reg587 <= (-reg520);
              reg588 <= "tunQPxo";
            end
          else
            begin
              reg587 <= "";
              reg588 <= ("TpO0p2CfO" & (~^($unsigned((+reg507)) == "U1OyDUtI0otlM2JAlNmcC")));
              reg589 <= $signed($signed((~&reg517[(1'h1):(1'h0)])));
              reg590 <= "gqAB";
            end
          reg591 <= {($signed(($unsigned(reg529) ?
                      $unsigned(reg499) : $signed((8'hb1)))) ?
                  reg504 : $unsigned($unsigned("SvO4qfzHfxiMBUBUP")))};
        end
      for (forvar592 = (1'h0); (forvar592 < (3'h4)); forvar592 = (forvar592 + (1'h1)))
        begin
          if (forvar525)
            begin
              reg593 <= {{{{$unsigned(reg573)},
                          ((reg588 << reg507) ~^ (reg573 ?
                              (8'hb7) : forvar496))}},
                  ((!$signed(reg500)) ?
                      (~^$signed((wire479 || reg568))) : {({reg531, reg497} ?
                              {reg559, forvar546} : $unsigned(reg527)),
                          $signed((forvar534 < reg543))})};
              reg594 <= $signed($unsigned({((~^forvar592) ?
                      (~&forvar571) : (reg508 << reg583)),
                  forvar534}));
              reg595 <= ("wVJD2kApAkfDtWv" ?
                  reg508[(3'h7):(3'h4)] : "LZUM2VFy0lG");
              reg596 <= ((^~($unsigned("ni7M3NBo6") ?
                      $unsigned("63JJZ") : ({reg531} ?
                          reg587 : $signed(forvar579)))) ?
                  "QCWbM7" : ($signed((((8'hb9) & (8'hb0)) ~^ "7X4eCpw")) > (^$signed((reg523 ~^ reg551)))));
              reg597 = $unsigned("0I0Y7EJZqPKACnzhhVMEx");
            end
          else
            begin
              reg593 <= "hCbZJggG22m";
              reg594 <= "sesDyAqIu4O9W5ZE69ZncQ";
              reg595 <= ((8'hb1) ?
                  $signed({($signed(reg554) ? reg593 : reg582)}) : ("NU5mX" ?
                      "zu2St0B3bnYp2yDa1b" : ($signed($unsigned(reg527)) ?
                          forvar496[(2'h2):(1'h1)] : wire494[(2'h2):(2'h2)])));
            end
          for (forvar598 = (1'h0); (forvar598 < (2'h2)); forvar598 = (forvar598 + (1'h1)))
            begin
              reg599 <= ("lCovUygWAwrJ2RccxZ" ?
                  $signed("92GTuOMY917qA3cu4I") : {{$unsigned($unsigned(reg529))},
                      $signed(reg594)});
              reg600 <= $signed({($signed($unsigned(reg560)) ?
                      $signed((forvar579 < reg550)) : (wire491[(4'hb):(4'hb)] && $signed(reg595))),
                  (wire578 != (~|((8'h9e) ? reg521 : reg498)))});
              reg601 <= (~&$signed((+$signed($signed(forvar570)))));
              reg602 <= $unsigned($signed("gB1LhCFh"));
            end
          reg603 <= {("vFFnFayzighIc" ?
                  reg509 : (reg563[(5'h10):(4'he)] ?
                      wire486[(2'h3):(2'h2)] : "T0eoxFVHKP"))};
        end
    end
  assign wire604 = $unsigned((("xz4xVAb33FwtirW91Jnq6z" <= ($unsigned(wire490) * {wire503})) ?
                       $signed("ufcK5JV2iMALQm") : "K"));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module374
#( parameter param473 = {({(^~((8'hb6) ? (8'hb8) : (8'ha1)))} ? {(&((8'hb8) ? (8'hbb) : (8'had))), (!(~&(8'ha1)))} : {(&((8'haf) ? (8'ha5) : (8'hbf)))})}
, parameter param474 = {(((7'h48) ? (param473 ? (param473 ? (7'h46) : param473) : (param473 ? param473 : (8'hb8))) : (~((7'h42) - param473))) ? {param473} : (({param473, (7'h42)} ? (param473 ? param473 : (8'h9e)) : param473) ? {((7'h43) > (8'h9d))} : (&(param473 ? param473 : param473)))), param473} )
(y, clk, wire379, wire378, wire377, wire376, wire375);
  output wire [(32'h4be):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire379;
  input wire signed [(5'h16):(1'h0)] wire378;
  input wire signed [(2'h3):(1'h0)] wire377;
  input wire [(4'hc):(1'h0)] wire376;
  input wire [(5'h11):(1'h0)] wire375;
  wire [(5'h14):(1'h0)] wire472;
  reg [(4'ha):(1'h0)] reg471 = (1'h0);
  reg [(2'h2):(1'h0)] reg470 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar469 = (1'h0);
  reg signed [(4'he):(1'h0)] reg468 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire467;
  wire [(3'h6):(1'h0)] wire466;
  wire signed [(3'h4):(1'h0)] wire465;
  wire [(5'h15):(1'h0)] wire464;
  wire signed [(5'h13):(1'h0)] wire463;
  wire [(5'h11):(1'h0)] wire462;
  reg signed [(5'h11):(1'h0)] reg461 = (1'h0);
  reg [(4'hd):(1'h0)] reg460 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg459 = (1'h0);
  reg [(3'h5):(1'h0)] reg458 = (1'h0);
  reg signed [(4'he):(1'h0)] reg457 = (1'h0);
  reg [(2'h3):(1'h0)] reg456 = (1'h0);
  reg [(4'he):(1'h0)] reg455 = (1'h0);
  reg [(5'h17):(1'h0)] reg454 = (1'h0);
  reg [(3'h5):(1'h0)] reg453 = (1'h0);
  reg [(4'h8):(1'h0)] forvar452 = (1'h0);
  reg [(4'ha):(1'h0)] reg452 = (1'h0);
  reg [(3'h4):(1'h0)] reg451 = (1'h0);
  reg [(5'h11):(1'h0)] reg450 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg448 = (1'h0);
  reg [(3'h4):(1'h0)] reg447 = (1'h0);
  reg [(5'h16):(1'h0)] reg446 = (1'h0);
  reg [(4'he):(1'h0)] forvar445 = (1'h0);
  reg [(4'h9):(1'h0)] reg444 = (1'h0);
  reg [(5'h13):(1'h0)] reg443 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg442 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg441 = (1'h0);
  reg [(3'h4):(1'h0)] forvar440 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg439 = (1'h0);
  reg [(5'h14):(1'h0)] reg438 = (1'h0);
  reg [(5'h11):(1'h0)] forvar437 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg436 = (1'h0);
  reg [(2'h2):(1'h0)] reg435 = (1'h0);
  reg [(5'h12):(1'h0)] reg434 = (1'h0);
  reg [(4'he):(1'h0)] reg433 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar432 = (1'h0);
  reg [(4'h9):(1'h0)] reg431 = (1'h0);
  reg [(3'h4):(1'h0)] reg430 = (1'h0);
  reg [(3'h5):(1'h0)] reg429 = (1'h0);
  reg [(2'h2):(1'h0)] reg428 = (1'h0);
  reg [(4'h8):(1'h0)] reg427 = (1'h0);
  reg [(2'h2):(1'h0)] forvar426 = (1'h0);
  reg [(4'h8):(1'h0)] reg425 = (1'h0);
  reg [(2'h3):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg423 = (1'h0);
  reg [(5'h14):(1'h0)] forvar422 = (1'h0);
  reg signed [(4'he):(1'h0)] reg421 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg420 = (1'h0);
  reg [(5'h14):(1'h0)] reg419 = (1'h0);
  reg [(4'hd):(1'h0)] reg418 = (1'h0);
  reg [(5'h16):(1'h0)] reg417 = (1'h0);
  reg [(5'h10):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar415 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar414 = (1'h0);
  reg signed [(4'he):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg412 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar411 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg410 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg409 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg408 = (1'h0);
  reg [(4'h8):(1'h0)] reg407 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg405 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar404 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg403 = (1'h0);
  reg [(4'hc):(1'h0)] forvar393 = (1'h0);
  reg [(4'h9):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg401 = (1'h0);
  reg [(3'h6):(1'h0)] reg400 = (1'h0);
  reg [(4'hd):(1'h0)] forvar399 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg397 = (1'h0);
  reg [(5'h15):(1'h0)] reg396 = (1'h0);
  reg [(4'hf):(1'h0)] reg395 = (1'h0);
  reg [(4'hf):(1'h0)] reg394 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg393 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg383 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar382 = (1'h0);
  reg [(5'h16):(1'h0)] reg392 = (1'h0);
  reg [(5'h10):(1'h0)] reg391 = (1'h0);
  reg [(5'h11):(1'h0)] forvar390 = (1'h0);
  reg [(3'h4):(1'h0)] reg389 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg388 = (1'h0);
  reg [(5'h12):(1'h0)] reg387 = (1'h0);
  reg signed [(4'he):(1'h0)] reg386 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg385 = (1'h0);
  reg [(4'hd):(1'h0)] reg384 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar383 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg382 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire381;
  wire [(4'hd):(1'h0)] wire380;
  assign y = {wire472,
                 reg471,
                 reg470,
                 forvar469,
                 reg468,
                 wire467,
                 wire466,
                 wire465,
                 wire464,
                 wire463,
                 wire462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 forvar452,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg447,
                 reg446,
                 forvar445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 forvar440,
                 reg439,
                 reg438,
                 forvar437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 forvar432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 forvar426,
                 reg425,
                 reg424,
                 reg423,
                 forvar422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 forvar415,
                 forvar414,
                 reg413,
                 reg412,
                 forvar411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 forvar404,
                 reg403,
                 forvar393,
                 reg402,
                 reg401,
                 reg400,
                 forvar399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg383,
                 forvar382,
                 reg392,
                 reg391,
                 forvar390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 forvar383,
                 reg382,
                 wire381,
                 wire380,
                 (1'h0)};
  assign wire380 = $signed(("KxH3D4XMqgfBILCllzUIZp" ^~ $unsigned((-$signed(wire376)))));
  assign wire381 = $unsigned(wire380[(3'h7):(3'h6)]);
  always
    @(posedge clk) begin
      if ("nJvsh2mOr")
        begin
          reg382 <= (!($signed((wire376[(1'h0):(1'h0)] ?
              wire375[(2'h3):(1'h1)] : (wire375 - wire376))) < $signed(((&wire381) & (wire380 * wire379)))));
          for (forvar383 = (1'h0); (forvar383 < (1'h1)); forvar383 = (forvar383 + (1'h1)))
            begin
              reg384 <= $signed($signed("uBF5ilmiZZA9afMw7RA"));
            end
          if (($unsigned(($signed((+reg382)) * (reg384 ^~ "u"))) ?
              forvar383 : (wire380 ?
                  {$signed((wire375 <= reg382)),
                      ((&reg384) ?
                          {(8'hb2),
                              wire377} : wire381[(5'h15):(5'h10)])} : (wire380[(2'h3):(2'h3)] >= (+$unsigned(wire379))))))
            begin
              reg385 <= $unsigned((wire376[(3'h5):(2'h2)] ?
                  reg382[(3'h4):(1'h0)] : (("RR5FQL" ? $signed((8'hb8)) : "c") ?
                      $unsigned(reg382[(5'h11):(4'hd)]) : $unsigned((+forvar383)))));
              reg386 <= $unsigned($signed($unsigned(forvar383[(3'h6):(3'h5)])));
              reg387 <= "vUz3NvPP0QVZdI7";
              reg388 <= {(("wNod" <= wire376) & {"cXXCiORV"}),
                  wire375[(3'h6):(1'h0)]};
              reg389 <= ($signed($unsigned($signed($signed(wire378)))) ?
                  (~"dtYJ") : wire377);
            end
          else
            begin
              reg385 = (-"fy");
              reg386 = "HG4rIHAxZTgPU";
              reg387 <= (wire377 ?
                  reg387[(4'hd):(3'h4)] : ($signed(reg384) ?
                      {(wire379 ? wire375 : (~^wire380))} : wire381));
              reg388 <= ({(~&$signed(((8'hba) + wire380))),
                      {(~(+wire380)),
                          ("B0ZmgIxg5sUEY1" ?
                              forvar383 : $signed(forvar383))}} ?
                  ($unsigned(($signed(reg385) <<< "9uSrJskzhFTtB8PWf")) >>> {($signed(reg389) && $unsigned(wire381))}) : "zlxMlR4hCUdE4");
            end
          for (forvar390 = (1'h0); (forvar390 < (1'h1)); forvar390 = (forvar390 + (1'h1)))
            begin
              reg391 <= $unsigned(("nBYiBa2M0eCNIk0" ?
                  (reg385 ?
                      wire380 : $unsigned("JEJEPFxEo8f5A4")) : (~^($signed((7'h42)) >= $signed((8'ha4))))));
              reg392 <= $signed(wire381[(4'hb):(4'h8)]);
            end
        end
      else
        begin
          for (forvar382 = (1'h0); (forvar382 < (2'h2)); forvar382 = (forvar382 + (1'h1)))
            begin
              reg383 <= wire381;
            end
          if ($unsigned(({$unsigned("bp2BJ1WRQdVfxFK4shrL"),
              (+(wire381 * reg384))} ^~ (((+forvar383) || (reg392 || forvar382)) < ($unsigned(wire375) ?
              (forvar382 < wire379) : $unsigned(wire379))))))
            begin
              reg384 <= reg392;
              reg385 <= $unsigned((^(~(8'hac))));
              reg386 = reg389[(3'h4):(2'h2)];
            end
          else
            begin
              reg384 <= ((|"Hgd24NGv9YJbZniPoAcSw") ?
                  reg384 : {("sCkZ2eD" <= ((wire381 ?
                          wire381 : reg392) + (+forvar382))),
                      (($unsigned(forvar382) ?
                          (reg384 ? wire378 : wire376) : (wire380 ?
                              reg385 : reg385)) <= reg386)});
              reg385 <= $unsigned((+(($unsigned((7'h47)) ^ {wire379, (7'h40)}) ?
                  (!(~^wire381)) : reg392)));
              reg386 <= (reg387 + wire381);
              reg387 <= ("gBZq8C7J5" ^~ "xU1Qr53i4");
              reg388 <= "FTp";
            end
          reg389 = "0CwuXfD53V9Ma8DBZX2ye";
        end
      if ((wire377 ?
          ($unsigned(((~|reg388) >> "7yg1AZ5XzriyY6mZk")) ?
              reg389 : ({(reg382 ?
                      wire376 : wire379)} * reg384[(4'hc):(1'h0)])) : $unsigned(wire377[(1'h1):(1'h1)])))
        begin
          if ((~(&($unsigned($signed(reg392)) ?
              "iFz" : $unsigned($unsigned(reg388))))))
            begin
              reg393 <= wire375;
              reg394 <= ((~^wire378) ?
                  ({$signed("riV7nSA0M1otN")} ?
                      $signed((+"fdukatTtp9SUOGY3HzpgM")) : "P") : reg387[(4'hf):(4'he)]);
              reg395 <= $unsigned($unsigned("By"));
            end
          else
            begin
              reg393 = (((((7'h44) ? reg391 : "m") ?
                  ("oqbDGOvYc4C7n" ?
                      forvar383 : (+reg382)) : $signed(reg384)) * $unsigned($unsigned($signed(reg386)))) - ((reg393 ^~ reg386) << $signed("qnewgY88PII30i3FecxVU")));
            end
          if ($unsigned(reg385))
            begin
              reg396 <= reg391;
              reg397 = reg395;
              reg398 = $signed(((wire377[(1'h1):(1'h0)] < $signed("yAqG1aaincfxE343MynJo7")) ?
                  (&(-(|wire375))) : "gOFDyZW1sale"));
            end
          else
            begin
              reg396 <= "ZwAg";
              reg397 <= "7EMB74";
              reg398 <= $unsigned(((8'hbb) & ({(7'h42)} * $unsigned("YYroXPimstyhvmmAfF"))));
            end
          for (forvar399 = (1'h0); (forvar399 < (3'h4)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg400 <= {$signed("ouNmHwlixcg")};
              reg401 <= (|$unsigned(forvar390));
            end
          reg402 <= ((&($unsigned(wire375[(3'h4):(2'h3)]) ?
              wire377 : "QNUFgvkn6")) > (reg394 ?
              "5ELgMP3Dv2SlUv6" : {forvar399}));
        end
      else
        begin
          for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 <= reg386[(4'he):(4'hd)];
              reg395 <= wire377[(1'h0):(1'h0)];
              reg396 <= {($unsigned(wire378) <= (+((forvar383 ^~ reg398) != reg402)))};
              reg397 <= $unsigned((reg384 ?
                  $unsigned($signed(wire381[(4'hc):(2'h3)])) : "4ESpWIcY02OmMM5I"));
              reg398 <= $signed(reg402);
            end
          for (forvar399 = (1'h0); (forvar399 < (2'h3)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg400 = (!(7'h46));
              reg401 <= (((reg394 >>> $signed((reg383 != (8'hb0)))) >>> reg392) ?
                  (^(~&"zah7ADT")) : ((^(~|$unsigned(reg387))) && "BitVi9Qm6"));
            end
          reg402 <= wire379[(1'h0):(1'h0)];
        end
      reg403 <= (-(!($signed(forvar383) ?
          (reg391[(4'hc):(2'h2)] ?
              reg383 : (8'hbf)) : (((8'hb9) & wire377) >> {forvar393}))));
      for (forvar404 = (1'h0); (forvar404 < (1'h0)); forvar404 = (forvar404 + (1'h1)))
        begin
          if ((|{"oDa4O2u3Yu0uA"}))
            begin
              reg405 <= $signed($signed($unsigned($unsigned(reg386))));
              reg406 <= ($unsigned("4O7aPVvJd") >>> reg397[(4'hf):(4'h9)]);
            end
          else
            begin
              reg405 <= $signed(((forvar399 >>> $unsigned((reg405 ?
                      forvar382 : reg392))) ?
                  "R99zaTFqeaPxLWwdpn0" : ((|reg398[(4'hd):(3'h7)]) ?
                      "0vKIJLybX5ONRP3qoI3WL" : reg396)));
              reg406 <= $signed($unsigned($signed($signed($unsigned(reg394)))));
              reg407 <= $signed($signed({($signed((8'hba)) ~^ (~reg391)),
                  $signed($unsigned(reg389))}));
              reg408 <= reg385;
              reg409 <= reg382[(5'h12):(5'h12)];
            end
        end
    end
  always
    @(posedge clk) begin
      if (((~&"4SAUz1cZs1d3") ?
          $unsigned("kQJKqCzJLbPEHP0Z") : {(reg392 ?
                  $signed({reg385, (8'hb2)}) : reg391[(5'h10):(2'h2)]),
              (8'haf)}))
        begin
          reg410 <= reg388;
          for (forvar411 = (1'h0); (forvar411 < (2'h3)); forvar411 = (forvar411 + (1'h1)))
            begin
              reg412 <= reg388;
              reg413 <= (|$unsigned((~&wire381[(4'h8):(4'h8)])));
            end
        end
      else
        begin
          reg410 <= $signed(reg397[(3'h7):(3'h7)]);
        end
      for (forvar414 = (1'h0); (forvar414 < (1'h1)); forvar414 = (forvar414 + (1'h1)))
        begin
          for (forvar415 = (1'h0); (forvar415 < (2'h2)); forvar415 = (forvar415 + (1'h1)))
            begin
              reg416 <= reg398;
              reg417 <= reg403;
              reg418 <= forvar399[(3'h5):(2'h2)];
            end
          if (({reg388[(1'h0):(1'h0)]} <<< $signed($unsigned($unsigned("WzoNmhTK")))))
            begin
              reg419 <= (+($unsigned(forvar382) + $signed("IfrrhBcegewWICf")));
              reg420 <= (-reg391[(2'h3):(2'h3)]);
              reg421 <= ($unsigned($unsigned(($unsigned((8'hb9)) ?
                  reg383 : reg395))) >>> "y1h");
            end
          else
            begin
              reg419 <= "BE";
              reg420 = {(^wire377), reg391[(4'h8):(1'h1)]};
              reg421 <= (!wire375[(3'h7):(2'h3)]);
            end
          for (forvar422 = (1'h0); (forvar422 < (1'h0)); forvar422 = (forvar422 + (1'h1)))
            begin
              reg423 <= {((!reg420) ?
                      wire381 : (forvar404[(2'h3):(1'h0)] ?
                          $unsigned($signed(reg418)) : (~&"DurovCF48IJ"))),
                  ((((~&(8'had)) ~^ "z9GlBdIsUkVi167kZZI7a") ?
                      $unsigned((~(7'h42))) : $signed($signed(forvar422))) <<< $signed(forvar399[(2'h3):(1'h0)]))};
              reg424 <= $unsigned(reg395);
              reg425 = {(^{reg409[(4'hb):(1'h1)]})};
            end
          for (forvar426 = (1'h0); (forvar426 < (2'h2)); forvar426 = (forvar426 + (1'h1)))
            begin
              reg427 <= ((wire380[(4'h8):(1'h0)] ?
                  "BYnCeb8FdsKP" : (~^forvar411[(3'h4):(1'h1)])) ^~ $signed(reg389));
              reg428 <= $signed(((({reg386} ? "dGUxaRZZO" : "Z0831sP") ?
                      reg423[(1'h0):(1'h0)] : (reg384 & $signed(reg409))) ?
                  ({$signed(reg427)} << (8'hac)) : forvar393[(3'h7):(3'h5)]));
              reg429 <= ((~^{($unsigned(reg406) ?
                      "rIyhfnKY9YszBgAkCn" : (^reg409)),
                  ($signed((8'hb6)) ?
                      (reg420 ?
                          (7'h48) : forvar399) : "ukbF")}) <= (-(((7'h46) == (^forvar383)) ?
                  reg386[(2'h2):(1'h1)] : $unsigned((forvar390 ~^ reg400)))));
            end
          reg430 <= $unsigned("vL9XrHL7OIU3aZ2QuXF");
        end
      reg431 <= reg400[(3'h6):(2'h3)];
      for (forvar432 = (1'h0); (forvar432 < (2'h3)); forvar432 = (forvar432 + (1'h1)))
        begin
          if (({((forvar383[(4'h9):(4'h9)] ?
                  (reg417 ?
                      reg405 : (8'haf)) : ((8'hae) <<< forvar399)) >>> reg407)} != "7"))
            begin
              reg433 = $unsigned(($unsigned($unsigned((reg427 >> forvar411))) ?
                  ({forvar422} ? "7mKIogVnCd7wyX6Skt2" : "I") : "wIAzDRpfd"));
              reg434 <= $signed((!((8'ha3) >= (forvar426 ?
                  {reg418} : "mX8f3p5i"))));
              reg435 <= $unsigned($signed($signed($unsigned((reg394 && reg413)))));
            end
          else
            begin
              reg433 <= $unsigned(({"PspKm3bJHVJ", reg408[(1'h1):(1'h1)]} ?
                  reg408 : (reg384 | $signed((reg409 + reg385)))));
              reg434 <= ((+(forvar422[(5'h10):(2'h3)] || forvar382)) ?
                  (-$unsigned(((~^reg389) ?
                      (-(8'hab)) : forvar432))) : "IG7D2FW8F4IinY3uyH70uO");
              reg435 <= (+({forvar411} ?
                  ("TNaq5JC11EDz" << $unsigned("iAUV")) : (reg402[(2'h3):(2'h3)] ?
                      "w0ZvnH4x30nDVYQxo" : reg406[(2'h2):(2'h2)])));
              reg436 <= (~|reg395);
            end
          for (forvar437 = (1'h0); (forvar437 < (2'h3)); forvar437 = (forvar437 + (1'h1)))
            begin
              reg438 <= "MCNY";
              reg439 <= (^~$unsigned("WFBRsiT3AN3PUP2S"));
            end
          for (forvar440 = (1'h0); (forvar440 < (2'h2)); forvar440 = (forvar440 + (1'h1)))
            begin
              reg441 = "9wzfTXsL";
              reg442 <= $signed($signed(((^~(reg441 ? forvar393 : (8'hb0))) ?
                  ($signed((8'hbc)) ?
                      (^reg382) : (~forvar399)) : "0YK7vSATi")));
              reg443 <= $signed(reg439);
              reg444 <= ($signed("7z6eHKCBR") | $signed($unsigned(reg405[(3'h7):(3'h7)])));
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed($signed(reg438[(5'h11):(2'h2)])))
        begin
          for (forvar445 = (1'h0); (forvar445 < (2'h3)); forvar445 = (forvar445 + (1'h1)))
            begin
              reg446 <= ("I5MQW6" ~^ reg427[(3'h6):(2'h2)]);
              reg447 <= ("mE1C53Irgm5R" != $signed($unsigned(($signed(reg382) >>> (~(8'hae))))));
              reg448 <= "AXUBuFQSbk";
              reg449 <= "H";
              reg450 <= reg403;
            end
          if ((forvar390[(1'h0):(1'h0)] ~^ reg408))
            begin
              reg451 <= $signed($signed("ealD6"));
              reg452 <= wire376[(4'h8):(3'h6)];
            end
          else
            begin
              reg451 <= forvar393[(3'h7):(3'h5)];
              reg452 <= {(($unsigned("A4") >= ($signed(forvar445) ?
                      (reg407 ^~ (8'hab)) : reg425[(3'h6):(2'h2)])) <<< reg388[(1'h1):(1'h0)]),
                  (7'h41)};
            end
        end
      else
        begin
          for (forvar445 = (1'h0); (forvar445 < (1'h0)); forvar445 = (forvar445 + (1'h1)))
            begin
              reg446 <= $signed("");
              reg447 = reg436[(4'hb):(1'h0)];
              reg448 <= {{(+((wire381 ? reg419 : reg382) ?
                          "hYS0pPz3s5M0EO8vdGE" : (-wire381)))}};
              reg449 <= (^$signed((~|wire375[(2'h2):(1'h1)])));
              reg450 <= $signed({(7'h45),
                  ("" || ({reg425} ?
                      (reg400 ^ reg447) : "w98tJmRhbRnqadVN5Tlo"))});
            end
          if ((((~&reg397[(1'h1):(1'h0)]) ?
              reg417 : "CvEl3L7UtsH1IZwsZ48") - {{(reg449 >> $unsigned(reg405))}}))
            begin
              reg451 <= $signed((&"sBRe"));
            end
          else
            begin
              reg451 <= $signed({wire377,
                  (forvar422[(5'h13):(4'h9)] >>> (8'h9c))});
            end
          for (forvar452 = (1'h0); (forvar452 < (2'h3)); forvar452 = (forvar452 + (1'h1)))
            begin
              reg453 <= $signed(reg387[(5'h11):(1'h0)]);
              reg454 <= reg436;
              reg455 <= ("mTQ" >>> $unsigned("LnmwGEZ5nPRGb00Xg4sTT"));
              reg456 <= "91WK9";
              reg457 <= "SYsoWeVcH7ig1B0mXmfs";
            end
          reg458 <= ((~$unsigned(((-reg428) >= $unsigned((8'hbf))))) ?
              "HUok9Wr3kywNTpV9" : ({{(forvar437 != reg393)}} ?
                  (forvar445 <= ({(8'had)} * "BJygP37n8gx2")) : ({$unsigned(reg446)} ^~ ((+reg438) - (8'hbf)))));
        end
      if ((~^((7'h40) ?
          (reg424 ?
              ("lJIKkrD6WBN64W5iE4G" >= "7lXJeSIUhSmNLQkVQJAI") : "oBO7LaQN5dKqlpA2p") : reg451)))
        begin
          reg459 <= "";
        end
      else
        begin
          if ((reg397[(5'h11):(4'hf)] >> (reg395[(3'h7):(1'h0)] ^ "l56Hkt")))
            begin
              reg459 <= (+reg393[(3'h5):(2'h2)]);
              reg460 <= "1epgy6EM8JuJIGMIXY2";
              reg461 <= (~wire378);
            end
          else
            begin
              reg459 <= (8'ha0);
              reg460 <= ($signed((((forvar437 ?
                  (8'ha0) : reg406) - $unsigned(reg452)) == ((reg448 ^~ wire375) || (^reg393)))) | $unsigned((|"uVnrkHXkMV9NQZAva0Rzmf")));
            end
        end
    end
  assign wire462 = reg424;
  assign wire463 = (7'h47);
  assign wire464 = {{(reg401 & $signed("AxobZgvDvkwabu"))},
                       $unsigned($signed((|reg458[(2'h3):(1'h0)])))};
  assign wire465 = (~&$signed((8'ha0)));
  assign wire466 = ($signed((~^reg433)) ?
                       {$signed((~^$signed(reg389)))} : $signed((^reg388[(4'he):(4'h8)])));
  assign wire467 = $signed($unsigned($signed({(!reg459), $signed(reg387)})));
  always
    @(posedge clk) begin
      reg468 <= "sAGiUXaJne2XDZ31GsxIu3";
      for (forvar469 = (1'h0); (forvar469 < (1'h0)); forvar469 = (forvar469 + (1'h1)))
        begin
          reg470 <= (wire462[(2'h3):(1'h1)] <= $signed(reg428[(1'h1):(1'h0)]));
          reg471 <= $unsigned($signed(((reg392[(4'h8):(1'h1)] <= reg420[(3'h6):(2'h3)]) ?
              (^~$unsigned(forvar414)) : ("qk7gUXff" == {reg384, forvar382}))));
        end
    end
  assign wire472 = (|"w2qKPInQv");
endmodule