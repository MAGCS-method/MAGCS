module top
#(parameter param485 = ((^~({{(7'h43)}, {(8'hac)}} ? ((8'hb4) << {(7'h42), (8'hae)}) : (+(^~(8'hb1))))) ^~ (((|(&(8'hbd))) ? ({(8'ha4)} ? {(8'hb0)} : ((8'hbb) <<< (8'hba))) : ((-(8'h9e)) ? ((8'ha4) ? (8'ha2) : (8'hae)) : ((8'ha5) ? (8'hb4) : (8'hb4)))) ? (({(8'ha6)} ? ((8'ha5) ? (8'hb9) : (8'ha8)) : ((8'hbe) - (7'h43))) ? {(8'haa), {(8'ha4), (8'ha9)}} : ((+(8'ha8)) != ((8'hb4) ? (8'hba) : (7'h43)))) : (({(8'hb6), (8'haf)} ? (+(8'haa)) : ((8'ha3) ? (7'h42) : (8'h9f))) ? (~|(|(7'h43))) : {((8'hac) ? (8'hba) : (8'hb7))}))), 
parameter param486 = param485)
(y, clk, wire308, wire307, wire306, wire305);
  output wire [(32'h8cd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire308;
  input wire signed [(2'h2):(1'h0)] wire307;
  input wire signed [(4'h9):(1'h0)] wire306;
  input wire signed [(2'h3):(1'h0)] wire305;
  wire signed [(5'h14):(1'h0)] wire484;
  wire signed [(4'hb):(1'h0)] wire465;
  wire [(3'h5):(1'h0)] wire464;
  wire [(4'hc):(1'h0)] wire463;
  wire [(4'h8):(1'h0)] wire394;
  wire signed [(2'h2):(1'h0)] wire393;
  wire [(5'h10):(1'h0)] wire392;
  wire signed [(5'h14):(1'h0)] wire391;
  wire [(4'hf):(1'h0)] wire390;
  wire signed [(5'h14):(1'h0)] wire388;
  wire signed [(5'h15):(1'h0)] wire387;
  wire [(4'hc):(1'h0)] wire372;
  wire [(5'h13):(1'h0)] wire352;
  reg [(3'h6):(1'h0)] reg483 = (1'h0);
  reg [(3'h5):(1'h0)] reg482 = (1'h0);
  reg [(5'h11):(1'h0)] reg480 = (1'h0);
  reg [(2'h3):(1'h0)] reg479 = (1'h0);
  reg signed [(4'he):(1'h0)] reg478 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg475 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg471 = (1'h0);
  reg [(4'he):(1'h0)] reg469 = (1'h0);
  reg [(5'h11):(1'h0)] reg468 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg467 = (1'h0);
  reg [(5'h11):(1'h0)] reg461 = (1'h0);
  reg [(5'h10):(1'h0)] reg460 = (1'h0);
  reg [(4'hf):(1'h0)] reg459 = (1'h0);
  reg [(3'h4):(1'h0)] reg457 = (1'h0);
  reg [(5'h12):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg454 = (1'h0);
  reg [(4'hb):(1'h0)] reg453 = (1'h0);
  reg [(4'hb):(1'h0)] reg452 = (1'h0);
  reg [(5'h13):(1'h0)] reg451 = (1'h0);
  reg [(5'h15):(1'h0)] reg450 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg447 = (1'h0);
  reg [(5'h12):(1'h0)] reg446 = (1'h0);
  reg [(4'hd):(1'h0)] reg445 = (1'h0);
  reg [(5'h14):(1'h0)] reg443 = (1'h0);
  reg [(2'h3):(1'h0)] reg440 = (1'h0);
  reg [(5'h13):(1'h0)] reg439 = (1'h0);
  reg [(4'hb):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg433 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg428 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg426 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg423 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg422 = (1'h0);
  reg [(4'he):(1'h0)] reg421 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg420 = (1'h0);
  reg [(4'hb):(1'h0)] reg418 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg415 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg413 = (1'h0);
  reg [(5'h11):(1'h0)] reg409 = (1'h0);
  reg [(5'h15):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg407 = (1'h0);
  reg [(5'h15):(1'h0)] reg403 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg397 = (1'h0);
  reg signed [(4'he):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg389 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg386 = (1'h0);
  reg [(4'hc):(1'h0)] reg385 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg374 = (1'h0);
  reg [(5'h10):(1'h0)] reg380 = (1'h0);
  reg [(4'hd):(1'h0)] reg369 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg366 = (1'h0);
  reg [(3'h7):(1'h0)] reg362 = (1'h0);
  reg [(5'h14):(1'h0)] reg361 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg359 = (1'h0);
  reg [(5'h13):(1'h0)] reg358 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg357 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg356 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg355 = (1'h0);
  reg [(4'hc):(1'h0)] reg354 = (1'h0);
  reg [(3'h7):(1'h0)] reg351 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg349 = (1'h0);
  reg [(5'h12):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg339 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg338 = (1'h0);
  reg [(2'h2):(1'h0)] reg335 = (1'h0);
  reg signed [(4'he):(1'h0)] reg334 = (1'h0);
  reg [(5'h14):(1'h0)] reg332 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg329 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg319 = (1'h0);
  reg [(2'h3):(1'h0)] reg327 = (1'h0);
  reg [(2'h2):(1'h0)] reg326 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg324 = (1'h0);
  reg [(4'hb):(1'h0)] reg322 = (1'h0);
  reg [(5'h14):(1'h0)] reg321 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg320 = (1'h0);
  reg [(4'ha):(1'h0)] reg318 = (1'h0);
  reg [(4'hd):(1'h0)] reg317 = (1'h0);
  reg [(4'h9):(1'h0)] reg311 = (1'h0);
  reg [(5'h13):(1'h0)] reg309 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar481 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg470 = (1'h0);
  reg [(5'h11):(1'h0)] forvar468 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg477 = (1'h0);
  reg [(3'h7):(1'h0)] reg476 = (1'h0);
  reg [(3'h4):(1'h0)] reg474 = (1'h0);
  reg [(4'he):(1'h0)] reg473 = (1'h0);
  reg [(4'hf):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar470 = (1'h0);
  reg [(2'h2):(1'h0)] reg466 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg462 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg458 = (1'h0);
  reg [(4'h8):(1'h0)] forvar457 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar458 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg456 = (1'h0);
  reg [(4'ha):(1'h0)] reg449 = (1'h0);
  reg [(5'h15):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg444 = (1'h0);
  reg [(4'hb):(1'h0)] reg442 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar441 = (1'h0);
  reg [(4'h9):(1'h0)] forvar438 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg436 = (1'h0);
  reg [(3'h4):(1'h0)] forvar435 = (1'h0);
  reg [(3'h5):(1'h0)] reg434 = (1'h0);
  reg [(4'hf):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg431 = (1'h0);
  reg [(4'hb):(1'h0)] forvar430 = (1'h0);
  reg [(5'h13):(1'h0)] reg429 = (1'h0);
  reg [(4'h8):(1'h0)] reg427 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg425 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg424 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar419 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg417 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg414 = (1'h0);
  reg [(5'h11):(1'h0)] forvar412 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg411 = (1'h0);
  reg [(4'h9):(1'h0)] reg410 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar406 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar405 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg404 = (1'h0);
  reg [(5'h13):(1'h0)] reg402 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg401 = (1'h0);
  reg [(5'h12):(1'h0)] forvar399 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg395 = (1'h0);
  reg [(5'h15):(1'h0)] forvar382 = (1'h0);
  reg [(4'hb):(1'h0)] reg381 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg384 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg383 = (1'h0);
  reg [(5'h10):(1'h0)] reg382 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar381 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg379 = (1'h0);
  reg [(3'h4):(1'h0)] reg378 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg377 = (1'h0);
  reg [(5'h11):(1'h0)] reg376 = (1'h0);
  reg [(3'h7):(1'h0)] reg375 = (1'h0);
  reg [(4'ha):(1'h0)] forvar374 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg373 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg370 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg368 = (1'h0);
  reg signed [(4'he):(1'h0)] reg365 = (1'h0);
  reg signed [(4'he):(1'h0)] reg364 = (1'h0);
  reg [(5'h15):(1'h0)] reg363 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar353 = (1'h0);
  reg [(4'hd):(1'h0)] forvar343 = (1'h0);
  reg [(5'h15):(1'h0)] reg350 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg348 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg347 = (1'h0);
  reg [(4'he):(1'h0)] reg346 = (1'h0);
  reg [(5'h15):(1'h0)] reg345 = (1'h0);
  reg [(4'h8):(1'h0)] reg344 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg343 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg340 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg337 = (1'h0);
  reg [(5'h13):(1'h0)] reg336 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar333 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg328 = (1'h0);
  reg [(3'h4):(1'h0)] forvar318 = (1'h0);
  reg [(4'h9):(1'h0)] reg314 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg325 = (1'h0);
  reg [(3'h4):(1'h0)] reg323 = (1'h0);
  reg [(4'hb):(1'h0)] forvar319 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg316 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg315 = (1'h0);
  reg [(4'hd):(1'h0)] forvar314 = (1'h0);
  reg [(2'h2):(1'h0)] reg313 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg312 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg310 = (1'h0);
  assign y = {wire484,
                 wire465,
                 wire464,
                 wire463,
                 wire394,
                 wire393,
                 wire392,
                 wire391,
                 wire390,
                 wire388,
                 wire387,
                 wire372,
                 wire352,
                 reg483,
                 reg482,
                 reg480,
                 reg479,
                 reg478,
                 reg475,
                 reg471,
                 reg469,
                 reg468,
                 reg467,
                 reg461,
                 reg460,
                 reg459,
                 reg457,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg447,
                 reg446,
                 reg445,
                 reg443,
                 reg440,
                 reg439,
                 reg437,
                 reg433,
                 reg428,
                 reg426,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg418,
                 reg415,
                 reg413,
                 reg409,
                 reg408,
                 reg407,
                 reg403,
                 reg400,
                 reg398,
                 reg397,
                 reg396,
                 reg389,
                 reg386,
                 reg385,
                 reg374,
                 reg380,
                 reg369,
                 reg367,
                 reg366,
                 reg362,
                 reg361,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg351,
                 reg349,
                 reg342,
                 reg341,
                 reg339,
                 reg338,
                 reg335,
                 reg334,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg319,
                 reg327,
                 reg326,
                 reg324,
                 reg322,
                 reg321,
                 reg320,
                 reg318,
                 reg317,
                 reg311,
                 reg309,
                 forvar481,
                 reg470,
                 forvar468,
                 reg477,
                 reg476,
                 reg474,
                 reg473,
                 reg472,
                 forvar470,
                 reg466,
                 reg462,
                 reg458,
                 forvar457,
                 forvar458,
                 reg456,
                 reg449,
                 reg448,
                 reg444,
                 reg442,
                 forvar441,
                 forvar438,
                 reg436,
                 forvar435,
                 reg434,
                 reg432,
                 reg431,
                 forvar430,
                 reg429,
                 reg427,
                 reg425,
                 reg424,
                 forvar419,
                 reg417,
                 forvar416,
                 reg414,
                 forvar412,
                 reg411,
                 reg410,
                 forvar406,
                 forvar405,
                 reg404,
                 reg402,
                 reg401,
                 forvar399,
                 reg395,
                 forvar382,
                 reg381,
                 reg384,
                 reg383,
                 reg382,
                 forvar381,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 forvar374,
                 reg373,
                 reg371,
                 reg370,
                 reg368,
                 reg365,
                 reg364,
                 reg363,
                 reg360,
                 forvar353,
                 forvar343,
                 reg350,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg340,
                 reg337,
                 reg336,
                 forvar333,
                 reg328,
                 forvar318,
                 reg314,
                 reg325,
                 reg323,
                 forvar319,
                 reg316,
                 reg315,
                 forvar314,
                 reg313,
                 reg312,
                 reg310,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((^~$unsigned(($unsigned(wire306[(3'h5):(2'h2)]) >> wire305))))
        begin
          if ((wire306 | wire307[(2'h2):(1'h0)]))
            begin
              reg309 <= wire305;
              reg310 = (|wire306);
              reg311 <= reg309;
              reg312 = $unsigned($unsigned({((wire308 ? wire307 : wire307) ?
                      wire305[(2'h3):(2'h2)] : wire307[(1'h1):(1'h0)]),
                  wire307[(2'h2):(1'h1)]}));
              reg313 = $signed(($unsigned($signed(wire307)) ?
                  wire305 : (reg312 != ($unsigned(wire308) != (wire308 ?
                      wire307 : reg312)))));
            end
          else
            begin
              reg309 <= (7'h41);
              reg311 <= $unsigned($unsigned($signed(wire308)));
            end
          for (forvar314 = (1'h0); (forvar314 < (1'h1)); forvar314 = (forvar314 + (1'h1)))
            begin
              reg315 = forvar314;
              reg316 = reg315[(2'h3):(1'h1)];
              reg317 <= $unsigned($signed((reg315 * ($unsigned(reg315) ?
                  (~|reg316) : (reg313 ? wire306 : forvar314)))));
              reg318 <= $unsigned($unsigned($unsigned(($unsigned(reg313) == (^~(8'haa))))));
            end
          for (forvar319 = (1'h0); (forvar319 < (1'h0)); forvar319 = (forvar319 + (1'h1)))
            begin
              reg320 <= reg313;
              reg321 <= ({reg315[(1'h0):(1'h0)],
                  {{$unsigned(forvar314)}}} > (~(~^$unsigned(reg313))));
              reg322 <= $unsigned($unsigned((8'hb7)));
            end
          if (wire308)
            begin
              reg323 = $signed(($unsigned($signed($signed(wire308))) ?
                  reg312 : ($unsigned($unsigned(reg321)) ?
                      (~|wire305) : {reg312, $signed(reg311)})));
              reg324 <= (&reg312);
            end
          else
            begin
              reg323 = {$signed((($unsigned(reg322) ?
                      reg315 : (&reg311)) & reg317))};
              reg325 = $unsigned(wire305);
              reg326 <= ($unsigned((($unsigned(reg317) ?
                      reg309[(3'h6):(1'h0)] : reg309) ?
                  reg310[(2'h3):(2'h2)] : {(8'ha0)})) <= $unsigned((!$unsigned((reg310 ^ reg320)))));
              reg327 <= (^~$unsigned((((^~reg310) ?
                  $unsigned(reg325) : $signed(forvar319)) ^ $signed({reg322,
                  reg310}))));
            end
        end
      else
        begin
          if ((reg320 && $signed(reg322)))
            begin
              reg309 <= reg321;
              reg311 <= reg325;
              reg312 = {reg312[(3'h7):(3'h7)],
                  (reg325 | $signed(reg320[(3'h4):(1'h0)]))};
              reg313 = $unsigned(wire306[(2'h3):(2'h2)]);
              reg314 = $signed($unsigned(reg321));
            end
          else
            begin
              reg309 <= (~|$signed(forvar314[(4'hb):(4'hb)]));
              reg310 = (~&($signed((wire308 != $signed((8'ha5)))) <<< $unsigned(({reg322} | $unsigned(reg322)))));
              reg312 = forvar319;
              reg317 <= wire305;
            end
          for (forvar318 = (1'h0); (forvar318 < (2'h3)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg319 <= wire308;
              reg320 <= forvar318[(3'h4):(1'h1)];
              reg323 = $unsigned(forvar314);
            end
          reg324 <= wire305[(2'h2):(1'h1)];
          if ($signed($unsigned($unsigned(reg316[(2'h2):(2'h2)]))))
            begin
              reg326 <= (~&($signed($signed($unsigned(reg322))) ?
                  forvar314[(2'h2):(1'h1)] : ((~|(~|wire308)) - reg326)));
              reg328 = (({wire308[(3'h5):(2'h2)], wire305} >= (^(~^(reg318 ?
                      reg319 : (8'hbf))))) ?
                  reg313 : ((reg318[(3'h4):(3'h4)] ?
                      (-(reg322 ?
                          reg313 : reg327)) : (reg327 ^~ $unsigned(wire307))) || $signed(((reg316 && reg311) == reg311[(4'h9):(3'h4)]))));
              reg329 <= (wire305 ?
                  reg317[(1'h1):(1'h1)] : $unsigned($unsigned($signed((reg325 ?
                      reg324 : (8'h9c))))));
              reg330 <= $unsigned(((&(wire306 ?
                      $unsigned(wire306) : $unsigned((8'ha6)))) ?
                  reg322[(4'ha):(4'ha)] : wire308[(1'h0):(1'h0)]));
            end
          else
            begin
              reg326 <= (~^forvar319);
            end
        end
      reg331 <= reg313[(1'h0):(1'h0)];
      reg332 <= $signed((reg316[(3'h5):(3'h4)] ?
          reg318 : (+$signed($unsigned(reg313)))));
      for (forvar333 = (1'h0); (forvar333 < (2'h2)); forvar333 = (forvar333 + (1'h1)))
        begin
          reg334 <= reg321;
          if ((~|$unsigned({(~(reg325 ? reg332 : reg315)),
              $unsigned((reg325 >>> (8'ha3)))})))
            begin
              reg335 <= (reg321 ?
                  (^reg321[(1'h1):(1'h0)]) : (reg325 >> reg309));
              reg336 = $unsigned($unsigned((forvar314 ?
                  ($signed(reg309) >> {forvar333,
                      reg323}) : reg315[(2'h2):(1'h1)])));
              reg337 = reg324;
            end
          else
            begin
              reg335 <= reg309[(1'h0):(1'h0)];
              reg338 <= (($signed($signed($signed(reg327))) >= reg327[(2'h2):(2'h2)]) ?
                  wire307 : ($signed(reg323[(1'h1):(1'h0)]) ?
                      {forvar319} : reg314[(3'h5):(2'h2)]));
              reg339 <= reg331;
              reg340 = reg336;
            end
          reg341 <= ((reg329 ?
              reg338[(1'h0):(1'h0)] : $unsigned(reg321)) >>> (~$unsigned(($unsigned(reg337) ?
              {reg312, reg336} : (reg323 ? forvar318 : reg331)))));
          reg342 <= $unsigned((($unsigned($signed(reg316)) ^ reg321) == (($signed(reg313) - (reg324 ?
              reg322 : forvar314)) && $unsigned($signed(reg332)))));
        end
    end
  always
    @(posedge clk) begin
      if (($signed((reg318[(4'ha):(4'ha)] != ($unsigned(reg341) < $unsigned(reg332)))) ?
          ((^((wire307 == wire308) ?
              (~^reg319) : (~reg320))) >> wire306) : $unsigned($unsigned(wire306))))
        begin
          if ((-$signed($signed($unsigned({reg321})))))
            begin
              reg343 = reg331;
              reg344 = (-$unsigned((((8'hb9) ?
                  (reg339 ?
                      wire305 : reg334) : (wire306 - reg338)) <= $unsigned($unsigned(wire308)))));
              reg345 = $signed(({reg334, reg320[(2'h3):(1'h0)]} ?
                  reg319 : ($unsigned(reg335) ?
                      ($unsigned(reg331) ?
                          $unsigned(reg342) : reg344) : $unsigned(reg332))));
              reg346 = ((wire305 + wire308) ?
                  (~&$unsigned($unsigned({reg344,
                      (8'ha5)}))) : ($unsigned($unsigned($unsigned(reg338))) ?
                      reg345 : reg341));
            end
          else
            begin
              reg343 = (reg330[(5'h10):(5'h10)] ?
                  (&$unsigned($unsigned((8'h9d)))) : (reg346 ?
                      $unsigned({$signed(reg343),
                          $unsigned(reg331)}) : wire306));
            end
          if ($unsigned((~&reg320)))
            begin
              reg347 = $unsigned({reg341});
              reg348 = $signed(wire305);
              reg349 <= {$unsigned(reg341)};
              reg350 = (((((reg334 * reg342) ?
                      $unsigned(reg342) : (reg344 ?
                          reg322 : wire305)) ^~ reg318[(3'h5):(1'h0)]) + (~&(~^(+reg349)))) ?
                  reg326 : $signed(reg318));
            end
          else
            begin
              reg349 <= (&(reg341 ?
                  ({$unsigned(wire305)} ?
                      ((^wire305) ?
                          (|reg350) : reg318) : wire307[(1'h1):(1'h1)]) : $unsigned($unsigned($signed(reg344)))));
            end
        end
      else
        begin
          for (forvar343 = (1'h0); (forvar343 < (2'h2)); forvar343 = (forvar343 + (1'h1)))
            begin
              reg344 = reg318;
              reg349 <= ($unsigned($unsigned($unsigned($unsigned(reg331)))) | ($unsigned(reg309) < $signed((~^(reg329 ~^ (8'hb1))))));
              reg351 <= $unsigned($signed(reg322));
            end
        end
    end
  assign wire352 = (reg332[(5'h10):(4'h9)] ?
                       ($signed((^{reg326, reg319})) ?
                           (+$signed((reg339 <<< reg332))) : {reg317}) : reg329);
  always
    @(posedge clk) begin
      for (forvar353 = (1'h0); (forvar353 < (3'h4)); forvar353 = (forvar353 + (1'h1)))
        begin
          if (($signed($unsigned((^~$unsigned(reg331)))) ?
              $unsigned(reg326[(2'h2):(2'h2)]) : reg349))
            begin
              reg354 <= $unsigned($signed(reg349[(3'h7):(3'h7)]));
              reg355 <= ((8'hb2) ?
                  (~^{$unsigned({(8'ha8)})}) : (&($signed($unsigned(reg329)) ?
                      $unsigned((^~reg322)) : $unsigned($unsigned(wire308)))));
              reg356 <= $unsigned((!(8'ha5)));
              reg357 <= reg311;
              reg358 <= (!$unsigned($unsigned(forvar353)));
            end
          else
            begin
              reg354 <= $unsigned((~^$unsigned(reg357[(1'h0):(1'h0)])));
              reg355 <= reg351;
              reg356 <= reg321;
            end
          if ({$signed($unsigned((~^(8'ha0))))})
            begin
              reg359 <= (reg355[(1'h1):(1'h1)] ?
                  ($signed({(wire306 ?
                          reg331 : (8'hb1))}) & ($unsigned(reg351) ?
                      ({forvar353, (8'hb3)} ?
                          reg357 : $unsigned(reg329)) : {reg327[(2'h2):(2'h2)],
                          reg324[(2'h2):(2'h2)]})) : reg324);
              reg360 = {$signed(((reg311 & {reg327}) ?
                      $unsigned(wire306) : $unsigned((~|reg321)))),
                  (|(&$unsigned((reg320 + reg357))))};
            end
          else
            begin
              reg360 = wire352;
              reg361 <= reg342[(5'h10):(3'h7)];
              reg362 <= $unsigned($unsigned($unsigned(($unsigned(reg321) ?
                  ((7'h42) || reg309) : $signed(reg324)))));
              reg363 = reg359;
              reg364 = reg359[(4'hd):(4'h9)];
            end
          if ($signed(reg354[(1'h1):(1'h1)]))
            begin
              reg365 = ($unsigned(($signed($unsigned(wire306)) ?
                      reg359 : {wire352, (|reg351)})) ?
                  reg317 : $unsigned($unsigned((8'hb9))));
              reg366 <= {($unsigned(reg351) ?
                      $signed($signed(((8'hbc) >> reg311))) : reg360),
                  (~&(-$unsigned((^~reg338))))};
              reg367 <= $unsigned(reg334);
              reg368 = $signed($unsigned({$unsigned(reg363),
                  (reg342[(4'he):(3'h5)] ?
                      (reg318 ? wire306 : reg338) : (!reg349))}));
            end
          else
            begin
              reg366 <= reg318[(2'h3):(2'h2)];
              reg367 <= ((+((~&(reg330 ? reg335 : reg324)) ?
                  $unsigned((reg365 ?
                      reg355 : forvar353)) : reg364[(4'h8):(2'h3)])) && reg324);
              reg369 <= {($signed($unsigned($unsigned((8'ha0)))) ?
                      (~reg355) : (((reg338 & reg361) ^~ (+reg330)) ?
                          $signed({reg357, reg317}) : (reg359 >> reg327))),
                  (-($signed({reg365, forvar353}) ?
                      ($signed(reg361) ?
                          $signed(reg324) : $signed(reg365)) : ($signed(reg329) == reg359)))};
              reg370 = $signed(reg339[(4'h9):(2'h3)]);
              reg371 = $unsigned((reg355[(2'h2):(2'h2)] ?
                  wire306 : $unsigned($unsigned(reg321))));
            end
        end
    end
  assign wire372 = {$signed($unsigned(reg326)), reg334};
  always
    @(posedge clk) begin
      if ((wire307[(1'h1):(1'h1)] ?
          $unsigned(($signed(reg319) > $unsigned({reg309,
              reg366}))) : {$signed(($unsigned(wire307) + reg309[(5'h10):(4'hd)])),
              (((reg335 ?
                  reg362 : reg327) == $signed(reg327)) & reg309[(5'h12):(4'h8)])}))
        begin
          reg373 = $signed($unsigned(reg324[(5'h13):(4'he)]));
          for (forvar374 = (1'h0); (forvar374 < (1'h0)); forvar374 = (forvar374 + (1'h1)))
            begin
              reg375 = reg356;
            end
          reg376 = reg367;
          if ($unsigned({reg351, $signed(reg330)}))
            begin
              reg377 = $unsigned(((^{reg330, $unsigned(reg309)}) ?
                  reg342 : (reg355 * $unsigned((-reg355)))));
              reg378 = ($unsigned($signed((-reg329[(3'h6):(1'h1)]))) == reg334);
              reg379 = ($signed((~&{$signed(reg375),
                  (&reg318)})) >>> $unsigned(reg355[(1'h0):(1'h0)]));
            end
          else
            begin
              reg380 <= (-(reg356 ?
                  $unsigned($unsigned((reg366 ?
                      reg351 : wire352))) : ($signed($signed(reg326)) ?
                      wire372[(2'h3):(1'h0)] : $unsigned($signed(reg375)))));
            end
          for (forvar381 = (1'h0); (forvar381 < (2'h2)); forvar381 = (forvar381 + (1'h1)))
            begin
              reg382 = $unsigned((!$signed($unsigned((reg320 ?
                  reg341 : reg332)))));
              reg383 = reg351[(2'h3):(2'h2)];
              reg384 = $unsigned(wire352);
            end
        end
      else
        begin
          reg374 <= ($unsigned(((((8'hb9) - wire372) ?
                      $signed((8'ha4)) : reg341) ?
                  $unsigned(reg351) : ($unsigned(reg338) ?
                      {reg382, reg341} : (+reg384)))) ?
              (((~|$unsigned((8'haa))) ?
                      (~|reg376) : $signed(reg383[(3'h4):(2'h3)])) ?
                  $signed($unsigned((8'ha5))) : ($signed({wire352,
                      wire306}) <<< (~|$unsigned(reg383)))) : {reg322});
          reg375 = $unsigned(($unsigned(reg329) ?
              {$signed($unsigned(reg369))} : $unsigned((&$unsigned(reg326)))));
          reg380 <= $unsigned(($unsigned(($unsigned(reg342) ?
              {reg384, reg383} : reg357)) <= (^reg309)));
          reg381 = $unsigned(($unsigned(wire352) >= (($unsigned(reg380) == reg354) > $unsigned(reg326))));
          for (forvar382 = (1'h0); (forvar382 < (2'h3)); forvar382 = (forvar382 + (1'h1)))
            begin
              reg385 <= {(reg324 ?
                      $unsigned(($signed(reg339) ?
                          $unsigned(reg379) : $signed(reg309))) : $unsigned($signed(reg349))),
                  $unsigned({$signed((reg374 - reg377))})};
              reg386 <= ($unsigned(reg374) ?
                  $unsigned(reg341) : $signed((wire307 ?
                      {$signed(reg369)} : reg374)));
            end
        end
    end
  assign wire387 = $unsigned((reg326[(1'h1):(1'h1)] ?
                       $unsigned($signed(reg335[(1'h0):(1'h0)])) : (+{(reg335 >>> reg317)})));
  assign wire388 = (|((~&(|reg356)) ?
                       reg332 : ($signed(wire306[(3'h5):(3'h5)]) ?
                           (^(~reg326)) : $unsigned((7'h40)))));
  always
    @(posedge clk) begin
      reg389 <= reg356[(3'h6):(3'h6)];
    end
  assign wire390 = (&($unsigned((^~(reg326 ?
                       reg334 : reg329))) >= reg321[(5'h11):(2'h3)]));
  assign wire391 = $unsigned(wire372);
  assign wire392 = reg389;
  assign wire393 = (!$unsigned(reg332));
  assign wire394 = (~|$signed($unsigned(wire390)));
  always
    @(posedge clk) begin
      reg395 = reg349;
      reg396 <= $unsigned(reg367);
      reg397 <= (({(((8'hbc) ?
              wire306 : wire352) - wire393)} >>> $unsigned((reg351[(3'h5):(2'h2)] ?
          (reg369 >> wire372) : $unsigned(reg335)))) || ((reg322 ?
              $signed((reg366 ?
                  reg334 : reg386)) : ((reg380 > (8'hbc)) & (~&reg334))) ?
          {reg334} : reg309));
      reg398 <= reg309[(4'hc):(3'h7)];
      for (forvar399 = (1'h0); (forvar399 < (2'h3)); forvar399 = (forvar399 + (1'h1)))
        begin
          reg400 <= $signed((reg324 ?
              $unsigned(reg338[(1'h1):(1'h1)]) : $signed(((~^reg321) <<< (&reg334)))));
          reg401 = $unsigned($signed(wire308[(4'hc):(3'h4)]));
          reg402 = (reg362[(3'h6):(1'h0)] ?
              (~|wire387[(4'hf):(1'h1)]) : {$signed(wire387[(5'h12):(4'ha)])});
          reg403 <= reg386[(3'h5):(1'h0)];
          reg404 = (reg366 ? reg389 : (!$signed((!$unsigned(wire305)))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar405 = (1'h0); (forvar405 < (1'h1)); forvar405 = (forvar405 + (1'h1)))
        begin
          for (forvar406 = (1'h0); (forvar406 < (1'h1)); forvar406 = (forvar406 + (1'h1)))
            begin
              reg407 <= $unsigned($unsigned((reg317 <<< ($signed(reg322) << $unsigned((8'h9f))))));
              reg408 <= $signed($unsigned($unsigned(reg354)));
              reg409 <= $signed((reg311 - {$unsigned((wire308 ^ reg349))}));
              reg410 = reg330;
              reg411 = $signed(reg374[(4'ha):(3'h5)]);
            end
          for (forvar412 = (1'h0); (forvar412 < (2'h2)); forvar412 = (forvar412 + (1'h1)))
            begin
              reg413 <= reg339;
              reg414 = reg326;
              reg415 <= reg361;
            end
          for (forvar416 = (1'h0); (forvar416 < (2'h3)); forvar416 = (forvar416 + (1'h1)))
            begin
              reg417 = reg317;
              reg418 <= reg374;
            end
          for (forvar419 = (1'h0); (forvar419 < (2'h3)); forvar419 = (forvar419 + (1'h1)))
            begin
              reg420 <= $unsigned((8'hae));
              reg421 <= {reg359};
              reg422 <= $unsigned($unsigned(reg322));
              reg423 <= (^~($unsigned(forvar416) ?
                  (&$signed((reg320 ?
                      wire393 : reg320))) : $unsigned($unsigned(reg356[(3'h5):(1'h1)]))));
              reg424 = $unsigned(reg386);
            end
          if ((reg422[(1'h1):(1'h0)] >>> $unsigned(reg326[(2'h2):(1'h0)])))
            begin
              reg425 = reg403;
              reg426 <= reg414;
              reg427 = (+reg426);
              reg428 <= $unsigned(((((~reg331) ? forvar405 : {reg408}) ?
                      $signed((reg403 ?
                          reg380 : reg418)) : (&$unsigned(reg362))) ?
                  wire391[(3'h4):(1'h1)] : (reg309 <= {$unsigned(reg425)})));
              reg429 = (($unsigned({$signed(reg338)}) ?
                      (reg332 <<< ((^~(8'ha8)) ?
                          (wire308 ?
                              reg354 : reg413) : (!forvar405))) : reg321[(4'hb):(3'h4)]) ?
                  $signed(wire308[(4'h8):(3'h7)]) : wire307[(2'h2):(2'h2)]);
            end
          else
            begin
              reg425 = reg330[(3'h5):(2'h3)];
              reg426 <= $signed((!{reg415, {(reg359 > reg342)}}));
            end
        end
      for (forvar430 = (1'h0); (forvar430 < (3'h4)); forvar430 = (forvar430 + (1'h1)))
        begin
          reg431 = ((reg411 ?
              ($unsigned((&wire392)) ?
                  reg396[(4'ha):(1'h0)] : {reg396}) : (-reg318)) ~^ $signed($unsigned(reg358)));
          reg432 = $unsigned(($signed(((~^reg341) ?
                  reg342 : reg408[(5'h13):(5'h10)])) ?
              reg358[(4'ha):(1'h1)] : ($unsigned(reg369) ?
                  reg320[(2'h3):(1'h1)] : (~$signed(reg367)))));
          reg433 <= ((~reg366) ?
              (8'ha3) : $signed((reg423[(3'h7):(3'h5)] & reg324[(4'he):(4'ha)])));
          reg434 = (($unsigned($unsigned((~&reg327))) ?
                  (~$signed($signed((8'had)))) : (reg427 ?
                      reg389 : $unsigned(wire391[(3'h7):(3'h5)]))) ?
              (8'hbc) : wire305);
        end
    end
  always
    @(posedge clk) begin
      for (forvar435 = (1'h0); (forvar435 < (3'h4)); forvar435 = (forvar435 + (1'h1)))
        begin
          reg436 = {{$unsigned((~&reg341[(1'h0):(1'h0)]))}};
          reg437 <= {$signed($unsigned(reg327)),
              $unsigned(forvar435[(2'h2):(1'h1)])};
          for (forvar438 = (1'h0); (forvar438 < (3'h4)); forvar438 = (forvar438 + (1'h1)))
            begin
              reg439 <= reg338;
              reg440 <= ($signed(($signed($unsigned(reg349)) & reg356)) ^~ ({(wire392[(1'h1):(1'h0)] <= $unsigned(reg380))} - reg385));
            end
          for (forvar441 = (1'h0); (forvar441 < (2'h3)); forvar441 = (forvar441 + (1'h1)))
            begin
              reg442 = {(reg321 <<< {$unsigned($unsigned(reg335)), reg326})};
              reg443 <= {(!(!reg334))};
              reg444 = $signed((^~((^$signed((8'ha6))) ^~ reg338)));
            end
        end
      reg445 <= ((~&reg374[(3'h7):(3'h5)]) ?
          ($signed(forvar441) * $unsigned(reg362)) : reg369);
      if ((reg400[(1'h0):(1'h0)] ?
          $unsigned(((~reg356) ?
              (~(reg389 ? reg408 : wire308)) : {(wire388 + reg418),
                  reg361})) : (+$unsigned((-$unsigned(reg433))))))
        begin
          if ($unsigned({wire394}))
            begin
              reg446 <= $unsigned((^(((reg409 <<< reg309) ~^ $signed(reg339)) & reg332[(3'h7):(1'h1)])));
              reg447 <= (~&reg442);
              reg448 = (reg422 ? $signed(reg439) : reg440);
            end
          else
            begin
              reg448 = $unsigned(($signed((reg319[(3'h6):(2'h2)] >>> reg385[(2'h2):(1'h0)])) ?
                  {forvar438, (8'ha0)} : $unsigned(($signed(reg369) ?
                      (wire392 - reg420) : reg396[(1'h0):(1'h0)]))));
              reg449 = $unsigned(wire308[(2'h3):(2'h3)]);
              reg450 <= wire392;
              reg451 <= reg330;
              reg452 <= $signed(((-$unsigned($signed(forvar438))) < $unsigned($signed((&reg309)))));
            end
          reg453 <= reg332[(3'h5):(2'h2)];
          if (((reg396[(3'h6):(2'h3)] ?
              (^$signed(reg449)) : $unsigned((reg413[(3'h4):(1'h0)] ?
                  {reg439, reg409} : reg357))) && (8'hb7)))
            begin
              reg454 <= ($signed(wire392) ?
                  $unsigned(($signed($unsigned(reg449)) ?
                      ((reg367 ? reg317 : reg338) ?
                          {reg356} : reg385) : ({reg329, reg398} ?
                          $signed(wire308) : reg362))) : (~|(~|(+reg407[(4'hd):(4'h9)]))));
              reg455 <= ($signed($unsigned((8'hbb))) ?
                  ($unsigned($signed($unsigned(reg318))) > (^(reg442 >> (reg329 & reg319)))) : $signed(reg361[(4'ha):(1'h1)]));
              reg456 = (~&reg334);
            end
          else
            begin
              reg454 <= (reg447 ?
                  (reg440 ~^ reg374) : (|reg326[(1'h1):(1'h0)]));
              reg456 = reg409;
              reg457 <= {((~((&reg447) ?
                      {wire352} : $signed(reg366))) > reg361[(4'h8):(2'h2)]),
                  wire392};
            end
          for (forvar458 = (1'h0); (forvar458 < (2'h3)); forvar458 = (forvar458 + (1'h1)))
            begin
              reg459 <= {reg413,
                  $unsigned((reg334 >> ($unsigned(reg367) ?
                      wire393 : reg420)))};
              reg460 <= (!wire390);
            end
        end
      else
        begin
          if ((reg407[(4'hd):(3'h4)] | reg357[(3'h5):(1'h1)]))
            begin
              reg448 = reg318[(3'h6):(3'h4)];
              reg449 = $unsigned((reg389[(3'h5):(3'h4)] ?
                  reg457 : $unsigned($unsigned({reg415, reg389}))));
            end
          else
            begin
              reg446 <= (reg455 ?
                  ({reg361} && $signed($unsigned(reg367))) : reg359);
              reg447 <= reg403;
              reg450 <= (~$unsigned($unsigned($signed((~&reg361)))));
            end
          reg456 = (reg361 ? reg329 : reg440[(2'h2):(1'h1)]);
          for (forvar457 = (1'h0); (forvar457 < (2'h3)); forvar457 = (forvar457 + (1'h1)))
            begin
              reg458 = wire394;
            end
          reg459 <= $signed(reg413);
        end
      reg461 <= ($unsigned($unsigned(reg322)) ?
          (reg459 ?
              ($signed(((8'ha6) ? wire372 : reg433)) ?
                  {reg436} : reg318[(4'ha):(2'h3)]) : ($unsigned($unsigned(reg403)) >> reg457)) : reg356);
      reg462 = ((|($signed($signed(reg324)) * reg446)) < ((wire305 ?
          wire352[(4'hf):(3'h7)] : (reg317 ?
              $unsigned(reg437) : (8'hac))) & (~|(((8'hb3) ^~ reg436) > (~^forvar458)))));
    end
  assign wire463 = $unsigned(($unsigned(reg341) ?
                       (($unsigned(reg324) >>> wire392[(1'h0):(1'h0)]) ?
                           reg433 : (reg361 ?
                               {reg403, reg339} : (reg355 ?
                                   reg420 : reg457))) : $unsigned((8'hbf))));
  assign wire464 = ((reg421[(3'h4):(3'h4)] ?
                           (reg318 ?
                               ((wire372 ? wire307 : (8'hbe)) ?
                                   reg453[(2'h3):(1'h1)] : (~&reg457)) : reg454[(4'h9):(3'h4)]) : wire352) ?
                       $unsigned($unsigned({$signed(reg421)})) : $unsigned(reg386[(4'hb):(2'h2)]));
  assign wire465 = (^~reg327);
  always
    @(posedge clk) begin
      reg466 = (8'hbc);
      reg467 <= reg317;
      if (($unsigned((!reg413[(4'hf):(3'h4)])) ^~ (reg437 != wire465[(4'h8):(3'h6)])))
        begin
          reg468 <= $signed((^(~|$unsigned(wire394[(3'h6):(2'h2)]))));
          reg469 <= ($signed(($unsigned(((8'hb0) & reg451)) ?
              reg322[(3'h6):(1'h1)] : $unsigned(reg408))) << $signed(reg443));
          for (forvar470 = (1'h0); (forvar470 < (1'h0)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 <= (&(reg452 != ($signed($signed(reg354)) > $signed($signed((8'h9c))))));
              reg472 = ({$unsigned(reg455),
                      ($signed((reg461 ? reg403 : wire392)) >= {(!wire393)})} ?
                  $signed(reg457[(1'h0):(1'h0)]) : (7'h44));
              reg473 = $signed((((wire308 ?
                      (reg366 ? reg332 : reg349) : $signed(reg469)) ?
                  (!$signed(reg471)) : reg413) > reg366));
              reg474 = (reg361[(4'hf):(4'ha)] ~^ reg334);
              reg475 <= $unsigned($signed($unsigned(wire372[(4'hc):(4'h8)])));
            end
          if (reg339)
            begin
              reg476 = $signed($unsigned(((8'haa) ?
                  $signed((reg386 | wire463)) : ({reg339, reg454} ?
                      $signed((8'hb9)) : $signed(reg447)))));
              reg477 = reg459;
              reg478 <= ((+(~^$signed((reg477 ?
                  reg440 : wire372)))) <<< reg331);
              reg479 <= $unsigned((reg374[(2'h2):(2'h2)] ?
                  wire464[(1'h0):(1'h0)] : reg466[(1'h0):(1'h0)]));
            end
          else
            begin
              reg476 = {{reg418, (reg330 * (|reg403))},
                  (reg322 ?
                      (reg459 ?
                          (reg342[(4'h9):(3'h4)] ?
                              $signed(reg398) : reg459) : reg475) : (8'ha2))};
            end
          reg480 <= $signed(reg329);
        end
      else
        begin
          for (forvar468 = (1'h0); (forvar468 < (1'h0)); forvar468 = (forvar468 + (1'h1)))
            begin
              reg470 = reg439;
              reg472 = $unsigned(reg445);
              reg473 = $signed(reg361);
            end
        end
      for (forvar481 = (1'h0); (forvar481 < (1'h1)); forvar481 = (forvar481 + (1'h1)))
        begin
          reg482 <= $unsigned(reg470[(2'h2):(2'h2)]);
        end
      reg483 <= reg447;
    end
  assign wire484 = (~|(reg469[(3'h4):(3'h4)] != $unsigned($unsigned(reg357[(2'h2):(1'h1)]))));
endmodule
