(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param3487 = ((((((7'h57) >= (8'hba)) == ((8'hb6) ? (8'ha3) : (8'hb8))) ^~ (~^((8'h9d) && (8'ha3)))) ? (+(~|((8'h9e) ? (8'hb5) : (8'ha7)))) : ((((7'h50) ? (8'hbb) : (7'h54)) ? ((8'hb9) ? (7'h4b) : (8'ha8)) : {(8'hb8), (8'haf), (8'had)}) ? ({(8'hb7)} > {(8'hb9), (8'hac), (8'hb0)}) : (+((7'h58) + (7'h54))))) ? {({((8'hbd) ? (8'had) : (8'hbd)), {(8'hb9), (8'hb0)}, {(7'h4f)}} ? (((7'h52) > (8'ha5)) >> (-(7'h50))) : (((7'h4d) ? (7'h51) : (8'hbc)) ? (~|(7'h54)) : (!(8'hb9)))), (((|(8'hb2)) ? (7'h49) : ((7'h4b) >= (8'hb7))) ? {((7'h54) ? (8'hb0) : (8'hab)), {(8'ha6)}} : (((8'ha8) ? (8'had) : (8'ha1)) ? (&(8'hab)) : ((8'hab) ? (8'hab) : (8'haf)))), (|(~^((8'hab) ? (8'ha3) : (8'ha7))))} : {(!((-(8'ha7)) ^~ (!(8'hab)))), {({(8'hac)} ? ((7'h4f) ? (8'ha3) : (8'ha9)) : (~&(8'hbb))), {{(7'h40), (8'hb8)}, ((8'h9c) < (7'h50)), ((8'hb9) ? (8'hbf) : (7'h50))}}, (({(8'hb7), (8'hb5), (8'hb6)} && (^~(7'h53))) >> (~((8'hb3) ? (7'h45) : (7'h4c))))}), 
parameter param3488 = (~&param3487))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h15d1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h19):(1'h0)] wire0;
  input wire [(5'h1e):(1'h0)] wire1;
  input wire [(5'h12):(1'h0)] wire2;
  input wire [(5'h13):(1'h0)] wire3;
  wire signed [(3'h7):(1'h0)] wire3485;
  wire signed [(3'h5):(1'h0)] wire1685;
  wire signed [(5'h1a):(1'h0)] wire1577;
  wire signed [(2'h2):(1'h0)] wire1576;
  wire [(4'hb):(1'h0)] wire1446;
  wire [(5'h15):(1'h0)] wire1444;
  reg [(5'h19):(1'h0)] reg1684 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1681 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1679 = (1'h0);
  reg [(5'h13):(1'h0)] reg1678 = (1'h0);
  reg [(4'h8):(1'h0)] reg1677 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1676 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1674 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1672 = (1'h0);
  reg [(4'h9):(1'h0)] reg1668 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1666 = (1'h0);
  reg [(3'h4):(1'h0)] reg1665 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1664 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1663 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1661 = (1'h0);
  reg [(5'h16):(1'h0)] reg1658 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1651 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1648 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1647 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1642 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1639 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1638 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1636 = (1'h0);
  reg [(3'h7):(1'h0)] reg1632 = (1'h0);
  reg [(3'h6):(1'h0)] reg1629 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1627 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1620 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1617 = (1'h0);
  reg [(3'h6):(1'h0)] reg1615 = (1'h0);
  reg [(4'hc):(1'h0)] reg1614 = (1'h0);
  reg [(3'h4):(1'h0)] reg1613 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1611 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1604 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1602 = (1'h0);
  reg [(4'hb):(1'h0)] reg1601 = (1'h0);
  reg [(5'h15):(1'h0)] reg1600 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1596 = (1'h0);
  reg [(5'h17):(1'h0)] reg1594 = (1'h0);
  reg [(5'h19):(1'h0)] reg1593 = (1'h0);
  reg [(3'h6):(1'h0)] reg1589 = (1'h0);
  reg [(4'hf):(1'h0)] reg1585 = (1'h0);
  reg [(4'h8):(1'h0)] reg1583 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1581 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1575 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1574 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1568 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1567 = (1'h0);
  reg [(2'h3):(1'h0)] reg1566 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1563 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1561 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1560 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1559 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1556 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1555 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1553 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1552 = (1'h0);
  reg [(3'h7):(1'h0)] reg1551 = (1'h0);
  reg [(5'h10):(1'h0)] reg1550 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1549 = (1'h0);
  reg [(4'he):(1'h0)] reg1547 = (1'h0);
  reg [(3'h6):(1'h0)] reg1545 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1544 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1541 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1536 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1533 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1532 = (1'h0);
  reg [(4'h9):(1'h0)] reg1530 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1528 = (1'h0);
  reg [(4'he):(1'h0)] reg1504 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1524 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1523 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1520 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1519 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1517 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1516 = (1'h0);
  reg [(4'h8):(1'h0)] reg1514 = (1'h0);
  reg [(3'h4):(1'h0)] reg1513 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1510 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1506 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1505 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1502 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1497 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1496 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1495 = (1'h0);
  reg [(4'hf):(1'h0)] reg1493 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1492 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1472 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1488 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1487 = (1'h0);
  reg [(4'hc):(1'h0)] reg1483 = (1'h0);
  reg [(5'h12):(1'h0)] reg1482 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1481 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1479 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1477 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1476 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1473 = (1'h0);
  reg [(4'he):(1'h0)] reg1471 = (1'h0);
  reg [(4'hf):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1466 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1465 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1464 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1459 = (1'h0);
  reg [(4'ha):(1'h0)] reg1457 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1456 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1453 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1451 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1447 = (1'h0);
  reg [(5'h16):(1'h0)] reg89 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg86 = (1'h0);
  reg [(5'h10):(1'h0)] reg84 = (1'h0);
  reg [(3'h5):(1'h0)] reg82 = (1'h0);
  reg [(5'h16):(1'h0)] reg81 = (1'h0);
  reg [(5'h11):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg78 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg75 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg67 = (1'h0);
  reg [(5'h17):(1'h0)] reg66 = (1'h0);
  reg [(3'h6):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg60 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg59 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg58 = (1'h0);
  reg [(4'hc):(1'h0)] reg57 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg56 = (1'h0);
  reg [(3'h7):(1'h0)] reg53 = (1'h0);
  reg [(4'hd):(1'h0)] reg51 = (1'h0);
  reg [(5'h1c):(1'h0)] reg50 = (1'h0);
  reg [(3'h7):(1'h0)] reg49 = (1'h0);
  reg [(5'h13):(1'h0)] reg43 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg46 = (1'h0);
  reg [(5'h1b):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg38 = (1'h0);
  reg [(4'hd):(1'h0)] reg31 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg28 = (1'h0);
  reg [(5'h15):(1'h0)] reg27 = (1'h0);
  reg [(5'h16):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg21 = (1'h0);
  reg [(5'h11):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg11 = (1'h0);
  reg [(4'hd):(1'h0)] reg10 = (1'h0);
  reg [(5'h10):(1'h0)] reg7 = (1'h0);
  reg [(4'ha):(1'h0)] reg5 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1683 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1682 = (1'h0);
  reg [(5'h15):(1'h0)] reg1680 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1675 = (1'h0);
  reg [(2'h3):(1'h0)] reg1673 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1671 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1670 = (1'h0);
  reg [(3'h7):(1'h0)] reg1669 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1664 = (1'h0);
  reg [(2'h3):(1'h0)] reg1667 = (1'h0);
  reg [(5'h10):(1'h0)] reg1662 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1660 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1659 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1657 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1656 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1655 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1654 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1653 = (1'h0);
  reg [(4'h9):(1'h0)] reg1652 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1650 = (1'h0);
  reg [(5'h12):(1'h0)] reg1649 = (1'h0);
  reg [(5'h14):(1'h0)] reg1646 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1645 = (1'h0);
  reg [(5'h13):(1'h0)] reg1644 = (1'h0);
  reg [(3'h7):(1'h0)] reg1643 = (1'h0);
  reg [(5'h18):(1'h0)] reg1641 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1640 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1637 = (1'h0);
  reg [(4'h8):(1'h0)] reg1635 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1634 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1633 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1631 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1630 = (1'h0);
  reg [(4'ha):(1'h0)] reg1628 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1626 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1625 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1624 = (1'h0);
  reg [(4'hd):(1'h0)] reg1623 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1622 = (1'h0);
  reg [(2'h2):(1'h0)] reg1621 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1619 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1618 = (1'h0);
  reg [(4'hd):(1'h0)] reg1616 = (1'h0);
  reg [(2'h3):(1'h0)] reg1612 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1610 = (1'h0);
  reg [(5'h15):(1'h0)] reg1609 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1608 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1607 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1606 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1605 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar1603 = (1'h0);
  reg [(5'h17):(1'h0)] reg1599 = (1'h0);
  reg [(3'h5):(1'h0)] reg1598 = (1'h0);
  reg [(4'hb):(1'h0)] reg1597 = (1'h0);
  reg [(4'hc):(1'h0)] reg1595 = (1'h0);
  reg [(4'hf):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1591 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1590 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1582 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1588 = (1'h0);
  reg [(4'he):(1'h0)] reg1587 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1586 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1584 = (1'h0);
  reg [(4'hd):(1'h0)] reg1582 = (1'h0);
  reg [(4'h8):(1'h0)] reg1580 = (1'h0);
  reg [(5'h14):(1'h0)] reg1579 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1578 = (1'h0);
  reg [(4'h9):(1'h0)] reg1573 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1572 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1571 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1570 = (1'h0);
  reg [(4'he):(1'h0)] reg1569 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1565 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1564 = (1'h0);
  reg [(5'h12):(1'h0)] reg1562 = (1'h0);
  reg [(5'h15):(1'h0)] reg1558 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1557 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1554 = (1'h0);
  reg [(5'h14):(1'h0)] reg1548 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1546 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1543 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1542 = (1'h0);
  reg [(5'h13):(1'h0)] reg1540 = (1'h0);
  reg [(5'h17):(1'h0)] reg1539 = (1'h0);
  reg [(4'h9):(1'h0)] reg1538 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1537 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1535 = (1'h0);
  reg [(3'h7):(1'h0)] reg1534 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1531 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1529 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1527 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1526 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1515 = (1'h0);
  reg [(5'h14):(1'h0)] reg1498 = (1'h0);
  reg [(4'h8):(1'h0)] reg1525 = (1'h0);
  reg [(5'h13):(1'h0)] reg1522 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1521 = (1'h0);
  reg [(3'h7):(1'h0)] reg1518 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1515 = (1'h0);
  reg [(4'hf):(1'h0)] reg1512 = (1'h0);
  reg [(3'h4):(1'h0)] reg1511 = (1'h0);
  reg [(4'h9):(1'h0)] reg1509 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1508 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1507 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1504 = (1'h0);
  reg [(5'h14):(1'h0)] reg1503 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1501 = (1'h0);
  reg [(4'hf):(1'h0)] reg1500 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1499 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1498 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1494 = (1'h0);
  reg [(5'h11):(1'h0)] reg1491 = (1'h0);
  reg [(5'h14):(1'h0)] reg1490 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1489 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar1485 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1484 = (1'h0);
  reg [(4'hd):(1'h0)] reg1486 = (1'h0);
  reg [(3'h7):(1'h0)] reg1485 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1484 = (1'h0);
  reg [(5'h14):(1'h0)] reg1480 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1478 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1475 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1474 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar1472 = (1'h0);
  reg [(5'h18):(1'h0)] reg1470 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1468 = (1'h0);
  reg [(5'h16):(1'h0)] reg1467 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1463 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1462 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1461 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1460 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1458 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1450 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1455 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1454 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1452 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1450 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1449 = (1'h0);
  reg [(2'h3):(1'h0)] reg1448 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg91 = (1'h0);
  reg [(4'hb):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg87 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg83 = (1'h0);
  reg [(5'h13):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg76 = (1'h0);
  reg [(3'h4):(1'h0)] forvar74 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar73 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg71 = (1'h0);
  reg [(5'h1b):(1'h0)] reg70 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg68 = (1'h0);
  reg [(5'h17):(1'h0)] reg65 = (1'h0);
  reg [(4'ha):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar54 = (1'h0);
  reg [(2'h3):(1'h0)] reg52 = (1'h0);
  reg [(4'ha):(1'h0)] reg48 = (1'h0);
  reg [(4'h9):(1'h0)] reg47 = (1'h0);
  reg [(4'hc):(1'h0)] reg45 = (1'h0);
  reg [(4'hb):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar43 = (1'h0);
  reg [(5'h19):(1'h0)] reg42 = (1'h0);
  reg [(5'h1f):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg39 = (1'h0);
  reg [(3'h4):(1'h0)] reg37 = (1'h0);
  reg [(5'h1e):(1'h0)] reg36 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg34 = (1'h0);
  reg signed [(4'he):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg32 = (1'h0);
  reg [(3'h5):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg29 = (1'h0);
  reg [(3'h5):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg23 = (1'h0);
  reg [(4'hf):(1'h0)] forvar22 = (1'h0);
  reg [(4'hc):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar17 = (1'h0);
  reg [(5'h1d):(1'h0)] reg16 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg15 = (1'h0);
  reg [(5'h11):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar9 = (1'h0);
  reg [(2'h3):(1'h0)] reg8 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar6 = (1'h0);
  reg [(5'h16):(1'h0)] forvar4 = (1'h0);
  assign y = {wire3485,
                 wire1685,
                 wire1577,
                 wire1576,
                 wire1446,
                 wire1444,
                 reg1684,
                 reg1681,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1674,
                 reg1672,
                 reg1668,
                 reg1666,
                 reg1665,
                 reg1664,
                 reg1663,
                 reg1661,
                 reg1658,
                 reg1651,
                 reg1648,
                 reg1647,
                 reg1642,
                 reg1639,
                 reg1638,
                 reg1636,
                 reg1632,
                 reg1629,
                 reg1627,
                 reg1620,
                 reg1617,
                 reg1615,
                 reg1614,
                 reg1613,
                 reg1611,
                 reg1604,
                 reg1602,
                 reg1601,
                 reg1600,
                 reg1596,
                 reg1594,
                 reg1593,
                 reg1589,
                 reg1585,
                 reg1583,
                 reg1581,
                 reg1575,
                 reg1574,
                 reg1568,
                 reg1567,
                 reg1566,
                 reg1563,
                 reg1561,
                 reg1560,
                 reg1559,
                 reg1556,
                 reg1555,
                 reg1553,
                 reg1552,
                 reg1551,
                 reg1550,
                 reg1549,
                 reg1547,
                 reg1545,
                 reg1544,
                 reg1541,
                 reg1536,
                 reg1533,
                 reg1532,
                 reg1530,
                 reg1528,
                 reg1504,
                 reg1524,
                 reg1523,
                 reg1520,
                 reg1519,
                 reg1517,
                 reg1516,
                 reg1514,
                 reg1513,
                 reg1510,
                 reg1506,
                 reg1505,
                 reg1502,
                 reg1497,
                 reg1496,
                 reg1495,
                 reg1493,
                 reg1492,
                 reg1472,
                 reg1488,
                 reg1487,
                 reg1483,
                 reg1482,
                 reg1481,
                 reg1479,
                 reg1477,
                 reg1476,
                 reg1473,
                 reg1471,
                 reg1469,
                 reg1466,
                 reg1465,
                 reg1464,
                 reg1459,
                 reg1457,
                 reg1456,
                 reg1453,
                 reg1451,
                 reg1447,
                 reg89,
                 reg86,
                 reg84,
                 reg82,
                 reg81,
                 reg79,
                 reg78,
                 reg75,
                 reg67,
                 reg66,
                 reg64,
                 reg63,
                 reg62,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg53,
                 reg51,
                 reg50,
                 reg49,
                 reg43,
                 reg46,
                 reg40,
                 reg38,
                 reg31,
                 reg28,
                 reg27,
                 reg25,
                 reg21,
                 reg20,
                 reg14,
                 reg11,
                 reg10,
                 reg7,
                 reg5,
                 reg1683,
                 reg1682,
                 reg1680,
                 reg1675,
                 reg1673,
                 reg1671,
                 reg1670,
                 reg1669,
                 forvar1664,
                 reg1667,
                 reg1662,
                 reg1660,
                 reg1659,
                 reg1657,
                 reg1656,
                 reg1655,
                 reg1654,
                 reg1653,
                 reg1652,
                 reg1650,
                 reg1649,
                 reg1646,
                 reg1645,
                 reg1644,
                 reg1643,
                 reg1641,
                 reg1640,
                 reg1637,
                 reg1635,
                 reg1634,
                 forvar1633,
                 forvar1631,
                 reg1630,
                 reg1628,
                 reg1626,
                 reg1625,
                 forvar1624,
                 reg1623,
                 reg1622,
                 reg1621,
                 forvar1619,
                 forvar1618,
                 reg1616,
                 reg1612,
                 reg1610,
                 reg1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 forvar1605,
                 forvar1603,
                 reg1599,
                 reg1598,
                 reg1597,
                 reg1595,
                 reg1592,
                 reg1591,
                 reg1590,
                 forvar1582,
                 reg1588,
                 reg1587,
                 reg1586,
                 reg1584,
                 reg1582,
                 reg1580,
                 reg1579,
                 reg1578,
                 reg1573,
                 forvar1572,
                 forvar1571,
                 reg1570,
                 reg1569,
                 forvar1565,
                 reg1564,
                 reg1562,
                 reg1558,
                 reg1557,
                 reg1554,
                 reg1548,
                 reg1546,
                 reg1543,
                 reg1542,
                 reg1540,
                 reg1539,
                 reg1538,
                 reg1537,
                 reg1535,
                 reg1534,
                 reg1531,
                 reg1529,
                 forvar1527,
                 reg1526,
                 reg1515,
                 reg1498,
                 reg1525,
                 reg1522,
                 forvar1521,
                 reg1518,
                 forvar1515,
                 reg1512,
                 reg1511,
                 reg1509,
                 reg1508,
                 reg1507,
                 forvar1504,
                 reg1503,
                 reg1501,
                 reg1500,
                 reg1499,
                 forvar1498,
                 reg1494,
                 reg1491,
                 reg1490,
                 reg1489,
                 forvar1485,
                 reg1484,
                 reg1486,
                 reg1485,
                 forvar1484,
                 reg1480,
                 reg1478,
                 reg1475,
                 reg1474,
                 forvar1472,
                 reg1470,
                 reg1468,
                 reg1467,
                 reg1463,
                 reg1462,
                 reg1461,
                 reg1460,
                 forvar1458,
                 forvar1450,
                 reg1455,
                 reg1454,
                 reg1452,
                 reg1450,
                 reg1449,
                 reg1448,
                 reg91,
                 reg90,
                 reg88,
                 reg87,
                 reg85,
                 reg83,
                 reg80,
                 reg77,
                 reg76,
                 forvar74,
                 forvar73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg65,
                 reg61,
                 reg55,
                 forvar54,
                 reg52,
                 reg48,
                 reg47,
                 reg45,
                 reg44,
                 forvar43,
                 reg42,
                 reg41,
                 reg39,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg30,
                 reg29,
                 reg26,
                 reg24,
                 reg23,
                 forvar22,
                 reg19,
                 reg18,
                 forvar17,
                 reg16,
                 reg15,
                 reg13,
                 reg12,
                 forvar9,
                 reg8,
                 forvar6,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (2'h2)); forvar4 = (forvar4 + (1'h1)))
        begin
          reg5 <= ((8'haf) >= ({($signed((8'hba)) <<< forvar4[(5'h12):(3'h6)])} * $signed($unsigned((wire1 >= wire2)))));
          for (forvar6 = (1'h0); (forvar6 < (1'h0)); forvar6 = (forvar6 + (1'h1)))
            begin
              reg7 <= forvar4;
              reg8 = reg7[(4'ha):(3'h5)];
            end
          for (forvar9 = (1'h0); (forvar9 < (3'h4)); forvar9 = (forvar9 + (1'h1)))
            begin
              reg10 <= forvar6;
              reg11 <= (~^$signed((!forvar6[(1'h0):(1'h0)])));
              reg12 = forvar9[(4'hd):(1'h0)];
              reg13 = $unsigned(wire3[(2'h2):(2'h2)]);
              reg14 <= reg5;
              reg15 = ((reg5 ?
                  {(~(wire3 ?
                          reg8 : reg5))} : (7'h57)) ~^ forvar9[(5'h10):(4'ha)]);
              reg16 = (($unsigned($unsigned($signed(forvar9))) ?
                  reg8 : $signed(((forvar6 >>> reg11) ^~ forvar6[(5'h10):(4'h8)]))) & $unsigned(reg15[(3'h5):(3'h5)]));
            end
          for (forvar17 = (1'h0); (forvar17 < (3'h4)); forvar17 = (forvar17 + (1'h1)))
            begin
              reg18 = {(forvar9 ?
                      {(reg15 ^~ wire3), (|(reg13 <= reg8))} : forvar9),
                  {$signed(reg13[(1'h1):(1'h1)]),
                      (-{((7'h4a) ? wire2 : wire3),
                          $signed(reg5),
                          $signed(reg15)}),
                      ($signed(reg13[(4'h8):(4'h8)]) ?
                          ((reg14 ?
                              reg15 : forvar6) - (^~reg5)) : {$unsigned(reg15)})}};
              reg19 = reg7;
              reg20 <= wire3[(4'h9):(2'h3)];
              reg21 <= reg13;
            end
          for (forvar22 = (1'h0); (forvar22 < (1'h1)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 = $signed(reg18);
              reg24 = reg13[(3'h5):(1'h0)];
              reg25 <= (7'h47);
              reg26 = ($signed(wire2) >>> {($unsigned(reg8[(2'h3):(1'h1)]) * (~^$signed(forvar4))),
                  ($unsigned(forvar17) > $unsigned(forvar9[(2'h3):(1'h0)]))});
              reg27 <= ($signed((-(~&{reg23}))) ?
                  (+$signed(reg7[(1'h1):(1'h1)])) : (!(((~^reg13) > reg11) ?
                      (^~reg21) : ((reg11 >> reg15) ?
                          (wire1 == wire3) : ((8'hb4) ? reg13 : (8'h9e))))));
              reg28 <= (7'h40);
              reg29 = $unsigned(reg10[(1'h0):(1'h0)]);
            end
        end
      if (((reg8 ?
              $signed($signed({reg14, reg27})) : (-((reg11 ?
                  reg26 : forvar22) >> (+reg26)))) ?
          ((reg26[(3'h4):(2'h2)] ?
              forvar6 : ($unsigned(forvar17) < (+reg13))) | reg26) : {wire1[(4'h9):(3'h4)],
              (~^{reg25, (reg27 ? (8'hbd) : (8'hb0))}),
              reg11[(4'hf):(4'hd)]}))
        begin
          reg30 = ($signed(forvar22) ?
              (reg5[(3'h5):(2'h2)] || ($signed((wire1 ?
                  (8'hbb) : wire3)) | reg24[(4'h8):(3'h6)])) : reg16[(3'h4):(3'h4)]);
          reg31 <= ({(forvar4 > {{reg12, reg8, reg28}}), reg21[(4'hf):(1'h1)]} ?
              (8'ha3) : (~|({$unsigned(reg25), reg30, reg10} ?
                  ($unsigned(reg15) >> reg7[(4'hc):(3'h5)]) : reg24)));
          reg32 = $unsigned(reg7);
          reg33 = $signed(reg30);
          if (reg8)
            begin
              reg34 = (reg25 ?
                  wire3[(5'h10):(3'h7)] : (($signed((reg16 || reg18)) ?
                          (~^forvar22[(4'hf):(3'h7)]) : (reg10[(3'h7):(1'h0)] ?
                              ((7'h56) ?
                                  wire2 : reg12) : reg23[(5'h11):(3'h7)])) ?
                      ($unsigned((reg8 ?
                          reg18 : reg11)) >> (|wire1[(4'he):(2'h3)])) : (((^~forvar22) ?
                              reg23 : $unsigned(reg8)) ?
                          $signed($signed(forvar9)) : ($signed(reg32) ?
                              $signed(forvar22) : $unsigned(reg14)))));
              reg35 = $unsigned({(reg24 & (((7'h4d) ^ reg27) ?
                      forvar9[(5'h1d):(4'hf)] : (wire3 ? reg23 : wire1))),
                  ((reg27 ? $signed(forvar9) : (~&reg26)) ?
                      $signed((reg21 ? reg10 : reg32)) : reg29)});
              reg36 = $signed({$unsigned(($signed((8'had)) && $signed(reg11))),
                  (reg29 ^ $unsigned((reg7 ^~ reg23))),
                  (((~reg10) ? wire3 : forvar9) ?
                      {$signed(wire2)} : ({reg23} ?
                          $signed(reg31) : (reg16 ? forvar9 : forvar6)))});
              reg37 = (~^(+$signed(reg7[(4'h8):(4'h8)])));
              reg38 <= reg18;
              reg39 = reg8;
            end
          else
            begin
              reg34 = ((~$unsigned(reg33)) > reg14);
              reg38 <= (reg20[(2'h3):(1'h1)] ~^ (reg14 ?
                  reg8[(2'h3):(1'h0)] : ($unsigned(reg10) ?
                      reg19 : (~&(reg36 ? reg19 : (7'h41))))));
              reg39 = reg18[(1'h0):(1'h0)];
              reg40 <= ($signed((-forvar22[(1'h1):(1'h0)])) ?
                  reg27 : $signed(($unsigned($signed(reg20)) ?
                      (!reg8[(2'h3):(1'h0)]) : {reg10,
                          $unsigned(wire2),
                          forvar9})));
              reg41 = ($unsigned((7'h45)) ?
                  {($unsigned((wire0 <= reg35)) ?
                          {((7'h56) ?
                                  reg34 : forvar9)} : ($signed(reg32) * reg29[(5'h1a):(5'h16)])),
                      (+reg40)} : (|(((reg5 != reg35) ?
                      forvar6 : forvar9[(4'ha):(4'h8)]) - $unsigned((reg28 >> reg32)))));
              reg42 = ((((forvar4[(5'h16):(2'h3)] - reg36) ?
                      ((|forvar17) >= {reg8,
                          (7'h49)}) : reg13[(4'hf):(4'he)]) == ($unsigned((reg38 <= reg11)) ?
                      reg16 : ($signed(forvar4) && (~reg10)))) ?
                  $signed((wire2[(3'h4):(1'h0)] ^~ $unsigned(reg36))) : (((8'hab) ?
                      (~((7'h41) ?
                          reg26 : reg7)) : $unsigned((+reg7))) >= $signed(forvar6)));
            end
          for (forvar43 = (1'h0); (forvar43 < (3'h6)); forvar43 = (forvar43 + (1'h1)))
            begin
              reg44 = {reg11[(4'h9):(4'h9)],
                  (+({$signed(reg12), forvar17[(4'ha):(3'h5)], (|(7'h48))} ?
                      $signed(((8'haa) == forvar9)) : reg37)),
                  (~^((!reg37) ?
                      (forvar6[(4'he):(4'h8)] ?
                          reg16[(2'h2):(2'h2)] : $signed(reg10)) : {$signed(forvar9)}))};
              reg45 = (&reg7);
              reg46 <= reg24[(2'h2):(1'h1)];
              reg47 = $signed((+(^~({forvar17} ?
                  (forvar9 << (8'hbc)) : (+(8'h9e))))));
              reg48 = $signed(reg42);
            end
        end
      else
        begin
          reg31 <= (((8'hb8) ?
              (~|$unsigned(reg39[(1'h0):(1'h0)])) : reg29[(5'h1b):(1'h1)]) + reg29);
          reg32 = reg20;
          reg33 = $signed((($signed($unsigned(reg34)) ?
                  reg8[(1'h0):(1'h0)] : $unsigned(reg29[(5'h1b):(5'h17)])) ?
              $signed($signed($signed(reg10))) : $signed($signed((reg46 << (7'h43))))));
          if ({(reg35[(2'h2):(1'h1)] ?
                  $unsigned(reg48[(3'h6):(2'h2)]) : (!(&$signed(reg11))))})
            begin
              reg34 = (!reg37);
              reg38 <= {$signed($unsigned(({forvar43,
                      (8'hb2)} == $unsigned(reg35)))),
                  reg39,
                  ((reg16 ?
                      (|$signed(reg20)) : reg20) <<< reg35[(1'h1):(1'h1)])};
              reg39 = ((~|(^~$unsigned($unsigned((7'h54))))) - $signed($unsigned($unsigned((-reg19)))));
              reg40 <= forvar4[(3'h7):(1'h1)];
            end
          else
            begin
              reg38 <= (reg31 != ((reg31[(4'ha):(4'ha)] ?
                      ($unsigned(forvar6) ?
                          (reg12 * reg48) : ((8'hb6) ~^ reg7)) : (8'had)) ?
                  (!($signed((8'h9f)) ^ reg30)) : (({wire3,
                          reg32} * reg25[(3'h7):(2'h3)]) ?
                      ((+reg12) ?
                          forvar6 : $unsigned(reg45)) : $unsigned($unsigned(forvar43)))));
              reg39 = reg25[(4'he):(4'h8)];
              reg40 <= (forvar6[(3'h5):(3'h4)] ?
                  $unsigned($unsigned($signed((-(7'h52))))) : {$signed($signed((reg23 ?
                          reg12 : reg21))),
                      (reg40[(3'h4):(3'h4)] - reg19[(2'h2):(1'h1)])});
              reg43 <= (-{wire3,
                  $unsigned($signed(reg28[(2'h2):(1'h1)])),
                  reg46});
              reg44 = (reg11 * (!(reg21 ?
                  (+forvar43[(1'h1):(1'h0)]) : ($unsigned(reg7) * {(8'hb5),
                      reg41}))));
              reg45 = ($signed({(~|(reg41 ? reg39 : reg31)),
                  reg47}) <= reg27[(2'h3):(1'h0)]);
              reg47 = reg31[(1'h1):(1'h0)];
            end
          reg49 <= (+($unsigned({wire1}) ?
              $unsigned(reg43[(4'h8):(1'h1)]) : $signed(wire0)));
          reg50 <= (7'h55);
          reg51 <= reg26[(3'h5):(3'h5)];
        end
      reg52 = $unsigned((^reg10));
    end
  always
    @(posedge clk) begin
      if (((~($signed($signed(reg5)) ? (8'ha1) : (~&(reg27 * reg40)))) ?
          (wire0[(4'h9):(3'h5)] | {reg10[(3'h4):(2'h2)],
              $signed(((8'hbe) * reg25)),
              (~reg49[(2'h2):(1'h0)])}) : ((((~&(8'haa)) | (^reg28)) ?
              ($signed(reg46) <= (~|reg21)) : ($unsigned(reg49) ?
                  reg5[(4'h8):(3'h5)] : (reg10 ?
                      reg28 : (8'hb2)))) > ($signed((reg20 >> (7'h4a))) >= reg11))))
        begin
          reg53 <= reg25[(4'ha):(3'h7)];
        end
      else
        begin
          reg53 <= reg10[(3'h7):(3'h5)];
        end
      for (forvar54 = (1'h0); (forvar54 < (3'h6)); forvar54 = (forvar54 + (1'h1)))
        begin
          if ($unsigned($unsigned((reg11[(4'h8):(3'h7)] ^ ($unsigned(wire1) * (wire2 ?
              reg50 : reg49))))))
            begin
              reg55 = (($signed($signed(reg49)) ?
                      $unsigned(reg7[(3'h4):(1'h1)]) : (+$unsigned((reg38 - reg38)))) ?
                  ($unsigned(((8'haa) ?
                      $signed(reg21) : $unsigned(reg21))) ~^ {$signed($unsigned(reg7)),
                      (|$signed(reg7))}) : {wire0});
              reg56 <= reg50;
            end
          else
            begin
              reg56 <= (^(~&$signed((reg53 == reg50))));
              reg57 <= $signed(wire3);
              reg58 <= ((!(~(((7'h40) * reg49) ? $unsigned((7'h4d)) : reg7))) ?
                  ({wire2} ?
                      ((8'hbf) ?
                          ($unsigned(reg5) ?
                              $signed((8'h9c)) : $unsigned(reg50)) : ($signed(reg27) != $unsigned(reg55))) : $unsigned($unsigned($signed(reg10)))) : $signed(reg31));
              reg59 <= (~|reg46);
              reg60 <= $unsigned((~|{$signed($unsigned((8'ha1))),
                  reg11[(4'h9):(3'h6)],
                  $unsigned((reg14 != reg58))}));
              reg61 = ($unsigned($signed($signed((reg60 ?
                  wire1 : forvar54)))) * (reg43[(4'hc):(4'hb)] ?
                  ($signed(reg20) * (~((8'hbf) >> reg25))) : reg43));
              reg62 <= (7'h40);
            end
          reg63 <= wire0[(3'h5):(2'h3)];
          if (reg20)
            begin
              reg64 <= wire1[(1'h1):(1'h0)];
              reg65 = (reg14 && $unsigned((|forvar54[(2'h2):(1'h0)])));
            end
          else
            begin
              reg64 <= reg20[(2'h3):(2'h3)];
              reg65 = $unsigned({reg64[(3'h6):(1'h0)],
                  $unsigned(reg57[(1'h0):(1'h0)]),
                  $signed((7'h4b))});
              reg66 <= wire1;
              reg67 <= {$signed(((reg62 ^ $unsigned(reg10)) ?
                      forvar54[(2'h3):(1'h1)] : $signed(((8'hbb) & reg62))))};
              reg68 = {($unsigned(reg49[(3'h4):(1'h0)]) ?
                      (reg28 <<< $unsigned((^~wire3))) : (|{(reg14 || (7'h51)),
                          $unsigned(reg10)})),
                  $signed(((reg61[(3'h5):(3'h5)] >>> (reg40 ?
                          (7'h53) : (8'ha1))) ?
                      $signed($signed(reg10)) : $signed((reg38 <= reg57)))),
                  $signed($signed((|(reg63 ? reg28 : (7'h47)))))};
            end
          reg69 = (|$signed($signed(reg65)));
          reg70 = (reg46 >> ($unsigned($signed(reg20[(4'hd):(3'h5)])) ?
              {reg10} : $unsigned(reg28)));
          if ($signed($unsigned(((~|(forvar54 | reg31)) - $signed($signed(reg40))))))
            begin
              reg71 = {reg69, reg46};
            end
          else
            begin
              reg71 = reg20;
              reg72 = ($signed(reg62[(3'h4):(3'h4)]) > $signed(reg58));
            end
        end
      for (forvar73 = (1'h0); (forvar73 < (2'h3)); forvar73 = (forvar73 + (1'h1)))
        begin
          for (forvar74 = (1'h0); (forvar74 < (3'h4)); forvar74 = (forvar74 + (1'h1)))
            begin
              reg75 <= $unsigned(reg31[(4'h8):(3'h7)]);
              reg76 = (({(reg72[(2'h3):(1'h1)] ?
                      reg69 : $signed(reg27))} >= {reg46[(3'h7):(1'h1)],
                  reg62,
                  ((reg7 ^~ reg68) || reg49)}) * reg56[(4'h8):(2'h2)]);
            end
          reg77 = ($unsigned(((~$signed(reg55)) ?
                  ($signed((8'h9c)) != $signed((7'h40))) : (reg76 ?
                      (reg38 ? reg75 : reg5) : (reg68 >> reg31)))) ?
              (reg49 ?
                  reg61[(2'h2):(2'h2)] : $unsigned(reg31)) : ((~reg38) || ({forvar54[(4'h9):(3'h7)],
                  ((7'h41) ? reg21 : forvar73),
                  (7'h54)} | reg61)));
          if (((($signed((reg51 ?
              wire0 : reg38)) >>> (7'h50)) & $signed({reg53})) <<< reg7))
            begin
              reg78 <= (~&$unsigned(reg75));
              reg79 <= (({reg28, (|$unsigned(wire0)), $unsigned(reg51)} ?
                  wire1 : (reg46[(3'h7):(3'h6)] ?
                      (^~$signed(wire2)) : $signed((reg64 >> reg7)))) ^~ ((~$signed($unsigned(reg31))) < (reg76 >= ((reg51 || (8'hac)) ?
                  (^reg63) : (reg20 <= reg58)))));
            end
          else
            begin
              reg80 = (!{$signed((^~(reg28 && reg56))),
                  $signed((^~reg20[(2'h3):(2'h3)]))});
              reg81 <= $signed((reg75 != {$unsigned($unsigned(reg75))}));
            end
          if ({reg10})
            begin
              reg82 <= ({reg25, (7'h41), $unsigned((~{reg14}))} ?
                  $unsigned(forvar74) : wire2[(4'h9):(3'h6)]);
            end
          else
            begin
              reg82 <= $unsigned((reg51 > $signed(((~^reg7) ?
                  (reg70 | reg38) : (reg76 <= reg28)))));
              reg83 = $unsigned($unsigned(reg56[(1'h0):(1'h0)]));
              reg84 <= $signed((~^{(~&$signed(reg76)),
                  (^(reg56 ? reg72 : (7'h56)))}));
              reg85 = (($unsigned((wire2[(2'h2):(1'h0)] & (^wire1))) ?
                  $unsigned((~(|(8'hbc)))) : $signed(($signed(reg76) < $unsigned(reg38)))) << (reg63[(4'h9):(2'h3)] >>> ({(~|reg55),
                  reg49[(1'h1):(1'h0)],
                  {reg78, reg50}} >>> (reg72[(2'h3):(2'h2)] ?
                  (reg65 ? forvar54 : (7'h45)) : $unsigned(reg59)))));
            end
          if ($unsigned((((~^$signed(reg49)) ?
                  ((reg62 >> reg77) - $unsigned(reg5)) : ((reg76 ?
                          reg11 : wire0) ?
                      reg80 : (reg51 ? reg56 : reg51))) ?
              (reg58 ?
                  reg49[(3'h6):(1'h1)] : $signed((~^reg38))) : {($unsigned(forvar54) ?
                      reg84 : (reg61 << reg40)),
                  (^wire2[(2'h3):(1'h0)])})))
            begin
              reg86 <= {(reg59[(2'h3):(2'h2)] ? (!reg65) : reg5),
                  $signed($unsigned($unsigned($unsigned(reg21))))};
              reg87 = reg82[(2'h2):(1'h0)];
              reg88 = $signed(forvar54);
            end
          else
            begin
              reg86 <= (reg75 ?
                  reg68[(4'hd):(3'h7)] : (reg63 << ((+{reg86, reg75, reg60}) ?
                      $unsigned($unsigned(reg82)) : (~&(reg14 ?
                          reg61 : reg43)))));
              reg87 = forvar54;
              reg88 = reg28[(1'h0):(1'h0)];
              reg89 <= ((^((~|reg86[(1'h1):(1'h1)]) ?
                  $unsigned($unsigned(reg7)) : (~^wire1[(4'ha):(3'h6)]))) == $unsigned($unsigned($signed((reg84 >>> (7'h48))))));
              reg90 = reg84[(3'h6):(2'h3)];
            end
        end
      reg91 = ($unsigned(($unsigned(reg62[(2'h3):(1'h1)]) ?
          $signed($signed(reg76)) : ((~(8'ha7)) <<< (reg90 ?
              reg71 : wire1)))) >= (-reg49[(1'h1):(1'h1)]));
    end
  module92 #() modinst1445 (.y(wire1444), .clk(clk), .wire96(reg14), .wire97(reg43), .wire94(reg21), .wire93(wire1), .wire95(reg38));
  assign wire1446 = (^~wire2[(5'h10):(2'h3)]);
  always
    @(posedge clk) begin
      if (reg84)
        begin
          reg1447 <= {$unsigned((^~($unsigned((8'h9c)) ^ (reg5 <<< reg84))))};
          reg1448 = (reg25 - (reg66[(1'h0):(1'h0)] ?
              (($signed(reg43) ?
                  (~&reg86) : ((7'h43) == reg40)) || reg59[(3'h5):(1'h1)]) : reg10[(4'h9):(2'h2)]));
          if ((8'ha8))
            begin
              reg1449 = $signed((!$unsigned(((~(7'h48)) ?
                  (~&reg1447) : reg62))));
              reg1450 = (+(~|wire0[(3'h6):(2'h2)]));
              reg1451 <= {$unsigned($signed((+wire2[(1'h0):(1'h0)]))),
                  reg38[(4'h9):(1'h1)],
                  ($signed(reg28) * ((reg51 != (~reg86)) ?
                      wire1446 : ((reg82 ? reg21 : reg5) + $unsigned(reg20))))};
              reg1452 = (reg28 ? reg57[(2'h2):(1'h0)] : $unsigned(reg56));
              reg1453 <= {reg67[(3'h7):(1'h1)], reg79[(4'hc):(4'hc)]};
              reg1454 = $signed({reg1447[(4'hf):(4'hd)],
                  ((^~reg78) ?
                      ((reg5 ? (8'hbf) : wire1) ?
                          reg25 : {reg10}) : $signed(reg57[(4'ha):(3'h6)])),
                  ((~|reg53[(3'h6):(3'h5)]) - reg1453[(5'h16):(5'h10)])});
              reg1455 = wire2[(4'ha):(4'ha)];
            end
          else
            begin
              reg1449 = reg53[(1'h1):(1'h0)];
              reg1451 <= ({{$signed((reg66 ? reg81 : wire1446)),
                          reg62[(1'h0):(1'h0)]},
                      ($signed(reg84) ?
                          $signed({reg25,
                              reg62,
                              reg60}) : $unsigned($unsigned(reg78))),
                      (reg1447 ?
                          reg89 : (reg84[(4'ha):(4'h8)] ?
                              reg75[(2'h3):(2'h2)] : reg11))} ?
                  reg81 : $signed(reg40));
              reg1453 <= (($signed((((7'h51) ? (7'h44) : reg20) ?
                  $signed((7'h56)) : (reg58 ?
                      wire1444 : (8'hb2)))) ^ reg89[(3'h6):(3'h6)]) ^ $signed((7'h4e)));
            end
          reg1456 <= {(7'h4e)};
        end
      else
        begin
          reg1448 = (-(~&$unsigned($signed((^~reg84)))));
          reg1449 = reg82;
          for (forvar1450 = (1'h0); (forvar1450 < (2'h2)); forvar1450 = (forvar1450 + (1'h1)))
            begin
              reg1452 = reg62;
              reg1453 <= reg1448[(2'h3):(1'h1)];
              reg1456 <= reg1451;
              reg1457 <= ((~&((((7'h4f) ~^ reg20) != reg58) <= $signed((reg66 ?
                      reg49 : reg31)))) ?
                  reg64 : $signed(reg51));
            end
          for (forvar1458 = (1'h0); (forvar1458 < (2'h3)); forvar1458 = (forvar1458 + (1'h1)))
            begin
              reg1459 <= (reg51[(4'hc):(2'h3)] ?
                  {reg49[(2'h3):(2'h3)],
                      wire1444,
                      (-$signed((reg21 >> reg89)))} : ($signed(reg5) ?
                      $unsigned((~&$unsigned(reg57))) : reg43));
              reg1460 = ({{((reg62 ? reg1456 : reg1449) ?
                          reg14 : (reg1457 ~^ reg1450))},
                  reg84[(2'h3):(2'h3)],
                  (^~reg51)} && (reg27[(4'hd):(4'hb)] < $signed((~&(-reg84)))));
              reg1461 = $unsigned((~(reg89[(2'h3):(1'h1)] || reg78[(5'h13):(3'h6)])));
              reg1462 = ((reg28 + {$unsigned($unsigned(wire3)),
                      $signed({reg84}),
                      reg49}) ?
                  (!{reg89[(3'h6):(3'h4)],
                      (wire3[(4'hf):(3'h7)] * $signed(reg50)),
                      ((wire1 || reg56) ?
                          reg1447[(5'h13):(1'h0)] : reg25[(5'h10):(3'h4)])}) : reg5);
            end
          reg1463 = $unsigned(reg1449);
        end
    end
  always
    @(posedge clk) begin
      if ($signed(reg25[(4'h9):(3'h6)]))
        begin
          if ((~^$signed((reg5[(1'h0):(1'h0)] ?
              $signed($signed(reg79)) : reg49[(3'h7):(3'h7)]))))
            begin
              reg1464 <= ((($unsigned((!reg1447)) ?
                      {(reg1456 ?
                              reg20 : (7'h58))} : ($unsigned(reg1457) - $signed(reg21))) ?
                  wire1[(5'h17):(4'hc)] : $signed(((^~wire2) * wire0))) ^ ((^~wire1444) ^ $unsigned(wire1444[(4'ha):(3'h7)])));
              reg1465 <= {(^~reg81[(3'h5):(2'h3)])};
              reg1466 <= reg1464;
              reg1467 = reg1464;
              reg1468 = reg43;
              reg1469 <= ({$unsigned((-reg81))} ?
                  $signed(reg27) : wire0[(2'h3):(2'h2)]);
              reg1470 = (~$unsigned(reg89[(5'h14):(1'h1)]));
            end
          else
            begin
              reg1464 <= {$unsigned(((reg43[(3'h4):(1'h0)] ?
                          (reg50 <<< wire1) : (reg28 ? reg1470 : (8'hb7))) ?
                      (reg62[(3'h6):(3'h4)] * $signed((8'ha8))) : reg78[(1'h1):(1'h1)]))};
              reg1467 = reg63;
              reg1469 <= $signed(reg1469);
              reg1471 <= reg1451;
            end
          for (forvar1472 = (1'h0); (forvar1472 < (2'h2)); forvar1472 = (forvar1472 + (1'h1)))
            begin
              reg1473 <= (&(!($unsigned((|reg57)) <<< reg79[(2'h2):(1'h1)])));
              reg1474 = (reg67[(3'h4):(3'h4)] ?
                  ({$unsigned((!reg1456)),
                      reg28[(1'h0):(1'h0)],
                      {reg86}} + reg14) : (~|$unsigned(reg56)));
              reg1475 = ($unsigned(reg49[(1'h1):(1'h1)]) ?
                  ($signed((^(reg7 <= reg31))) && (~&(((7'h4e) ?
                          reg62 : reg31) ?
                      (wire3 ?
                          reg82 : reg82) : (8'ha6)))) : reg84[(4'hf):(3'h7)]);
              reg1476 <= $unsigned($unsigned(reg59[(1'h0):(1'h0)]));
              reg1477 <= reg1474;
              reg1478 = $unsigned((((8'ha9) ?
                      $signed({reg1469,
                          (8'hba),
                          reg51}) : reg1451[(5'h1b):(5'h13)]) ?
                  {($signed(reg56) ^ (7'h52))} : reg1465[(5'h15):(2'h2)]));
              reg1479 <= ((~|reg1470) >= (&$unsigned((~&$signed(wire1446)))));
            end
          reg1480 = (($unsigned($signed(reg56)) << (8'ha2)) ?
              $unsigned((({reg1474} <= (^~wire0)) ?
                  (8'hbe) : {(~&reg1473)})) : (reg21[(5'h14):(5'h13)] ?
                  ((^~(reg86 * reg58)) < reg1478[(1'h1):(1'h0)]) : $unsigned(reg31[(4'h9):(2'h2)])));
          reg1481 <= (|wire1[(5'h1d):(5'h19)]);
          reg1482 <= ($signed({reg1467}) * ((({wire3, reg57, (8'hb4)} ?
                  ((7'h49) * reg58) : reg1471) ?
              reg1457 : $unsigned($unsigned(wire3))) || wire2[(4'he):(3'h7)]));
          reg1483 <= reg63[(5'h1b):(4'hc)];
          for (forvar1484 = (1'h0); (forvar1484 < (1'h1)); forvar1484 = (forvar1484 + (1'h1)))
            begin
              reg1485 = ((($signed((8'hbb)) ?
                      $unsigned((reg82 <= reg1464)) : (&reg21[(5'h10):(1'h1)])) ?
                  $unsigned({(reg1467 ?
                          reg53 : reg78)}) : reg14[(5'h11):(5'h10)]) > (reg1447[(3'h7):(3'h5)] >= (~^$unsigned($unsigned(reg1469)))));
              reg1486 = ((reg10 * (~&reg66[(4'he):(4'h8)])) ?
                  reg1447 : $signed(reg1478[(3'h4):(1'h0)]));
              reg1487 <= $signed($signed($signed($unsigned(reg63[(5'h19):(1'h1)]))));
              reg1488 <= $unsigned(reg59[(2'h2):(1'h0)]);
            end
        end
      else
        begin
          if ((reg7 != reg1470[(5'h18):(2'h3)]))
            begin
              reg1467 = (reg67 ?
                  ((($signed(reg1459) ?
                          reg1459[(4'hb):(1'h0)] : reg1466[(4'h8):(2'h3)]) ?
                      reg49[(3'h4):(2'h3)] : $unsigned((reg1456 + reg75))) == $unsigned($unsigned({reg66}))) : $signed((-{$unsigned(reg1479)})));
              reg1468 = $signed(reg1488);
              reg1469 <= (($signed($signed($unsigned((8'hbe)))) & reg75[(1'h1):(1'h0)]) & (~|$unsigned((&(~&reg58)))));
              reg1471 <= reg62;
              reg1472 <= $unsigned(reg89[(3'h4):(1'h1)]);
            end
          else
            begin
              reg1467 = (-($signed(((^(7'h4b)) ?
                      $signed(reg1472) : $unsigned(reg1488))) ?
                  ({reg1475[(5'h16):(5'h10)]} ?
                      $unsigned((8'hba)) : $signed(((8'h9f) ?
                          wire1 : reg1467))) : reg1459));
              reg1469 <= ((((|((8'ha0) <<< (8'had))) ?
                          reg1465 : (~&$signed(reg56))) ?
                      reg67[(2'h3):(2'h2)] : {(reg1474[(5'h1c):(5'h16)] ?
                              reg1474 : $unsigned(reg1477)),
                          ($signed(reg89) ? (reg62 - reg28) : wire1446)}) ?
                  reg11 : (reg1465[(4'h8):(2'h2)] << reg20));
              reg1470 = ($unsigned((^~$unsigned($unsigned(reg1457)))) < (8'hb8));
              reg1471 <= ($unsigned(reg21[(1'h0):(1'h0)]) ?
                  {$unsigned(reg1456),
                      (~^(&(reg49 << (8'hb2)))),
                      $unsigned(((reg1459 == reg63) == reg1470[(4'ha):(3'h6)]))} : $unsigned((^$signed($unsigned(reg11)))));
              reg1472 <= ((~|reg1482[(2'h2):(1'h0)]) ?
                  $signed(((~^wire1446) <<< $unsigned($unsigned(reg1469)))) : (|{wire2[(3'h6):(3'h4)],
                      reg60,
                      (reg1478 ? reg1485 : (+reg66))}));
              reg1474 = (~|reg1473[(4'h8):(4'h8)]);
              reg1475 = reg79;
            end
          if ((reg1472 <<< $unsigned({reg5})))
            begin
              reg1478 = (^$unsigned((8'hb2)));
              reg1479 <= ((|($unsigned($unsigned(reg1483)) >> reg62)) ?
                  (~|$signed((!(~^reg5)))) : $signed((~$signed((8'hb2)))));
              reg1481 <= (wire1 ?
                  $signed(reg79) : ({((reg1472 + reg50) ?
                          wire1444 : (!reg11))} ^~ $unsigned(reg64[(3'h4):(1'h0)])));
              reg1482 <= reg62;
              reg1484 = ($unsigned((reg1487[(1'h0):(1'h0)] <<< ($unsigned(reg1483) | $signed((7'h4b))))) ^~ (|$unsigned({(~|reg1457),
                  reg1479})));
            end
          else
            begin
              reg1478 = $unsigned((^$unsigned(reg84[(2'h3):(2'h2)])));
            end
          for (forvar1485 = (1'h0); (forvar1485 < (1'h1)); forvar1485 = (forvar1485 + (1'h1)))
            begin
              reg1487 <= ($unsigned((reg64[(3'h5):(3'h5)] >> $signed((7'h49)))) != wire3[(3'h4):(1'h0)]);
              reg1489 = ((reg1482[(4'hd):(2'h3)] >> ($signed($unsigned(reg1465)) ?
                      ($unsigned(reg1479) ?
                          (|(8'ha8)) : $unsigned(reg64)) : {(reg1484 ?
                              reg40 : (8'hac)),
                          $unsigned(reg78)})) ?
                  $unsigned((|$signed($signed((8'ha8))))) : $unsigned($signed($signed({reg31}))));
              reg1490 = ({$unsigned($signed($unsigned((7'h58)))),
                  (&$unsigned(reg11[(5'h10):(2'h3)])),
                  (|{reg1482[(4'h8):(3'h7)],
                      $signed(reg1472)})} <= ({((reg49 >>> reg1483) ?
                          reg1479 : reg25)} ?
                  reg66 : reg20));
            end
          if (reg50[(4'he):(4'he)])
            begin
              reg1491 = $unsigned((($unsigned((reg1490 <= reg1484)) ?
                  $unsigned($unsigned(wire2)) : $unsigned((~^reg49))) - wire2));
              reg1492 <= reg66;
              reg1493 <= $unsigned({$unsigned({reg1469[(3'h5):(1'h1)]}),
                  reg46[(4'h9):(3'h5)],
                  (reg1488[(3'h7):(3'h6)] ^ (~|reg1477[(3'h6):(1'h1)]))});
              reg1494 = $signed({(((reg10 ?
                          (8'ha9) : reg1480) - reg59[(1'h0):(1'h0)]) ?
                      ((reg28 ^~ reg58) != (reg28 ?
                          reg49 : reg31)) : $signed($signed(reg1487))),
                  reg60,
                  reg86});
            end
          else
            begin
              reg1492 <= ((^~(reg1473[(2'h3):(2'h3)] ?
                  (+(!reg84)) : (8'h9e))) && ($signed(({reg28,
                  reg1475,
                  reg1465} >> (reg1474 ?
                  reg1466 : reg5))) ^ ($signed($signed((7'h43))) ?
                  (^(&reg1469)) : ($signed(reg1486) ?
                      (~&(7'h4c)) : {reg79, reg86}))));
              reg1493 <= wire1;
            end
          reg1495 <= reg1476;
          reg1496 <= (-($signed((~&reg53)) ?
              wire1 : $unsigned($signed({reg1487, reg56}))));
          reg1497 <= reg7[(4'hf):(4'h8)];
        end
      if ($unsigned((reg1488 ?
          $signed({(wire1 == reg75)}) : ($signed(reg1474[(5'h11):(4'h8)]) ?
              (!reg10[(4'hb):(1'h1)]) : forvar1472[(5'h10):(4'h9)]))))
        begin
          for (forvar1498 = (1'h0); (forvar1498 < (3'h4)); forvar1498 = (forvar1498 + (1'h1)))
            begin
              reg1499 = (({$signed($signed(reg11)),
                      reg1485[(3'h4):(1'h1)],
                      {reg1492}} ?
                  ((reg1457 & (+reg1492)) <= reg1492[(2'h2):(2'h2)]) : ((reg1474 & (reg11 ?
                      forvar1498 : reg25)) ^~ $signed((^reg1494)))) >> (reg43[(4'he):(1'h0)] ?
                  reg1457[(2'h2):(2'h2)] : $unsigned(reg1472)));
              reg1500 = (forvar1485[(2'h3):(2'h2)] ?
                  ((~|$signed(reg14[(5'h10):(2'h3)])) ~^ ((^~{reg58,
                      reg84}) * $signed((+reg1470)))) : $signed(reg1470[(4'hb):(2'h3)]));
              reg1501 = reg1482;
              reg1502 <= reg82[(2'h2):(1'h0)];
              reg1503 = (7'h40);
            end
          for (forvar1504 = (1'h0); (forvar1504 < (1'h0)); forvar1504 = (forvar1504 + (1'h1)))
            begin
              reg1505 <= ($unsigned((+(|(reg56 ? reg1453 : wire0)))) ?
                  (reg11[(4'hd):(3'h6)] ?
                      reg1475[(3'h5):(3'h5)] : $unsigned($signed((reg62 ?
                          reg64 : reg49)))) : reg1465[(5'h1b):(1'h1)]);
              reg1506 <= $unsigned((($unsigned(reg78) ~^ {(reg1493 << reg60)}) ?
                  ((-reg1500) ? reg1488 : reg1470[(5'h18):(4'ha)]) : ((reg1480 ?
                          $unsigned(reg81) : reg1503[(3'h5):(1'h0)]) ?
                      ($unsigned(reg10) ?
                          (reg1457 ? reg1475 : reg1497) : (reg27 ?
                              reg66 : reg1469)) : $signed(reg59[(2'h2):(1'h1)]))));
              reg1507 = reg1502;
              reg1508 = $signed($signed($unsigned((&reg1469[(3'h6):(1'h1)]))));
            end
          if (reg1481)
            begin
              reg1509 = (reg1469[(3'h5):(2'h2)] ?
                  reg1508[(2'h2):(2'h2)] : reg21[(4'hb):(4'h9)]);
              reg1510 <= ((reg1484[(4'hb):(3'h6)] ?
                  reg7 : ($signed((reg1501 >>> (8'ha6))) ^~ ((reg1478 | reg5) ?
                      (^~reg56) : ((7'h54) ? reg1474 : reg27)))) * ({({reg40,
                              reg53} ?
                          (7'h51) : reg84),
                      reg46} ?
                  ((~&reg59[(3'h6):(2'h3)]) ?
                      (~{reg1506, reg89, reg62}) : ((reg81 ?
                              reg1473 : reg1505) ?
                          $unsigned(reg1475) : forvar1504)) : $unsigned(reg46)));
              reg1511 = ((+$unsigned(((reg81 ? (8'hb1) : reg60) ?
                      {reg27} : ((8'ha1) ? reg1480 : reg1476)))) ?
                  (($unsigned((reg53 >> reg62)) != ((wire0 ?
                      reg1505 : (7'h4a)) << $signed(reg20))) + $unsigned({(!wire1446),
                      wire0[(5'h16):(3'h4)],
                      reg1457[(4'h9):(1'h1)]})) : (((~^(reg21 ?
                          wire3 : reg1481)) >> (reg27[(4'hf):(1'h0)] <<< reg1474)) ?
                      wire1[(5'h1a):(3'h6)] : {(reg1474[(4'h8):(3'h7)] + $signed(reg1459)),
                          ($unsigned(reg1478) ?
                              (forvar1484 ?
                                  reg57 : reg63) : (forvar1484 | reg75)),
                          reg79}));
              reg1512 = $unsigned($unsigned(reg1447[(4'ha):(3'h6)]));
            end
          else
            begin
              reg1510 <= reg1476;
              reg1511 = (|(((~|(~^(7'h54))) <<< ($signed((8'ha8)) ?
                      $unsigned(reg1489) : (~reg31))) ?
                  (-$signed(reg1478)) : (+reg1499)));
              reg1513 <= (reg11 ^~ $unsigned((reg1473 ?
                  $unsigned(wire2) : (!reg63))));
              reg1514 <= (~^$signed(({((8'hb8) ~^ reg1471)} ?
                  (~^$signed(reg1484)) : {(+reg78)})));
            end
          for (forvar1515 = (1'h0); (forvar1515 < (2'h2)); forvar1515 = (forvar1515 + (1'h1)))
            begin
              reg1516 <= {((7'h50) == reg1464)};
              reg1517 <= (({$unsigned(reg1479[(3'h4):(2'h3)])} ?
                      forvar1485[(3'h5):(1'h1)] : (reg75[(2'h2):(1'h0)] ~^ $unsigned((reg1451 ?
                          reg1491 : wire3)))) ?
                  reg28 : (+$signed(reg59[(3'h4):(3'h4)])));
              reg1518 = reg1494[(4'ha):(4'h8)];
              reg1519 <= (({$unsigned((reg50 ? reg1465 : (8'hbd)))} ?
                      $signed(reg57[(3'h6):(3'h4)]) : (((+reg1490) >> reg79[(3'h6):(2'h3)]) | reg1510[(5'h16):(5'h10)])) ?
                  ((+(reg64 ? $unsigned(reg31) : (reg1508 ~^ reg1506))) ?
                      (reg1512 * (+{reg78, wire3})) : reg1507) : reg50);
            end
          reg1520 <= ((reg1496 ? reg1451[(4'h8):(2'h2)] : $signed(reg60)) ?
              reg51 : ({{(reg1484 ?
                          reg1512 : reg1490)}} || $unsigned(($unsigned(reg1517) ~^ {reg1470}))));
          for (forvar1521 = (1'h0); (forvar1521 < (2'h3)); forvar1521 = (forvar1521 + (1'h1)))
            begin
              reg1522 = (reg1471[(2'h2):(1'h1)] && ((&$signed({forvar1472})) ?
                  $signed((reg40 ?
                      reg1480 : forvar1504[(5'h15):(2'h2)])) : (!$unsigned((reg75 ^ (8'h9f))))));
              reg1523 <= {((~&reg1457) <= $unsigned($unsigned($unsigned(reg21))))};
              reg1524 <= (reg1471 ~^ (8'h9d));
              reg1525 = $unsigned(((($signed(reg1470) >> $signed(reg1509)) ?
                      $unsigned(reg28) : (~^reg56[(1'h1):(1'h0)])) ?
                  ($signed((~reg1508)) != $signed((8'hb5))) : reg1519));
            end
        end
      else
        begin
          if (reg1471)
            begin
              reg1498 = $unsigned(reg1484[(4'hb):(3'h4)]);
              reg1502 <= (|(forvar1504[(4'h9):(3'h5)] - ($unsigned(reg1512) < (7'h4d))));
            end
          else
            begin
              reg1502 <= {{($unsigned({reg79, reg40}) || reg1502),
                      ((-forvar1484[(1'h1):(1'h0)]) && (reg86[(2'h2):(1'h0)] + reg1485)),
                      reg1469[(2'h2):(2'h2)]}};
              reg1503 = $signed((-(({reg1480, reg75, reg40} ?
                  (8'hb4) : (reg1494 & reg1487)) & $signed((^~reg46)))));
              reg1504 <= wire1446;
              reg1505 <= $signed($signed(reg89[(3'h6):(3'h4)]));
              reg1506 <= reg14;
            end
          reg1507 = $signed(((^~({reg20, reg1476} < ((7'h4c) ?
                  reg1484 : reg82))) ?
              $signed((~^reg59[(3'h5):(2'h3)])) : reg63[(5'h10):(3'h5)]));
          reg1510 <= reg1465;
          reg1511 = $signed((reg1487[(4'hc):(4'h8)] == $signed({$unsigned(reg1481),
              {reg43, reg1473, reg1498},
              reg60})));
          reg1513 <= reg1480;
          reg1515 = (|((+$unsigned($unsigned(reg1501))) ?
              (^~((~&reg1477) ?
                  (reg1516 ? wire0 : reg82) : reg56)) : $signed(reg1495)));
        end
      reg1526 = ($unsigned($unsigned(($signed(reg1451) >> $signed(reg1502)))) ?
          reg1471[(4'he):(1'h0)] : (reg1494[(4'hd):(2'h3)] ?
              ($unsigned($signed((8'ha1))) * {$signed(reg1481),
                  (reg1484 ? reg1482 : reg1494)}) : (~&{(reg46 != reg1447),
                  (reg21 ? reg1491 : forvar1484),
                  (reg27 ~^ reg1475)})));
      for (forvar1527 = (1'h0); (forvar1527 < (3'h5)); forvar1527 = (forvar1527 + (1'h1)))
        begin
          if (reg1495)
            begin
              reg1528 <= reg1484;
              reg1529 = {$unsigned({{$unsigned(reg89),
                          (~|reg84),
                          reg1525[(1'h0):(1'h0)]}}),
                  $signed($signed(reg1525))};
            end
          else
            begin
              reg1528 <= $unsigned({$unsigned((((8'hb0) ?
                      reg1465 : reg1459) ^~ $signed(forvar1527))),
                  $signed((reg14 & (+reg89))),
                  $unsigned(reg60[(5'h13):(3'h5)])});
              reg1529 = (($signed(({reg1503, (8'hb3)} ?
                      (reg79 == reg1526) : (^reg1528))) ?
                  $signed({$unsigned(reg60)}) : (reg1497[(1'h1):(1'h0)] ?
                      wire1446 : reg81[(3'h5):(1'h1)])) + (!(~^((|(7'h4f)) ?
                  wire0 : reg1464[(1'h0):(1'h0)]))));
              reg1530 <= $signed(((($signed(reg11) ?
                          (reg58 * reg1511) : reg63[(2'h2):(2'h2)]) ?
                      (+reg1447) : reg1508[(5'h11):(2'h3)]) ?
                  (($signed((8'haf)) << reg1493) && $unsigned((reg1494 ?
                      reg60 : reg1473))) : $unsigned((forvar1485[(3'h6):(3'h5)] ?
                      {reg56, reg1482, reg78} : (~^reg1526)))));
            end
          if ((((reg82 ?
                  reg1497[(3'h4):(1'h0)] : $signed((~&(7'h56)))) | $unsigned($unsigned((reg27 <= reg1469)))) ?
              ((reg1488[(4'hb):(3'h4)] ?
                      ((reg1484 & reg1519) ?
                          (~^reg1478) : (7'h44)) : reg1510[(5'h19):(2'h2)]) ?
                  (~{$unsigned(reg1477),
                      reg14,
                      forvar1527[(3'h4):(2'h3)]}) : (~|((reg1495 | reg86) ^ (reg1496 || reg7)))) : $unsigned({(&((7'h46) ?
                      (7'h4e) : reg1525)),
                  $unsigned((~|reg1516))})))
            begin
              reg1531 = $unsigned(reg49[(3'h4):(2'h2)]);
            end
          else
            begin
              reg1531 = {$unsigned(((^reg1484) ? reg78 : $unsigned({wire1})))};
              reg1532 <= reg1495;
              reg1533 <= {reg1482[(4'hc):(1'h1)]};
            end
        end
      if ({$signed(($signed((~^forvar1485)) << ((reg14 ?
              reg1507 : reg31) | (forvar1521 ? reg21 : reg1500))))})
        begin
          reg1534 = reg1481;
        end
      else
        begin
          reg1534 = reg1489[(3'h4):(1'h0)];
          reg1535 = $unsigned((8'hbc));
          if (reg40[(3'h5):(3'h5)])
            begin
              reg1536 <= ((^$signed({{reg1528, reg49, reg79}, (~&reg1475)})) ?
                  (((&$signed(reg51)) ?
                      (~^reg1535) : (+reg79)) != ($unsigned((~&(7'h4b))) ?
                      ((+(7'h4b)) ?
                          $unsigned(reg1513) : reg11[(5'h11):(3'h6)]) : (~^$signed(reg79)))) : (reg1495[(3'h6):(3'h5)] ?
                      ($unsigned({reg1465, reg38}) ?
                          ($unsigned(reg1492) * $unsigned(reg10)) : reg1499[(1'h0):(1'h0)]) : ((+$signed(reg1486)) ?
                          reg1477[(3'h7):(3'h7)] : $signed((!reg1492)))));
              reg1537 = ({(((reg1457 ? reg1532 : reg1475) << (+reg1535)) ?
                          (~&((7'h49) ?
                              reg1533 : reg86)) : wire3[(4'hc):(3'h5)])} ?
                  reg1511 : (({{forvar1521, (8'hac)}} >> {$signed((8'hae)),
                      reg1506,
                      {reg1507,
                          (7'h4f)}}) << (~^((+reg82) >>> $signed(reg1479)))));
              reg1538 = (reg1507 ? $unsigned(forvar1504) : reg51);
              reg1539 = $unsigned(reg58);
              reg1540 = reg1499[(2'h2):(1'h1)];
            end
          else
            begin
              reg1537 = $signed((!reg64[(1'h0):(1'h0)]));
              reg1541 <= reg1506[(2'h2):(1'h0)];
              reg1542 = reg1475;
              reg1543 = $unsigned(reg1491[(4'hf):(1'h1)]);
              reg1544 <= {((-(~^forvar1485[(5'h14):(2'h2)])) >= ((~|reg1512[(4'hc):(4'ha)]) ?
                      $signed((-reg1459)) : $unsigned(reg28))),
                  $unsigned((^$signed((7'h54)))),
                  {$signed((!{wire2, reg86}))}};
              reg1545 <= (8'ha5);
            end
          if (reg1465[(5'h12):(4'h9)])
            begin
              reg1546 = reg28;
              reg1547 <= $unsigned((|$unsigned($signed(((8'h9f) ?
                  (7'h57) : reg1518)))));
              reg1548 = reg21[(5'h11):(1'h1)];
              reg1549 <= {{reg1484[(4'hb):(1'h0)]},
                  (+$signed((7'h46))),
                  ($signed($unsigned(reg1514)) >> ($unsigned(reg1494) ?
                      ((~&reg1516) == ((8'haa) ?
                          reg1526 : reg1514)) : (reg67[(4'hb):(3'h7)] ?
                          reg1533 : $signed(reg1503))))};
            end
          else
            begin
              reg1547 <= $signed((!$signed(reg1457)));
            end
        end
      reg1550 <= ($signed(reg1519[(5'h17):(4'ha)]) == $signed({(reg28[(1'h1):(1'h1)] ?
              (~&reg1480) : $signed((8'h9c)))}));
    end
  always
    @(posedge clk) begin
      if (reg1506)
        begin
          reg1551 <= reg79[(3'h5):(3'h4)];
          if (($unsigned((^(&$unsigned(reg7)))) >= $unsigned((($signed(reg1456) ~^ (~|reg78)) >= (~reg59)))))
            begin
              reg1552 <= (-reg59);
              reg1553 <= {$unsigned(reg20),
                  (8'ha7),
                  $unsigned($unsigned(($signed(reg53) >= $signed(reg40))))};
              reg1554 = {reg1553[(2'h3):(2'h3)],
                  reg1506[(2'h2):(1'h0)],
                  (reg1492 ?
                      ((^{reg1466, reg1523}) ?
                          reg1551[(3'h5):(1'h0)] : wire1444) : {reg1492[(1'h1):(1'h0)],
                          reg1530,
                          {reg56[(1'h1):(1'h0)], reg5[(4'h8):(3'h6)]}})};
              reg1555 <= {reg1483};
              reg1556 <= (^(~|(8'hbc)));
              reg1557 = $signed(($unsigned((-(reg1520 != reg40))) ?
                  {(reg1519 >= $signed(reg27)),
                      ((reg49 ? reg1555 : reg27) ?
                          $signed(reg1483) : (7'h48))} : reg62));
              reg1558 = ($unsigned(reg1533) & (|{reg1466}));
            end
          else
            begin
              reg1554 = (reg1558 ? reg1520 : reg50);
              reg1555 <= $signed({(-$unsigned($signed(reg1483)))});
              reg1556 <= wire1[(4'h8):(3'h7)];
              reg1557 = (^~(^~(+(~|$unsigned(reg53)))));
              reg1559 <= reg1533[(3'h5):(1'h0)];
              reg1560 <= reg59;
            end
        end
      else
        begin
          if (((+$signed($unsigned({(8'hb2), reg1464}))) ?
              ((^$unsigned((reg59 ? reg1555 : reg1451))) ?
                  $unsigned($signed(reg1516[(5'h13):(3'h4)])) : $unsigned($unsigned((reg1451 ~^ (7'h55))))) : (7'h56)))
            begin
              reg1554 = ((reg43 ?
                      (~|{$signed(reg1541)}) : {((-(8'hac)) ?
                              $signed(reg1469) : ((8'hb8) && reg1453)),
                          ($signed(reg1495) ? (&reg1456) : (^reg10))}) ?
                  {reg1459,
                      $unsigned(reg1514),
                      $unsigned((^(^~reg60)))} : reg1477[(3'h6):(1'h0)]);
              reg1557 = (~^$unsigned($unsigned($unsigned(reg1560[(4'he):(4'hb)]))));
              reg1558 = (reg57[(4'h9):(3'h6)] <= ((7'h50) + (~&((7'h4b) == (reg1502 ?
                  reg67 : reg1536)))));
            end
          else
            begin
              reg1554 = ((^$unsigned($unsigned((reg1544 ?
                      reg1555 : reg1488)))) ?
                  $signed(reg81) : reg1528[(2'h2):(2'h2)]);
              reg1557 = $signed($signed(($unsigned($signed(reg1516)) ?
                  (+$signed(reg1481)) : ((reg62 ?
                      (8'h9e) : reg10) ^ reg1519[(5'h14):(2'h2)]))));
              reg1558 = (($unsigned(reg1451[(2'h3):(1'h1)]) ~^ reg21[(4'h9):(3'h5)]) ?
                  $unsigned($signed(reg1465)) : (reg1466 + ((|(reg1488 ?
                          reg79 : reg43)) ?
                      reg43[(1'h1):(1'h1)] : $unsigned(reg1547[(3'h4):(1'h1)]))));
              reg1559 <= reg1524[(5'h15):(2'h2)];
              reg1560 <= $unsigned($signed({(8'ha1),
                  $unsigned((~reg28)),
                  (reg1506 >>> reg75[(1'h1):(1'h1)])}));
              reg1561 <= reg1487;
              reg1562 = reg60;
            end
          reg1563 <= ((reg27[(5'h15):(4'hb)] ^~ reg1530[(2'h2):(1'h0)]) ?
              reg78 : ($unsigned((reg14[(1'h0):(1'h0)] ?
                      (reg84 >> reg1557) : ((8'ha2) & reg1547))) ?
                  (~&(!(8'haf))) : ((|$unsigned(reg1493)) || ((reg89 ^~ reg1545) | reg1514))));
          reg1564 = $unsigned({reg1451[(4'hb):(2'h3)], reg1544});
          for (forvar1565 = (1'h0); (forvar1565 < (1'h0)); forvar1565 = (forvar1565 + (1'h1)))
            begin
              reg1566 <= (($unsigned(reg1544[(3'h5):(1'h1)]) ?
                      reg1557[(5'h10):(4'hd)] : ($signed((reg1476 | (7'h48))) + (~|(~^reg1487)))) ?
                  $unsigned((~&wire0[(5'h12):(5'h12)])) : $unsigned((reg89[(5'h16):(4'h8)] == ((reg1492 ?
                      (7'h49) : (7'h44)) <<< $signed(reg50)))));
              reg1567 <= ((-$signed((8'ha2))) ?
                  ((8'ha4) ?
                      (&($signed(reg79) >= (wire1444 ?
                          reg1562 : wire1))) : reg1502) : (wire1444[(3'h6):(2'h2)] ?
                      $signed(reg1497) : (!(~&$unsigned(reg1564)))));
              reg1568 <= reg1481[(5'h1a):(5'h10)];
              reg1569 = ($signed($unsigned((7'h47))) <= (^($signed($signed(reg1476)) != (reg14 <= reg1488))));
            end
        end
      reg1570 = (~&($unsigned($unsigned(reg1555)) ?
          ((reg1466[(3'h4):(1'h0)] ?
              $unsigned(reg1567) : (reg1466 ?
                  (8'hb9) : (7'h46))) == $unsigned((8'had))) : $signed(reg1528[(2'h3):(1'h1)])));
      for (forvar1571 = (1'h0); (forvar1571 < (2'h2)); forvar1571 = (forvar1571 + (1'h1)))
        begin
          for (forvar1572 = (1'h0); (forvar1572 < (2'h2)); forvar1572 = (forvar1572 + (1'h1)))
            begin
              reg1573 = reg1560[(4'hd):(4'h8)];
              reg1574 <= $unsigned($unsigned((reg1504[(4'hd):(3'h4)] ?
                  reg1456[(3'h5):(1'h0)] : reg1559[(4'hc):(2'h3)])));
              reg1575 <= reg62[(3'h6):(2'h2)];
            end
        end
    end
  assign wire1576 = $signed(reg27);
  assign wire1577 = $signed($unsigned($unsigned(reg1568)));
  always
    @(posedge clk) begin
      reg1578 = reg63;
      reg1579 = reg1466;
      reg1580 = $unsigned($unsigned(($unsigned($unsigned((7'h4a))) << ({reg1519,
          reg1487} || (~^reg79)))));
      if ($signed($unsigned(($unsigned((reg1550 ?
          reg1513 : reg1516)) >>> ({reg1541, reg66} == (wire0 ^~ reg1523))))))
        begin
          if ($unsigned((!(($signed((7'h50)) ? (reg1549 ^ (8'h9c)) : wire2) ?
              reg1520 : (8'haa)))))
            begin
              reg1581 <= $unsigned($unsigned(($unsigned((reg1513 ?
                  reg1567 : reg1506)) ^ reg57)));
              reg1582 = (&reg58[(1'h0):(1'h0)]);
              reg1583 <= ($signed((reg67[(4'ha):(4'h8)] <<< reg1510)) - $signed(reg20[(4'he):(4'ha)]));
              reg1584 = wire1[(3'h7):(3'h7)];
              reg1585 <= (8'hb3);
              reg1586 = ($unsigned($signed((|$unsigned(wire1)))) ?
                  $signed((7'h46)) : {((~&(-reg1497)) ?
                          reg57[(4'hc):(3'h6)] : (~&(reg1550 ?
                              (7'h45) : reg1551)))});
              reg1587 = $signed($signed({$signed((+(8'ha9))),
                  {(7'h4e), $signed((8'ha6)), reg1493},
                  ($signed(reg1545) << $signed(reg1520))}));
            end
          else
            begin
              reg1581 <= reg1504;
              reg1583 <= (^~reg1504[(1'h0):(1'h0)]);
              reg1585 <= ($signed(reg50[(5'h11):(4'ha)]) ?
                  ({reg1582[(2'h2):(1'h0)],
                          ((~(8'hbf)) ?
                              {reg1578, wire3, (8'hb8)} : (reg1510 << reg79))} ?
                      reg1523 : reg5) : (({$signed((8'hbf)),
                              (reg1513 <= reg31),
                              reg1456} ?
                          ((~reg1497) - ((7'h54) != reg1559)) : ((reg25 ?
                              reg1520 : (7'h4b)) ~^ (!reg1559))) ?
                      ($signed($signed((8'had))) << ({reg84, reg1566} ?
                          reg1580[(3'h5):(3'h5)] : (reg1496 | reg1575))) : $unsigned((7'h42))));
            end
          reg1588 = {reg49[(3'h6):(2'h3)],
              ((&((&reg1453) ? (!(7'h4c)) : reg1568)) ~^ (~^{$signed((8'hb5)),
                  $unsigned(reg1506)})),
              $unsigned($signed($signed(reg1549)))};
        end
      else
        begin
          reg1581 <= $unsigned({(8'hb0), reg1513});
          for (forvar1582 = (1'h0); (forvar1582 < (2'h2)); forvar1582 = (forvar1582 + (1'h1)))
            begin
              reg1584 = ((((&reg1492) > reg40[(4'he):(4'h9)]) ?
                  (reg1556 ?
                      (reg46[(3'h4):(1'h0)] >> reg20) : $signed($signed((8'ha7)))) : {($signed(reg49) >> (!reg25)),
                      {((7'h4d) > (7'h44)), (reg1574 >>> (8'hac))}}) * reg1549);
              reg1586 = {{wire1576, (|reg1516), (reg79 - reg64)},
                  (+(reg1530 ?
                      reg1583 : {reg53, (reg1514 ? wire1446 : (8'hbc))})),
                  reg43};
              reg1587 = (7'h40);
              reg1589 <= $signed($unsigned(reg1553));
              reg1590 = $unsigned($unsigned(reg1553));
              reg1591 = (~&$signed((reg5[(3'h7):(3'h5)] ?
                  (-$signed(reg1493)) : $signed(reg1590[(1'h1):(1'h1)]))));
              reg1592 = $signed((wire1576[(2'h2):(1'h1)] >>> (((reg50 > (8'hb5)) << reg86[(3'h7):(3'h6)]) ?
                  ({reg1587} || $signed(reg1563)) : ((reg1545 >>> reg1544) ?
                      (reg62 == reg11) : $signed((8'had))))));
            end
          reg1593 <= $unsigned($signed(reg78[(1'h0):(1'h0)]));
          if ((-(((((8'h9e) <<< reg21) - (reg1520 ?
                  wire1576 : reg11)) + (-(reg1533 ? wire1577 : (7'h4e)))) ?
              (wire1[(5'h1e):(5'h19)] | $unsigned($unsigned(reg1516))) : $unsigned(reg1506))))
            begin
              reg1594 <= reg21[(3'h5):(3'h5)];
            end
          else
            begin
              reg1595 = (^~reg1536);
              reg1596 <= (wire3[(1'h1):(1'h0)] <<< {(reg1556[(2'h2):(1'h0)] ?
                      (~$unsigned((8'hba))) : ($signed((7'h4f)) ?
                          reg1582[(3'h6):(2'h2)] : reg1551))});
              reg1597 = (+reg1520);
              reg1598 = (($unsigned(((reg1483 ? reg79 : reg1575) ?
                      $unsigned(reg1496) : reg1585)) ?
                  (&reg1466[(2'h3):(2'h2)]) : $signed($unsigned($signed(wire0)))) && reg1556[(5'h13):(4'h8)]);
              reg1599 = $unsigned($signed((reg1556 + $unsigned((~reg1457)))));
              reg1600 <= (8'hb6);
              reg1601 <= (({reg43,
                      (~(^~reg81)),
                      $unsigned($unsigned(reg1497))} && {wire1446[(2'h3):(1'h1)],
                      ({reg27} == reg1497[(4'h9):(3'h4)])}) ?
                  ($signed((reg1592[(2'h2):(1'h1)] ?
                          (reg1600 ? reg1536 : reg1559) : $unsigned(reg59))) ?
                      {($signed(reg1599) ?
                              $signed(reg1587) : {reg25, reg1591, reg1582}),
                          (reg1547 ?
                              $unsigned(reg1582) : (&(7'h45)))} : $signed($unsigned(reg86[(1'h0):(1'h0)]))) : (^(((+reg1451) != reg1591[(4'hd):(4'ha)]) ?
                      $unsigned($signed(reg1597)) : reg1457)));
            end
          reg1602 <= $signed(wire2);
          for (forvar1603 = (1'h0); (forvar1603 < (3'h4)); forvar1603 = (forvar1603 + (1'h1)))
            begin
              reg1604 <= $unsigned((&(($unsigned(reg1583) | (reg1520 ^ reg75)) || $unsigned({reg1588}))));
            end
          for (forvar1605 = (1'h0); (forvar1605 < (3'h5)); forvar1605 = (forvar1605 + (1'h1)))
            begin
              reg1606 = (~|(8'hb6));
              reg1607 = ($signed(reg1563) ?
                  $unsigned((+({reg25, reg1457, reg1523} ?
                      (~&reg14) : reg1479[(4'h9):(1'h0)]))) : (|reg1496));
              reg1608 = (~(($signed((8'ha4)) > $unsigned((reg1456 ?
                      reg75 : reg1590))) ?
                  (reg1594[(5'h11):(4'ha)] ?
                      reg1604 : reg1549) : ((reg14[(5'h13):(3'h7)] + $unsigned(reg1513)) ?
                      $signed((^~reg40)) : $signed(reg1536[(3'h7):(3'h7)]))));
              reg1609 = (|(reg1556[(2'h3):(2'h3)] || {{forvar1605,
                      $signed(reg1584),
                      $unsigned(reg27)}}));
              reg1610 = (!reg1550);
              reg1611 <= (reg1465[(5'h13):(4'hd)] != ((reg57[(3'h5):(3'h4)] ^~ {((8'had) ?
                          reg1541 : reg1579)}) ?
                  (reg1530 <= $signed((&reg11))) : reg1602));
            end
        end
      if ($unsigned($signed((7'h54))))
        begin
          reg1612 = $unsigned((&($signed($signed(wire1444)) ?
              reg1556[(4'h9):(3'h4)] : $signed({reg1477, (8'ha8), reg31}))));
        end
      else
        begin
          if (reg1582[(4'hd):(4'hd)])
            begin
              reg1612 = ((^reg1602) ?
                  ((reg1587[(3'h6):(3'h5)] ?
                          ((|reg1602) < $signed(reg1611)) : (8'h9d)) ?
                      ($signed(reg1609[(3'h5):(1'h0)]) >= {$unsigned(reg1533),
                          {reg1523,
                              reg1547}}) : $unsigned({(reg1493 & forvar1605)})) : (~$unsigned($unsigned($unsigned(reg1578)))));
              reg1613 <= reg1496;
              reg1614 <= ((($unsigned((^~reg1466)) ?
                      $signed(reg1481[(4'h8):(3'h6)]) : ((-wire1446) ?
                          reg62 : (reg1532 * reg53))) ?
                  ($unsigned(reg1597[(2'h3):(1'h1)]) <<< reg1544[(4'h8):(2'h3)]) : $unsigned(reg1451[(5'h15):(3'h6)])) != $signed({reg1598[(3'h5):(3'h5)]}));
              reg1615 <= reg1482[(4'hc):(2'h3)];
              reg1616 = (!(((reg1523[(5'h10):(3'h5)] == reg1541[(1'h0):(1'h0)]) ?
                  reg1520[(5'h1c):(5'h1b)] : ((reg89 ?
                      reg1583 : reg1594) < (reg7 >= reg1615))) ~^ {(!(reg1549 ?
                      (8'haf) : reg1482))}));
            end
          else
            begin
              reg1613 <= (((~&{$unsigned(wire3), $unsigned(reg1602)}) ?
                      (((reg1544 ?
                          wire1444 : reg1607) - reg1579[(1'h0):(1'h0)]) * $unsigned((reg50 & reg66))) : ((reg62 ?
                          (~|reg50) : (reg1477 & reg1581)) || ({reg1465,
                              reg1600,
                              reg82} ?
                          (reg1544 ?
                              reg1590 : reg1582) : reg1559[(5'h10):(1'h1)]))) ?
                  reg1602 : (reg21[(3'h6):(2'h3)] ~^ ($signed($unsigned((8'hb1))) ?
                      ({reg63} ?
                          $unsigned(reg1608) : (8'ha9)) : ((reg1532 <<< reg1517) >= ((8'hac) >>> reg1532)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg1617 <= (|$unsigned((((~(8'h9c)) << $unsigned(reg53)) ?
          ((reg1585 * reg1459) ~^ {(7'h47),
              reg1497,
              reg1514}) : reg1456[(1'h0):(1'h0)])));
      for (forvar1618 = (1'h0); (forvar1618 < (2'h3)); forvar1618 = (forvar1618 + (1'h1)))
        begin
          for (forvar1619 = (1'h0); (forvar1619 < (3'h4)); forvar1619 = (forvar1619 + (1'h1)))
            begin
              reg1620 <= (~(-(7'h40)));
              reg1621 = reg1552;
            end
          reg1622 = ((&reg57) ?
              (-{$signed($unsigned(reg1602)),
                  {(reg1472 < reg1510)},
                  reg1581[(1'h1):(1'h0)]}) : (reg1585[(4'h8):(1'h1)] ?
                  ($signed($signed(reg1532)) ^~ (|reg1589)) : $signed(((reg1465 || reg14) ~^ (reg1553 * reg1556)))));
          reg1623 = (~$signed(reg53));
          for (forvar1624 = (1'h0); (forvar1624 < (3'h4)); forvar1624 = (forvar1624 + (1'h1)))
            begin
              reg1625 = reg1514;
              reg1626 = ((reg1456 ?
                      (($unsigned(reg1560) <<< $unsigned(reg1550)) ?
                          (-reg62[(1'h0):(1'h0)]) : reg1516[(4'hf):(3'h4)]) : (((reg1545 ?
                              reg86 : reg1560) ?
                          $unsigned(reg1566) : (~reg1466)) || (~&$signed(reg1533)))) ?
                  $signed(reg1476[(4'hc):(4'hc)]) : $signed($signed(((reg1451 ?
                      reg1620 : (7'h4e)) == ((8'hb3) ? (8'h9c) : reg1502)))));
              reg1627 <= {{(reg46[(2'h3):(2'h3)] <= ($unsigned(reg82) ?
                          $unsigned((8'hab)) : ((7'h4c) <<< reg1620))),
                      (8'hb4),
                      (7'h54)},
                  reg60[(5'h13):(3'h4)],
                  $signed(reg43[(3'h4):(1'h0)])};
              reg1628 = reg1617[(4'hc):(3'h6)];
              reg1629 <= $signed(((8'hae) | $signed($signed(reg1487[(4'h8):(4'h8)]))));
              reg1630 = ($unsigned(($signed(reg1492[(1'h0):(1'h0)]) == $signed($signed(reg43)))) ?
                  $unsigned(reg1544[(5'h14):(3'h7)]) : (reg1519 ?
                      reg40[(5'h14):(5'h14)] : $unsigned($signed((reg1472 ?
                          forvar1618 : reg1514)))));
            end
          for (forvar1631 = (1'h0); (forvar1631 < (3'h6)); forvar1631 = (forvar1631 + (1'h1)))
            begin
              reg1632 <= (reg10[(1'h0):(1'h0)] | $unsigned($unsigned((|{reg1623}))));
            end
          for (forvar1633 = (1'h0); (forvar1633 < (2'h3)); forvar1633 = (forvar1633 + (1'h1)))
            begin
              reg1634 = ($unsigned(reg1520[(3'h4):(2'h3)]) > reg1517);
              reg1635 = (reg1553 ? reg1627 : $signed((+reg1630)));
              reg1636 <= $signed(($unsigned(($signed((8'ha3)) >= $unsigned(reg1479))) ?
                  (-$signed({reg1623, reg86})) : reg43[(4'h8):(3'h4)]));
              reg1637 = (~reg1636);
              reg1638 <= (!$unsigned((reg1473[(2'h2):(1'h1)] ?
                  $unsigned((reg79 >>> reg1636)) : (|{reg67,
                      (8'h9c),
                      reg11}))));
              reg1639 <= {reg1482[(2'h2):(1'h0)]};
            end
          if (reg1524[(4'hc):(3'h5)])
            begin
              reg1640 = ($signed(reg53) ? reg75 : reg51[(4'hb):(4'hb)]);
              reg1641 = $unsigned((reg1465 | $unsigned((&$unsigned((7'h4c))))));
              reg1642 <= ((((-(reg1516 >= reg62)) << (reg1583 ?
                          (~&reg1453) : $unsigned(reg1635))) ?
                      reg1629 : (&{$signed(reg1524),
                          $unsigned(reg56),
                          $signed(reg1504)})) ?
                  $signed($unsigned((-reg1510[(5'h13):(1'h0)]))) : $signed(reg1634[(2'h2):(1'h1)]));
              reg1643 = ((~^(^((reg1629 ? reg1561 : reg1502) ^ {reg1481}))) ?
                  (($unsigned({reg1472}) >= $signed({(8'haf),
                      (8'hb9),
                      reg1551})) == $unsigned((reg67 >>> $unsigned(reg1611)))) : (8'ha6));
            end
          else
            begin
              reg1642 <= reg1473;
              reg1643 = $signed((~&(^~reg1622[(2'h2):(1'h0)])));
              reg1644 = (((reg1536 >>> $unsigned(reg1626[(2'h2):(2'h2)])) - reg1517[(3'h5):(1'h1)]) ?
                  reg27 : (reg1628[(1'h1):(1'h1)] ?
                      $signed((~&$unsigned(reg50))) : $unsigned((~&(reg1506 ?
                          reg1528 : wire1576)))));
              reg1645 = $signed(((^~(^~$unsigned((7'h51)))) != $signed($signed(reg1568[(3'h7):(2'h2)]))));
              reg1646 = ((7'h44) <<< $unsigned($signed((~^reg20))));
              reg1647 <= (&((~|reg1476) == (~|{(~reg1567)})));
            end
        end
      if (reg89[(4'ha):(1'h1)])
        begin
          reg1648 <= {(~reg1504), reg1641[(5'h17):(3'h5)]};
          reg1649 = ($unsigned($signed($signed(reg10))) ?
              (7'h56) : (|$unsigned((^(~|reg1481)))));
          reg1650 = $signed((reg78 ? reg57 : reg1472[(3'h4):(2'h3)]));
          reg1651 <= (($unsigned($signed(reg1647[(4'hd):(4'ha)])) ?
                  reg1561 : (&reg1549)) ?
              (^~((^~reg1541[(4'hb):(4'h8)]) ?
                  ((reg60 ? reg1476 : reg84) << (reg1640 ?
                      (8'ha5) : reg89)) : ((forvar1631 ?
                      reg1520 : reg1447) <= (!reg86)))) : reg1627);
          reg1652 = ($unsigned((~($signed(reg78) & reg1496[(4'h9):(2'h3)]))) * reg1594);
          if (reg1568)
            begin
              reg1653 = (7'h56);
              reg1654 = $signed(reg1602[(3'h7):(1'h0)]);
              reg1655 = ({$signed(({reg1482, reg1632} >= (8'ha2))),
                  (((reg1477 ?
                      reg1466 : reg1623) || (-reg20)) >> (~$unsigned(reg1620)))} << (~((~{reg1504,
                      (8'hb4)}) ?
                  $signed((reg43 ? reg53 : reg1583)) : $signed((reg1550 ?
                      reg1471 : (8'ha6))))));
              reg1656 = ((~^$signed(reg1601[(3'h5):(2'h2)])) == {(reg1567 == reg38)});
              reg1657 = $unsigned(($unsigned(($unsigned(reg1555) << $unsigned(reg1651))) & ((((8'hb6) ?
                          reg1514 : (8'h9d)) ?
                      $signed(reg1532) : $signed(reg1504)) ?
                  reg1637[(2'h3):(2'h2)] : (reg1530[(4'h9):(4'h8)] ?
                      reg1649[(4'h8):(3'h4)] : (^reg1634)))));
            end
          else
            begin
              reg1658 <= (~&reg5);
              reg1659 = forvar1633;
              reg1660 = reg43[(5'h12):(3'h4)];
            end
          if (reg1496[(3'h4):(2'h3)])
            begin
              reg1661 <= reg57[(4'hb):(1'h0)];
              reg1662 = $signed({({{reg1658},
                      reg5[(3'h7):(3'h4)]} < $signed($signed(reg27)))});
              reg1663 <= (reg10[(4'h9):(3'h6)] ?
                  (wire3 ~^ $unsigned(($unsigned(reg1659) < $signed(reg43)))) : ((~{(~|reg21),
                          reg27[(5'h13):(4'ha)]}) ?
                      {reg1519[(3'h5):(2'h2)],
                          $unsigned((reg1472 < forvar1618)),
                          reg59} : ($unsigned(reg1623[(1'h1):(1'h0)]) < reg1495)));
            end
          else
            begin
              reg1662 = reg1640[(4'hd):(4'h8)];
              reg1663 <= ($signed((^$signed({reg1649,
                  (8'hb2)}))) + (~|$unsigned(($unsigned(reg1634) ^ reg1451))));
              reg1664 <= reg57[(3'h5):(1'h0)];
              reg1665 <= ((reg1632[(3'h7):(2'h2)] ?
                      (^$signed((reg1545 ? reg1664 : reg1502))) : reg1581) ?
                  ($signed(($signed(reg1556) ?
                      (reg1530 + reg1566) : $signed(reg1643))) >>> {$signed(reg1495),
                      $unsigned(reg1553),
                      ($unsigned(reg1620) != (reg1544 != reg40))}) : $unsigned($unsigned($unsigned((^reg1487)))));
              reg1666 <= (~&$signed((($unsigned((8'ha7)) <<< (reg1471 < reg1602)) ?
                  $unsigned({reg1639, reg53, reg1658}) : {((7'h52) >>> reg58),
                      $signed(reg1640)})));
              reg1667 = (~&(^~(+{reg86[(3'h4):(2'h3)],
                  (reg1510 << (7'h45)),
                  $unsigned(reg1487)})));
              reg1668 <= (~|$unsigned((($unsigned(reg1464) ?
                  $unsigned(reg1492) : ((7'h50) ?
                      reg57 : reg1634)) ^ (8'hb8))));
            end
        end
      else
        begin
          reg1648 <= (reg1658 != $signed((7'h55)));
          if ({(wire3 ?
                  {(reg1506 << reg5),
                      (8'hac),
                      {$signed((8'hab)),
                          ((7'h41) ? reg1666 : wire0),
                          (!reg1466)}} : (({reg1545,
                      wire1444} * (reg1514 || reg1466)) & $unsigned((8'hb6)))),
              ({$signed((reg89 & forvar1633))} ~^ ((reg1551 <= (reg1594 ?
                  reg53 : reg66)) != $unsigned(forvar1624[(3'h7):(2'h2)])))})
            begin
              reg1651 <= $unsigned((~&($unsigned(((8'hbe) >= reg1532)) ?
                  $unsigned((reg1510 ? reg1488 : reg40)) : {reg1596})));
              reg1658 <= $signed($unsigned(reg89[(2'h2):(1'h0)]));
              reg1661 <= reg1666[(2'h2):(1'h0)];
              reg1662 = (^({{(reg1506 & reg1583),
                          (reg5 ~^ reg1488),
                          $signed(reg1567)},
                      reg1600[(4'hd):(1'h0)],
                      reg1459[(1'h1):(1'h0)]} ?
                  (~|(7'h40)) : (reg1488[(4'h9):(1'h0)] ?
                      (~|reg1622[(5'h13):(4'h8)]) : (~&$unsigned(reg21)))));
            end
          else
            begin
              reg1651 <= ((8'h9c) ? (-reg1523) : reg1620[(5'h10):(4'h9)]);
              reg1658 <= $unsigned($unsigned((reg1611[(3'h4):(3'h4)] | reg1502[(3'h7):(2'h2)])));
              reg1661 <= reg1652;
            end
          reg1663 <= (7'h50);
          for (forvar1664 = (1'h0); (forvar1664 < (3'h4)); forvar1664 = (forvar1664 + (1'h1)))
            begin
              reg1667 = reg1666;
              reg1669 = (~&(^$signed(((reg1465 > reg1541) ?
                  reg1630[(2'h3):(1'h1)] : reg1549[(5'h19):(5'h18)]))));
              reg1670 = (+(^(reg43[(4'he):(4'hb)] ?
                  $signed(reg1481) : reg1560)));
              reg1671 = (~&wire2[(4'hf):(4'hf)]);
              reg1672 <= ((~&(reg59[(2'h2):(2'h2)] | reg49[(3'h5):(2'h2)])) ~^ $signed((($signed(reg1541) << $signed(reg53)) ?
                  wire1444[(5'h14):(4'h8)] : reg1600)));
              reg1673 = ((8'hae) ? {(7'h4b)} : (reg59 ? reg67 : reg1550));
            end
          if ($unsigned(((({reg1566, reg1613} ?
              $unsigned(reg1641) : $signed(reg1645)) ~^ $signed((reg1459 ?
              (8'hbc) : reg1664))) != reg1551)))
            begin
              reg1674 <= $unsigned(($unsigned(({reg67} - $signed((8'ha2)))) ?
                  $unsigned((^~$unsigned(reg1563))) : $unsigned((((7'h4e) * reg1505) >> {reg1545,
                      reg1669}))));
              reg1675 = (+((reg1628 ? reg1574 : (+{reg1566})) ?
                  ($signed($signed(reg1669)) >= $signed((forvar1619 | reg50))) : ($unsigned(reg75) < (8'haf))));
            end
          else
            begin
              reg1674 <= $unsigned(reg49);
              reg1676 <= ((reg49[(3'h4):(2'h3)] == (((reg1667 & reg1465) ?
                      $signed(reg1464) : forvar1633[(4'h8):(3'h4)]) ?
                  reg1530 : {$signed(reg1472)})) <= $unsigned(({reg1456} << {$signed(reg81)})));
              reg1677 <= reg1642;
              reg1678 <= {{$signed((^$signed(reg1629)))}};
              reg1679 <= reg1472;
            end
          if (reg1647)
            begin
              reg1680 = reg46[(2'h3):(2'h3)];
              reg1681 <= reg1552;
              reg1682 = reg78;
              reg1683 = ((&(($unsigned(reg1620) ?
                      (reg1544 ^~ (8'ha9)) : $signed(reg1532)) << {(reg81 ?
                          reg1479 : (7'h45))})) ?
                  reg1497 : ($unsigned($unsigned($unsigned(reg43))) >> $signed((7'h57))));
              reg1684 <= ($unsigned(((&reg1650[(3'h7):(3'h6)]) ?
                      reg1552[(5'h12):(4'h9)] : reg1636[(4'he):(4'hd)])) ?
                  reg1647 : (7'h51));
            end
          else
            begin
              reg1680 = (reg1497 ?
                  $signed(forvar1631) : {$unsigned((&(&reg1504))), reg1589});
              reg1681 <= (~&($unsigned(reg7[(2'h2):(2'h2)]) ?
                  ((reg27 ? $unsigned((8'ha1)) : (reg1497 >= reg1635)) ?
                      (((8'hb7) ? reg1611 : reg46) ?
                          $signed(reg1614) : (reg1447 ?
                              reg86 : reg1510)) : ((7'h41) & ((8'hbc) + reg1651))) : $unsigned(((reg1683 <= reg1497) ?
                      (7'h56) : (-reg1514)))));
              reg1682 = ((($unsigned($unsigned((8'hba))) ?
                      $signed((reg1672 && reg1496)) : {(reg1671 ?
                              reg28 : reg1662),
                          (reg1502 ? reg64 : reg1645),
                          reg1594}) ?
                  $signed(reg57[(4'h9):(2'h3)]) : {((!reg1621) - (7'h4b)),
                      (!(8'hbf))}) || reg31[(4'ha):(2'h3)]);
              reg1683 = {{reg27}};
              reg1684 <= $signed((-{reg1650}));
            end
        end
    end
  assign wire1685 = $unsigned(((&(+(~reg1553))) ?
                        $signed($signed(reg27)) : (~^reg1642[(2'h2):(1'h0)])));
  module1686 #() modinst3486 (.wire1688(reg1575), .wire1687(reg1453), .wire1692(reg89), .clk(clk), .wire1691(reg1517), .wire1689(reg1479), .wire1690(reg1469), .y(wire3485));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1686
#(parameter param3483 = ((~{(((8'h9d) << (8'hbd)) ? ((8'hab) ? (8'hbd) : (7'h52)) : (-(7'h53))), {((8'hbb) > (7'h44)), {(7'h46), (8'ha5)}, (~^(8'ha0))}}) << {((8'hbc) ? (~&{(7'h55)}) : ({(7'h4f), (7'h4c), (8'hb9)} ? ((8'hab) ? (8'hb5) : (8'ha9)) : (&(8'hbf))))}), 
parameter param3484 = (param3483 > {(-(param3483 ? param3483 : param3483)), ((^~((8'hbd) != param3483)) || param3483)}))
(y, clk, wire1687, wire1688, wire1689, wire1690, wire1691, wire1692);
  output wire [(32'h23dd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h18):(1'h0)] wire1687;
  input wire [(5'h18):(1'h0)] wire1688;
  input wire [(5'h1c):(1'h0)] wire1689;
  input wire [(4'hf):(1'h0)] wire1690;
  input wire signed [(3'h6):(1'h0)] wire1691;
  input wire signed [(4'he):(1'h0)] wire1692;
  wire signed [(5'h19):(1'h0)] wire1693;
  wire signed [(5'h19):(1'h0)] wire1694;
  wire [(4'hc):(1'h0)] wire2946;
  wire [(2'h2):(1'h0)] wire2948;
  wire signed [(5'h1a):(1'h0)] wire3036;
  wire signed [(4'h9):(1'h0)] wire3070;
  wire [(5'h19):(1'h0)] wire3096;
  wire signed [(5'h11):(1'h0)] wire3147;
  wire signed [(4'hd):(1'h0)] wire3148;
  wire signed [(5'h14):(1'h0)] wire3268;
  wire [(5'h1f):(1'h0)] wire3364;
  wire [(5'h10):(1'h0)] wire3405;
  wire [(4'hb):(1'h0)] wire3406;
  wire [(5'h10):(1'h0)] wire3407;
  wire signed [(4'h9):(1'h0)] wire3408;
  wire signed [(5'h15):(1'h0)] wire3409;
  wire [(5'h11):(1'h0)] wire3410;
  wire [(5'h1d):(1'h0)] wire3479;
  wire [(5'h15):(1'h0)] wire3481;
  reg signed [(5'h1c):(1'h0)] reg3478 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3476 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3475 = (1'h0);
  reg [(4'he):(1'h0)] reg3471 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3469 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3466 = (1'h0);
  reg [(3'h6):(1'h0)] reg3465 = (1'h0);
  reg [(4'hd):(1'h0)] reg3464 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3463 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3462 = (1'h0);
  reg [(4'hb):(1'h0)] reg3461 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3460 = (1'h0);
  reg [(5'h11):(1'h0)] reg3457 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3454 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3449 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3448 = (1'h0);
  reg [(5'h17):(1'h0)] reg3447 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3443 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3439 = (1'h0);
  reg [(5'h15):(1'h0)] reg3438 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3437 = (1'h0);
  reg [(5'h18):(1'h0)] reg3436 = (1'h0);
  reg [(4'h9):(1'h0)] reg3435 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3434 = (1'h0);
  reg [(5'h13):(1'h0)] reg3431 = (1'h0);
  reg [(3'h5):(1'h0)] reg3430 = (1'h0);
  reg [(4'ha):(1'h0)] reg3428 = (1'h0);
  reg [(4'hf):(1'h0)] reg3420 = (1'h0);
  reg [(4'hd):(1'h0)] reg3419 = (1'h0);
  reg [(5'h14):(1'h0)] reg3417 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3416 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3415 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3414 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3412 = (1'h0);
  reg [(5'h16):(1'h0)] reg3411 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3404 = (1'h0);
  reg [(4'hc):(1'h0)] reg3403 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3402 = (1'h0);
  reg [(4'h9):(1'h0)] reg3400 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3396 = (1'h0);
  reg [(5'h11):(1'h0)] reg3395 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3392 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3384 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3383 = (1'h0);
  reg [(4'hc):(1'h0)] reg3376 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3380 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3374 = (1'h0);
  reg [(4'hc):(1'h0)] reg3373 = (1'h0);
  reg [(3'h6):(1'h0)] reg3372 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3370 = (1'h0);
  reg [(5'h18):(1'h0)] reg3367 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3362 = (1'h0);
  reg [(4'hc):(1'h0)] reg3361 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3359 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3354 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3351 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3349 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3348 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3346 = (1'h0);
  reg [(3'h6):(1'h0)] reg3345 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3344 = (1'h0);
  reg [(3'h4):(1'h0)] reg3343 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3341 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3340 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3338 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3337 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3334 = (1'h0);
  reg [(3'h7):(1'h0)] reg3333 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3332 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3324 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3323 = (1'h0);
  reg [(3'h5):(1'h0)] reg3322 = (1'h0);
  reg [(5'h17):(1'h0)] reg3316 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3312 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3311 = (1'h0);
  reg [(4'h9):(1'h0)] reg3310 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3309 = (1'h0);
  reg [(4'h8):(1'h0)] reg3308 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3304 = (1'h0);
  reg [(3'h6):(1'h0)] reg3300 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3298 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3297 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3296 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3295 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3293 = (1'h0);
  reg [(5'h11):(1'h0)] reg3288 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3284 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3280 = (1'h0);
  reg [(4'h8):(1'h0)] reg3277 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3273 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3267 = (1'h0);
  reg [(3'h7):(1'h0)] reg3266 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3265 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3262 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3261 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3258 = (1'h0);
  reg [(5'h14):(1'h0)] reg3257 = (1'h0);
  reg [(4'he):(1'h0)] reg3253 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3250 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3249 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3248 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3246 = (1'h0);
  reg [(4'hd):(1'h0)] reg3244 = (1'h0);
  reg [(4'hf):(1'h0)] reg3243 = (1'h0);
  reg [(4'hc):(1'h0)] reg3240 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3239 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3238 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3237 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3236 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3235 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3234 = (1'h0);
  reg [(5'h13):(1'h0)] reg3232 = (1'h0);
  reg [(4'h9):(1'h0)] reg3230 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3228 = (1'h0);
  reg [(4'hb):(1'h0)] reg3226 = (1'h0);
  reg [(4'hc):(1'h0)] reg3222 = (1'h0);
  reg [(5'h15):(1'h0)] reg3220 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3218 = (1'h0);
  reg [(4'h8):(1'h0)] reg3215 = (1'h0);
  reg [(4'ha):(1'h0)] reg3212 = (1'h0);
  reg [(2'h3):(1'h0)] reg3208 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3206 = (1'h0);
  reg [(5'h14):(1'h0)] reg3205 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3192 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3189 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3200 = (1'h0);
  reg [(5'h10):(1'h0)] reg3198 = (1'h0);
  reg [(5'h17):(1'h0)] reg3194 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3190 = (1'h0);
  reg [(5'h14):(1'h0)] reg3188 = (1'h0);
  reg [(3'h6):(1'h0)] reg3184 = (1'h0);
  reg [(5'h11):(1'h0)] reg3183 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3180 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3176 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3173 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3172 = (1'h0);
  reg [(5'h18):(1'h0)] reg3170 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3169 = (1'h0);
  reg [(5'h1b):(1'h0)] reg3168 = (1'h0);
  reg [(4'he):(1'h0)] reg3166 = (1'h0);
  reg [(5'h11):(1'h0)] reg3165 = (1'h0);
  reg [(4'h8):(1'h0)] reg3163 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3161 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3155 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3154 = (1'h0);
  reg [(5'h18):(1'h0)] reg3152 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3150 = (1'h0);
  reg [(5'h18):(1'h0)] reg3144 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3142 = (1'h0);
  reg [(5'h18):(1'h0)] reg3135 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3134 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3132 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3131 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3128 = (1'h0);
  reg [(3'h4):(1'h0)] reg3124 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3122 = (1'h0);
  reg [(5'h18):(1'h0)] reg3118 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3116 = (1'h0);
  reg [(5'h13):(1'h0)] reg3113 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3110 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3109 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3107 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3106 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3102 = (1'h0);
  reg [(2'h3):(1'h0)] reg3101 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3099 = (1'h0);
  reg [(4'ha):(1'h0)] reg3098 = (1'h0);
  reg [(3'h5):(1'h0)] reg3095 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3094 = (1'h0);
  reg [(5'h12):(1'h0)] reg3093 = (1'h0);
  reg [(3'h4):(1'h0)] reg3089 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3085 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3081 = (1'h0);
  reg [(2'h3):(1'h0)] reg3080 = (1'h0);
  reg [(5'h11):(1'h0)] reg3079 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3077 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3075 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3073 = (1'h0);
  reg [(3'h4):(1'h0)] reg3071 = (1'h0);
  reg [(3'h5):(1'h0)] reg3067 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3065 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3063 = (1'h0);
  reg [(3'h7):(1'h0)] reg3059 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3058 = (1'h0);
  reg [(4'h9):(1'h0)] reg3038 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3047 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3046 = (1'h0);
  reg [(5'h16):(1'h0)] reg3043 = (1'h0);
  reg [(5'h19):(1'h0)] reg3041 = (1'h0);
  reg [(4'h9):(1'h0)] reg3039 = (1'h0);
  reg [(5'h15):(1'h0)] reg3035 = (1'h0);
  reg [(2'h3):(1'h0)] reg3033 = (1'h0);
  reg [(5'h18):(1'h0)] reg3032 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3031 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3030 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3027 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3026 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3024 = (1'h0);
  reg [(5'h14):(1'h0)] reg3023 = (1'h0);
  reg [(5'h14):(1'h0)] reg3022 = (1'h0);
  reg [(5'h17):(1'h0)] reg3020 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3018 = (1'h0);
  reg [(3'h6):(1'h0)] reg3015 = (1'h0);
  reg [(5'h11):(1'h0)] reg3012 = (1'h0);
  reg [(5'h16):(1'h0)] reg3011 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3009 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3005 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3004 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3003 = (1'h0);
  reg [(5'h15):(1'h0)] reg3002 = (1'h0);
  reg [(2'h2):(1'h0)] reg3001 = (1'h0);
  reg [(4'h8):(1'h0)] reg2999 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2997 = (1'h0);
  reg [(5'h12):(1'h0)] reg2993 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2991 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2987 = (1'h0);
  reg [(4'hf):(1'h0)] reg2983 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2981 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2980 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2975 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2974 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2972 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2969 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2967 = (1'h0);
  reg [(5'h14):(1'h0)] reg2951 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2965 = (1'h0);
  reg [(4'hf):(1'h0)] reg2962 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2960 = (1'h0);
  reg [(5'h13):(1'h0)] reg2955 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2954 = (1'h0);
  reg [(3'h5):(1'h0)] reg2952 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2950 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2949 = (1'h0);
  reg [(2'h2):(1'h0)] reg3477 = (1'h0);
  reg [(5'h15):(1'h0)] reg3474 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar3473 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3472 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3470 = (1'h0);
  reg [(5'h13):(1'h0)] reg3468 = (1'h0);
  reg [(3'h7):(1'h0)] reg3467 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3459 = (1'h0);
  reg [(2'h3):(1'h0)] reg3458 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar3456 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3455 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3453 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar3452 = (1'h0);
  reg [(2'h3):(1'h0)] reg3451 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3450 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3446 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3445 = (1'h0);
  reg [(4'hc):(1'h0)] reg3444 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3442 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3441 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3440 = (1'h0);
  reg [(4'he):(1'h0)] reg3433 = (1'h0);
  reg [(2'h3):(1'h0)] reg3432 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3429 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3427 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3426 = (1'h0);
  reg [(4'he):(1'h0)] reg3425 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar3424 = (1'h0);
  reg [(4'hf):(1'h0)] reg3423 = (1'h0);
  reg [(4'hf):(1'h0)] reg3422 = (1'h0);
  reg [(4'hb):(1'h0)] reg3421 = (1'h0);
  reg [(2'h3):(1'h0)] reg3418 = (1'h0);
  reg [(3'h4):(1'h0)] reg3413 = (1'h0);
  reg [(5'h13):(1'h0)] reg3401 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3399 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3398 = (1'h0);
  reg [(4'h8):(1'h0)] reg3397 = (1'h0);
  reg [(4'hd):(1'h0)] reg3394 = (1'h0);
  reg [(2'h2):(1'h0)] reg3393 = (1'h0);
  reg [(5'h16):(1'h0)] reg3391 = (1'h0);
  reg [(5'h11):(1'h0)] reg3390 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3389 = (1'h0);
  reg [(5'h11):(1'h0)] reg3389 = (1'h0);
  reg [(5'h15):(1'h0)] reg3388 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3387 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3386 = (1'h0);
  reg [(2'h2):(1'h0)] reg3385 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3382 = (1'h0);
  reg [(5'h12):(1'h0)] reg3381 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3379 = (1'h0);
  reg [(2'h3):(1'h0)] reg3378 = (1'h0);
  reg [(5'h18):(1'h0)] reg3377 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar3376 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3375 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3371 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3369 = (1'h0);
  reg [(5'h12):(1'h0)] reg3368 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3366 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3365 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3339 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3332 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3363 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3360 = (1'h0);
  reg [(2'h2):(1'h0)] reg3358 = (1'h0);
  reg [(4'h9):(1'h0)] reg3357 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3356 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3355 = (1'h0);
  reg [(4'hb):(1'h0)] reg3353 = (1'h0);
  reg [(5'h13):(1'h0)] reg3352 = (1'h0);
  reg [(3'h6):(1'h0)] reg3350 = (1'h0);
  reg [(4'hd):(1'h0)] reg3347 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3342 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar3339 = (1'h0);
  reg [(2'h3):(1'h0)] reg3336 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3335 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3331 = (1'h0);
  reg [(5'h19):(1'h0)] reg3330 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3329 = (1'h0);
  reg [(4'h8):(1'h0)] reg3328 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3327 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3326 = (1'h0);
  reg [(4'hb):(1'h0)] reg3325 = (1'h0);
  reg [(4'hc):(1'h0)] reg3321 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3320 = (1'h0);
  reg [(5'h16):(1'h0)] reg3319 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3318 = (1'h0);
  reg [(4'hc):(1'h0)] reg3317 = (1'h0);
  reg [(5'h15):(1'h0)] reg3315 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3314 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3313 = (1'h0);
  reg [(2'h2):(1'h0)] reg3302 = (1'h0);
  reg [(4'hc):(1'h0)] reg3307 = (1'h0);
  reg [(3'h4):(1'h0)] reg3306 = (1'h0);
  reg [(4'h9):(1'h0)] reg3305 = (1'h0);
  reg [(4'hd):(1'h0)] reg3303 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar3302 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3301 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3299 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3294 = (1'h0);
  reg [(3'h7):(1'h0)] reg3292 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3291 = (1'h0);
  reg [(4'hd):(1'h0)] reg3290 = (1'h0);
  reg [(5'h16):(1'h0)] reg3289 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3287 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3286 = (1'h0);
  reg [(3'h4):(1'h0)] reg3285 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3283 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar3282 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3281 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3279 = (1'h0);
  reg [(2'h3):(1'h0)] reg3278 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3276 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3275 = (1'h0);
  reg [(5'h10):(1'h0)] reg3274 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3272 = (1'h0);
  reg [(5'h13):(1'h0)] forvar3271 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3270 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar3269 = (1'h0);
  reg [(5'h15):(1'h0)] reg3264 = (1'h0);
  reg [(3'h5):(1'h0)] reg3263 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3260 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3259 = (1'h0);
  reg [(5'h19):(1'h0)] reg3256 = (1'h0);
  reg [(5'h10):(1'h0)] reg3255 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3254 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3252 = (1'h0);
  reg [(4'h8):(1'h0)] reg3251 = (1'h0);
  reg [(4'he):(1'h0)] reg3247 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3245 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3242 = (1'h0);
  reg [(4'hd):(1'h0)] reg3241 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar3233 = (1'h0);
  reg [(4'h8):(1'h0)] reg3231 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3229 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3227 = (1'h0);
  reg [(5'h14):(1'h0)] reg3225 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3224 = (1'h0);
  reg [(5'h14):(1'h0)] reg3223 = (1'h0);
  reg [(4'hb):(1'h0)] reg3221 = (1'h0);
  reg [(5'h12):(1'h0)] reg3213 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3219 = (1'h0);
  reg [(5'h14):(1'h0)] reg3217 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg3216 = (1'h0);
  reg [(5'h1d):(1'h0)] reg3214 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3213 = (1'h0);
  reg [(4'ha):(1'h0)] reg3211 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3210 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3209 = (1'h0);
  reg [(2'h3):(1'h0)] reg3207 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3204 = (1'h0);
  reg [(5'h15):(1'h0)] reg3203 = (1'h0);
  reg [(4'he):(1'h0)] reg3199 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3196 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3202 = (1'h0);
  reg [(3'h5):(1'h0)] reg3201 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3199 = (1'h0);
  reg [(3'h6):(1'h0)] reg3197 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3196 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3195 = (1'h0);
  reg [(5'h10):(1'h0)] reg3193 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3192 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3191 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3189 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3187 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3186 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3185 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3182 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3181 = (1'h0);
  reg [(5'h14):(1'h0)] forvar3179 = (1'h0);
  reg [(5'h11):(1'h0)] reg3178 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3177 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3175 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3174 = (1'h0);
  reg [(5'h18):(1'h0)] reg3171 = (1'h0);
  reg [(5'h19):(1'h0)] reg3167 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3164 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3162 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3160 = (1'h0);
  reg [(2'h2):(1'h0)] reg3159 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3158 = (1'h0);
  reg [(4'h9):(1'h0)] reg3157 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3156 = (1'h0);
  reg [(4'hc):(1'h0)] reg3153 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar3151 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3149 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3146 = (1'h0);
  reg [(5'h13):(1'h0)] reg3145 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3143 = (1'h0);
  reg [(4'hf):(1'h0)] reg3141 = (1'h0);
  reg [(3'h7):(1'h0)] reg3140 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar3139 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar3138 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3137 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3136 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3133 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3130 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3129 = (1'h0);
  reg [(5'h14):(1'h0)] forvar3127 = (1'h0);
  reg [(4'hf):(1'h0)] reg3126 = (1'h0);
  reg [(5'h10):(1'h0)] reg3125 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3123 = (1'h0);
  reg [(5'h15):(1'h0)] reg3121 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3120 = (1'h0);
  reg [(4'he):(1'h0)] reg3119 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3117 = (1'h0);
  reg [(4'h9):(1'h0)] reg3115 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3114 = (1'h0);
  reg [(5'h1f):(1'h0)] reg3112 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar3111 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg3108 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3105 = (1'h0);
  reg [(5'h13):(1'h0)] reg3104 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3103 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg3100 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar3097 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar3092 = (1'h0);
  reg [(5'h13):(1'h0)] reg3091 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3090 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3088 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3087 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3086 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3084 = (1'h0);
  reg [(5'h1c):(1'h0)] reg3083 = (1'h0);
  reg [(5'h17):(1'h0)] reg3082 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3078 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3076 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3074 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3072 = (1'h0);
  reg [(4'ha):(1'h0)] reg3069 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar3068 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg3066 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3064 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3062 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3061 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar3060 = (1'h0);
  reg [(4'hd):(1'h0)] reg3048 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3046 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3039 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg3057 = (1'h0);
  reg [(5'h1e):(1'h0)] reg3056 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3055 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3054 = (1'h0);
  reg [(5'h19):(1'h0)] reg3053 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3052 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3051 = (1'h0);
  reg [(4'hc):(1'h0)] reg3050 = (1'h0);
  reg [(2'h3):(1'h0)] reg3049 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3048 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3045 = (1'h0);
  reg [(5'h14):(1'h0)] reg3044 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3042 = (1'h0);
  reg [(4'hb):(1'h0)] reg3040 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar3038 = (1'h0);
  reg [(5'h13):(1'h0)] reg3037 = (1'h0);
  reg [(4'h8):(1'h0)] reg3034 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3028 = (1'h0);
  reg [(5'h18):(1'h0)] reg3029 = (1'h0);
  reg [(5'h13):(1'h0)] reg3028 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3025 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar3021 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3019 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3017 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3016 = (1'h0);
  reg [(4'h8):(1'h0)] reg3014 = (1'h0);
  reg [(4'hb):(1'h0)] reg3013 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3010 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3008 = (1'h0);
  reg [(4'hc):(1'h0)] reg3007 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3006 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3000 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2998 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2996 = (1'h0);
  reg [(5'h17):(1'h0)] reg2995 = (1'h0);
  reg [(4'he):(1'h0)] forvar2994 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2992 = (1'h0);
  reg [(4'hf):(1'h0)] reg2990 = (1'h0);
  reg [(5'h19):(1'h0)] reg2989 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2988 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2986 = (1'h0);
  reg [(5'h11):(1'h0)] reg2985 = (1'h0);
  reg [(3'h6):(1'h0)] reg2984 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2982 = (1'h0);
  reg [(3'h4):(1'h0)] reg2979 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2978 = (1'h0);
  reg [(2'h2):(1'h0)] reg2977 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2976 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2973 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2971 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2970 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2968 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2956 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2966 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2964 = (1'h0);
  reg [(3'h7):(1'h0)] reg2963 = (1'h0);
  reg [(5'h16):(1'h0)] reg2961 = (1'h0);
  reg [(3'h7):(1'h0)] reg2959 = (1'h0);
  reg [(4'h8):(1'h0)] reg2958 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2957 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar2956 = (1'h0);
  reg [(5'h16):(1'h0)] reg2953 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2951 = (1'h0);
  assign y = {wire1693,
                 wire1694,
                 wire2946,
                 wire2948,
                 wire3036,
                 wire3070,
                 wire3096,
                 wire3147,
                 wire3148,
                 wire3268,
                 wire3364,
                 wire3405,
                 wire3406,
                 wire3407,
                 wire3408,
                 wire3409,
                 wire3410,
                 wire3479,
                 wire3481,
                 reg3478,
                 reg3476,
                 reg3475,
                 reg3471,
                 reg3469,
                 reg3466,
                 reg3465,
                 reg3464,
                 reg3463,
                 reg3462,
                 reg3461,
                 reg3460,
                 reg3457,
                 reg3454,
                 reg3449,
                 reg3448,
                 reg3447,
                 reg3443,
                 reg3439,
                 reg3438,
                 reg3437,
                 reg3436,
                 reg3435,
                 reg3434,
                 reg3431,
                 reg3430,
                 reg3428,
                 reg3420,
                 reg3419,
                 reg3417,
                 reg3416,
                 reg3415,
                 reg3414,
                 reg3412,
                 reg3411,
                 reg3404,
                 reg3403,
                 reg3402,
                 reg3400,
                 reg3396,
                 reg3395,
                 reg3392,
                 reg3384,
                 reg3383,
                 reg3376,
                 reg3380,
                 reg3374,
                 reg3373,
                 reg3372,
                 reg3370,
                 reg3367,
                 reg3362,
                 reg3361,
                 reg3359,
                 reg3354,
                 reg3351,
                 reg3349,
                 reg3348,
                 reg3346,
                 reg3345,
                 reg3344,
                 reg3343,
                 reg3341,
                 reg3340,
                 reg3338,
                 reg3337,
                 reg3334,
                 reg3333,
                 reg3332,
                 reg3324,
                 reg3323,
                 reg3322,
                 reg3316,
                 reg3312,
                 reg3311,
                 reg3310,
                 reg3309,
                 reg3308,
                 reg3304,
                 reg3300,
                 reg3298,
                 reg3297,
                 reg3296,
                 reg3295,
                 reg3293,
                 reg3288,
                 reg3284,
                 reg3280,
                 reg3277,
                 reg3273,
                 reg3267,
                 reg3266,
                 reg3265,
                 reg3262,
                 reg3261,
                 reg3258,
                 reg3257,
                 reg3253,
                 reg3250,
                 reg3249,
                 reg3248,
                 reg3246,
                 reg3244,
                 reg3243,
                 reg3240,
                 reg3239,
                 reg3238,
                 reg3237,
                 reg3236,
                 reg3235,
                 reg3234,
                 reg3232,
                 reg3230,
                 reg3228,
                 reg3226,
                 reg3222,
                 reg3220,
                 reg3218,
                 reg3215,
                 reg3212,
                 reg3208,
                 reg3206,
                 reg3205,
                 reg3192,
                 reg3189,
                 reg3200,
                 reg3198,
                 reg3194,
                 reg3190,
                 reg3188,
                 reg3184,
                 reg3183,
                 reg3180,
                 reg3176,
                 reg3173,
                 reg3172,
                 reg3170,
                 reg3169,
                 reg3168,
                 reg3166,
                 reg3165,
                 reg3163,
                 reg3161,
                 reg3155,
                 reg3154,
                 reg3152,
                 reg3150,
                 reg3144,
                 reg3142,
                 reg3135,
                 reg3134,
                 reg3132,
                 reg3131,
                 reg3128,
                 reg3124,
                 reg3122,
                 reg3118,
                 reg3116,
                 reg3113,
                 reg3110,
                 reg3109,
                 reg3107,
                 reg3106,
                 reg3102,
                 reg3101,
                 reg3099,
                 reg3098,
                 reg3095,
                 reg3094,
                 reg3093,
                 reg3089,
                 reg3085,
                 reg3081,
                 reg3080,
                 reg3079,
                 reg3077,
                 reg3075,
                 reg3073,
                 reg3071,
                 reg3067,
                 reg3065,
                 reg3063,
                 reg3059,
                 reg3058,
                 reg3038,
                 reg3047,
                 reg3046,
                 reg3043,
                 reg3041,
                 reg3039,
                 reg3035,
                 reg3033,
                 reg3032,
                 reg3031,
                 reg3030,
                 reg3027,
                 reg3026,
                 reg3024,
                 reg3023,
                 reg3022,
                 reg3020,
                 reg3018,
                 reg3015,
                 reg3012,
                 reg3011,
                 reg3009,
                 reg3005,
                 reg3004,
                 reg3003,
                 reg3002,
                 reg3001,
                 reg2999,
                 reg2997,
                 reg2993,
                 reg2991,
                 reg2987,
                 reg2983,
                 reg2981,
                 reg2980,
                 reg2975,
                 reg2974,
                 reg2972,
                 reg2969,
                 reg2967,
                 reg2951,
                 reg2965,
                 reg2962,
                 reg2960,
                 reg2955,
                 reg2954,
                 reg2952,
                 reg2950,
                 reg2949,
                 reg3477,
                 reg3474,
                 forvar3473,
                 reg3472,
                 reg3470,
                 reg3468,
                 reg3467,
                 forvar3459,
                 reg3458,
                 forvar3456,
                 reg3455,
                 reg3453,
                 forvar3452,
                 reg3451,
                 reg3450,
                 reg3446,
                 forvar3445,
                 reg3444,
                 reg3442,
                 reg3441,
                 reg3440,
                 reg3433,
                 reg3432,
                 reg3429,
                 reg3427,
                 forvar3426,
                 reg3425,
                 forvar3424,
                 reg3423,
                 reg3422,
                 reg3421,
                 reg3418,
                 reg3413,
                 reg3401,
                 reg3399,
                 forvar3398,
                 reg3397,
                 reg3394,
                 reg3393,
                 reg3391,
                 reg3390,
                 forvar3389,
                 reg3389,
                 reg3388,
                 reg3387,
                 reg3386,
                 reg3385,
                 reg3382,
                 reg3381,
                 reg3379,
                 reg3378,
                 reg3377,
                 forvar3376,
                 reg3375,
                 reg3371,
                 reg3369,
                 reg3368,
                 reg3366,
                 forvar3365,
                 reg3339,
                 forvar3332,
                 reg3363,
                 reg3360,
                 reg3358,
                 reg3357,
                 reg3356,
                 reg3355,
                 reg3353,
                 reg3352,
                 reg3350,
                 reg3347,
                 reg3342,
                 forvar3339,
                 reg3336,
                 reg3335,
                 reg3331,
                 reg3330,
                 reg3329,
                 reg3328,
                 reg3327,
                 reg3326,
                 reg3325,
                 reg3321,
                 reg3320,
                 reg3319,
                 forvar3318,
                 reg3317,
                 reg3315,
                 reg3314,
                 reg3313,
                 reg3302,
                 reg3307,
                 reg3306,
                 reg3305,
                 reg3303,
                 forvar3302,
                 reg3301,
                 reg3299,
                 reg3294,
                 reg3292,
                 forvar3291,
                 reg3290,
                 reg3289,
                 reg3287,
                 reg3286,
                 reg3285,
                 reg3283,
                 forvar3282,
                 forvar3281,
                 reg3279,
                 reg3278,
                 reg3276,
                 reg3275,
                 reg3274,
                 forvar3272,
                 forvar3271,
                 reg3270,
                 forvar3269,
                 reg3264,
                 reg3263,
                 reg3260,
                 reg3259,
                 reg3256,
                 reg3255,
                 reg3254,
                 reg3252,
                 reg3251,
                 reg3247,
                 reg3245,
                 reg3242,
                 reg3241,
                 forvar3233,
                 reg3231,
                 reg3229,
                 reg3227,
                 reg3225,
                 reg3224,
                 reg3223,
                 reg3221,
                 reg3213,
                 reg3219,
                 reg3217,
                 reg3216,
                 reg3214,
                 forvar3213,
                 reg3211,
                 reg3210,
                 reg3209,
                 reg3207,
                 forvar3204,
                 reg3203,
                 reg3199,
                 reg3196,
                 reg3202,
                 reg3201,
                 forvar3199,
                 reg3197,
                 forvar3196,
                 reg3195,
                 reg3193,
                 forvar3192,
                 reg3191,
                 forvar3189,
                 reg3187,
                 reg3186,
                 reg3185,
                 reg3182,
                 reg3181,
                 forvar3179,
                 reg3178,
                 reg3177,
                 reg3175,
                 reg3174,
                 reg3171,
                 reg3167,
                 reg3164,
                 reg3162,
                 reg3160,
                 reg3159,
                 reg3158,
                 reg3157,
                 reg3156,
                 reg3153,
                 forvar3151,
                 forvar3149,
                 reg3146,
                 reg3145,
                 reg3143,
                 reg3141,
                 reg3140,
                 forvar3139,
                 forvar3138,
                 reg3137,
                 reg3136,
                 reg3133,
                 reg3130,
                 reg3129,
                 forvar3127,
                 reg3126,
                 reg3125,
                 reg3123,
                 reg3121,
                 forvar3120,
                 reg3119,
                 reg3117,
                 reg3115,
                 reg3114,
                 reg3112,
                 forvar3111,
                 reg3108,
                 reg3105,
                 reg3104,
                 reg3103,
                 reg3100,
                 forvar3097,
                 forvar3092,
                 reg3091,
                 reg3090,
                 reg3088,
                 reg3087,
                 reg3086,
                 reg3084,
                 reg3083,
                 reg3082,
                 reg3078,
                 reg3076,
                 reg3074,
                 reg3072,
                 reg3069,
                 forvar3068,
                 reg3066,
                 reg3064,
                 reg3062,
                 forvar3061,
                 forvar3060,
                 reg3048,
                 forvar3046,
                 forvar3039,
                 reg3057,
                 reg3056,
                 reg3055,
                 reg3054,
                 reg3053,
                 reg3052,
                 reg3051,
                 reg3050,
                 reg3049,
                 forvar3048,
                 reg3045,
                 reg3044,
                 reg3042,
                 reg3040,
                 forvar3038,
                 reg3037,
                 reg3034,
                 forvar3028,
                 reg3029,
                 reg3028,
                 reg3025,
                 forvar3021,
                 reg3019,
                 reg3017,
                 reg3016,
                 reg3014,
                 reg3013,
                 forvar3010,
                 reg3008,
                 reg3007,
                 reg3006,
                 forvar3000,
                 reg2998,
                 reg2996,
                 reg2995,
                 forvar2994,
                 reg2992,
                 reg2990,
                 reg2989,
                 reg2988,
                 reg2986,
                 reg2985,
                 reg2984,
                 reg2982,
                 reg2979,
                 forvar2978,
                 reg2977,
                 reg2976,
                 reg2973,
                 reg2971,
                 forvar2970,
                 forvar2968,
                 reg2956,
                 reg2966,
                 reg2964,
                 reg2963,
                 reg2961,
                 reg2959,
                 reg2958,
                 reg2957,
                 forvar2956,
                 reg2953,
                 forvar2951,
                 (1'h0)};
  assign wire1693 = ($unsigned(((wire1689 > $signed((8'hab))) ?
                        ((wire1689 < (7'h57)) ?
                            wire1692 : $signed(wire1690)) : ({wire1692,
                            wire1691,
                            wire1690} != {wire1690,
                            wire1687,
                            wire1690}))) != (~|(wire1689 ?
                        (wire1692[(3'h4):(1'h0)] ?
                            (wire1689 ?
                                wire1689 : wire1687) : (+wire1687)) : ($unsigned(wire1689) * (wire1690 ?
                            wire1692 : wire1688)))));
  assign wire1694 = wire1690[(4'h9):(4'h8)];
  module1695 #() modinst2947 (wire2946, clk, wire1688, wire1694, wire1687, wire1693);
  assign wire2948 = $unsigned((+wire1688[(2'h3):(2'h3)]));
  always
    @(posedge clk) begin
      reg2949 <= ((8'hac) ? (|(!$unsigned($unsigned(wire1692)))) : wire1692);
      reg2950 <= $signed($unsigned($signed(wire2946[(3'h5):(2'h3)])));
      if (wire1690)
        begin
          for (forvar2951 = (1'h0); (forvar2951 < (3'h4)); forvar2951 = (forvar2951 + (1'h1)))
            begin
              reg2952 <= $unsigned(wire1694);
              reg2953 = (8'hae);
              reg2954 <= {($unsigned(({wire1692} ?
                          {wire1693, wire2946} : {wire1691})) ?
                      $unsigned($signed($unsigned(wire2946))) : (^wire1687[(5'h11):(3'h6)]))};
            end
          reg2955 <= $unsigned(((~|$signed($signed(reg2953))) || wire1691[(3'h5):(3'h4)]));
          for (forvar2956 = (1'h0); (forvar2956 < (1'h1)); forvar2956 = (forvar2956 + (1'h1)))
            begin
              reg2957 = reg2949;
              reg2958 = $signed($unsigned((&reg2950[(4'hb):(4'h8)])));
              reg2959 = forvar2956[(4'ha):(4'h9)];
              reg2960 <= ($unsigned($unsigned($unsigned(forvar2956[(5'h17):(1'h0)]))) >>> reg2958);
              reg2961 = $unsigned((8'hb5));
              reg2962 <= ($signed(reg2955[(4'h9):(2'h3)]) ?
                  wire1693[(3'h6):(2'h2)] : $signed(wire1694));
            end
          reg2963 = $unsigned(reg2953);
          if (wire1687[(2'h2):(1'h0)])
            begin
              reg2964 = $unsigned((forvar2951[(3'h6):(3'h5)] ?
                  $unsigned($unsigned($signed(forvar2951))) : (~|{reg2961[(4'hb):(3'h6)],
                      reg2952,
                      (wire1693 * reg2958)})));
            end
          else
            begin
              reg2965 <= reg2963;
            end
          reg2966 = (~|(($signed(((7'h51) ? reg2962 : reg2964)) ?
              {wire2946} : reg2958[(3'h6):(1'h0)]) < ({wire1691[(1'h1):(1'h1)],
              $unsigned(wire1692)} * ($signed(reg2955) ?
              {wire1688} : $unsigned(wire1694)))));
        end
      else
        begin
          if (forvar2951)
            begin
              reg2951 <= (7'h54);
              reg2953 = (!(reg2959[(1'h1):(1'h0)] * ($unsigned(reg2950[(3'h7):(3'h4)]) | ({wire1688,
                  reg2949} ^ (wire1694 >> (7'h50))))));
              reg2954 <= (^{$signed({(~&reg2966),
                      $signed(reg2965),
                      $signed(wire2948)})});
            end
          else
            begin
              reg2953 = $unsigned({((!$signed(reg2954)) == (8'ha1)), wire1694});
              reg2956 = {($unsigned((-(8'hbb))) ?
                      $unsigned(wire1691) : reg2965[(3'h7):(1'h1)])};
              reg2957 = $unsigned((((7'h48) >> ((wire1688 ^ (8'hae)) ?
                      reg2960[(3'h7):(3'h5)] : wire1694)) ?
                  wire1691[(2'h3):(2'h3)] : $signed($unsigned($signed(reg2950)))));
              reg2960 <= (((~(~^{reg2965, wire1692, wire2948})) ?
                      (($signed(wire1689) <<< (!reg2957)) ?
                          reg2953 : (!$signed(reg2955))) : $unsigned({reg2952[(3'h4):(3'h4)],
                          (wire2948 < wire1690),
                          $signed((8'hbe))})) ?
                  ($unsigned($unsigned((reg2956 ? reg2963 : reg2957))) ?
                      {$unsigned((^reg2964)),
                          ($signed((8'ha9)) ^ (~reg2957))} : {forvar2951[(5'h15):(4'ha)],
                          $unsigned($unsigned(wire2948)),
                          (~(reg2964 ? (8'hac) : wire1690))}) : wire1687);
              reg2961 = (wire2948[(1'h0):(1'h0)] ?
                  reg2960 : (reg2963 ?
                      (7'h4d) : $unsigned(reg2963[(1'h1):(1'h0)])));
              reg2963 = $signed(((^~(((8'hbe) ?
                      forvar2951 : wire1691) == ((7'h48) ?
                      wire1689 : (8'hbb)))) ?
                  $unsigned($signed(forvar2956)) : reg2965[(3'h4):(1'h0)]));
              reg2965 <= $signed($signed(({reg2965[(3'h4):(3'h4)],
                  wire1693,
                  $signed((8'ha9))} - wire1687)));
            end
        end
      reg2967 <= ((8'hb2) >>> ((({wire1687, (8'h9c)} <<< (reg2962 ?
              reg2950 : reg2951)) ?
          wire2948 : $unsigned(reg2951)) >>> wire1694[(5'h11):(4'hb)]));
      for (forvar2968 = (1'h0); (forvar2968 < (3'h5)); forvar2968 = (forvar2968 + (1'h1)))
        begin
          reg2969 <= (~^(({wire2948[(1'h1):(1'h1)]} && $unsigned($signed(wire2946))) ?
              $unsigned(reg2963) : (8'hbb)));
          for (forvar2970 = (1'h0); (forvar2970 < (3'h4)); forvar2970 = (forvar2970 + (1'h1)))
            begin
              reg2971 = $unsigned((((((8'haa) ? wire2946 : wire2946) ?
                      (7'h4f) : $signed(reg2960)) ?
                  $signed($signed(reg2965)) : ((7'h48) ?
                      $unsigned(reg2961) : (~&reg2963))) == (forvar2968[(3'h7):(3'h6)] <<< wire1687)));
              reg2972 <= (~|wire1692);
              reg2973 = ((~&(reg2951 ?
                      wire1690[(4'hd):(3'h6)] : $unsigned((-reg2951)))) ?
                  (8'hb2) : reg2963[(1'h1):(1'h0)]);
              reg2974 <= $signed($unsigned($unsigned((reg2973 ~^ $signed(reg2960)))));
              reg2975 <= wire1688;
            end
          reg2976 = (reg2972[(1'h0):(1'h0)] == (((!(reg2974 >= (8'h9e))) ^ ({reg2958,
                      reg2965,
                      reg2955} ?
                  {reg2972, wire1689} : reg2966)) ?
              (^~reg2953[(5'h10):(5'h10)]) : (reg2957[(4'hc):(1'h1)] & $signed($signed(reg2960)))));
          reg2977 = (~^$signed((~&(&$signed(forvar2968)))));
        end
      for (forvar2978 = (1'h0); (forvar2978 < (3'h4)); forvar2978 = (forvar2978 + (1'h1)))
        begin
          if ($unsigned(((reg2964[(2'h2):(1'h1)] ?
              $signed($signed(reg2958)) : ({(7'h58)} ^ reg2959[(3'h5):(3'h5)])) <= (-$signed($unsigned(reg2973))))))
            begin
              reg2979 = forvar2951;
              reg2980 <= ((~reg2951) ?
                  (reg2966 ^ $signed({reg2969,
                      (reg2977 ?
                          reg2953 : reg2954)})) : $unsigned({reg2957[(1'h0):(1'h0)],
                      (8'hb1)}));
              reg2981 <= reg2965[(1'h1):(1'h1)];
              reg2982 = {($signed((&((7'h58) || forvar2970))) ?
                      (wire2946[(1'h1):(1'h1)] ?
                          reg2963 : $signed($signed(forvar2978))) : {reg2975,
                          $signed($unsigned(wire1691)),
                          reg2958[(2'h2):(1'h1)]}),
                  ((!$signed((reg2972 ? reg2955 : reg2961))) >> reg2964),
                  reg2954};
            end
          else
            begin
              reg2979 = $unsigned({(((!reg2969) == {reg2958}) ?
                      wire1687 : reg2960)});
              reg2980 <= reg2966;
              reg2982 = (wire1692[(1'h1):(1'h0)] < $unsigned(($unsigned((~&reg2965)) > (~|reg2976))));
              reg2983 <= {reg2952[(3'h5):(2'h3)]};
              reg2984 = (|wire1692[(3'h6):(3'h5)]);
              reg2985 = $unsigned((~|{$unsigned((forvar2951 ?
                      reg2976 : (7'h58)))}));
            end
          if ($signed((&($unsigned((reg2985 ?
              reg2958 : (7'h44))) < $signed(wire1690[(1'h0):(1'h0)])))))
            begin
              reg2986 = (7'h50);
              reg2987 <= (reg2967[(5'h1a):(5'h19)] ?
                  (reg2955 ?
                      $unsigned(($unsigned(wire2946) ?
                          (8'ha0) : {reg2986,
                              (7'h4c),
                              reg2977})) : $unsigned(reg2975[(3'h5):(3'h4)])) : $unsigned($signed(($signed(wire1693) ?
                      reg2950[(3'h4):(2'h3)] : (reg2955 * reg2986)))));
              reg2988 = $unsigned((+($unsigned((reg2949 >> reg2951)) ?
                  forvar2951[(5'h17):(2'h2)] : reg2980[(2'h3):(2'h2)])));
              reg2989 = ($signed((reg2981 <= $unsigned(reg2984[(3'h4):(1'h1)]))) ?
                  $unsigned((~reg2953[(1'h0):(1'h0)])) : reg2969[(2'h2):(1'h0)]);
            end
          else
            begin
              reg2987 <= $signed((~|reg2973[(1'h1):(1'h0)]));
              reg2988 = ($signed(reg2954) ?
                  (-$unsigned($unsigned({(7'h4d),
                      reg2981}))) : ($signed((forvar2968[(4'hb):(1'h1)] ?
                          ((8'ha0) ? reg2982 : (8'ha6)) : $unsigned(reg2974))) ?
                      (~$unsigned((reg2963 ?
                          reg2971 : reg2975))) : $signed((-$signed((8'hbd))))));
              reg2989 = reg2986;
              reg2990 = reg2961;
              reg2991 <= (~&(reg2955[(5'h13):(4'ha)] ?
                  ((!$signed((8'hb8))) - ({wire2948, reg2966} ?
                      reg2985 : {reg2966, reg2983, reg2984})) : reg2973));
              reg2992 = $unsigned((~reg2988[(3'h5):(1'h0)]));
            end
          reg2993 <= ((|(^~reg2961[(2'h3):(1'h1)])) + $signed((8'h9d)));
          for (forvar2994 = (1'h0); (forvar2994 < (1'h0)); forvar2994 = (forvar2994 + (1'h1)))
            begin
              reg2995 = reg2980[(5'h12):(1'h1)];
              reg2996 = (~forvar2994);
              reg2997 <= (^$signed(wire1690));
              reg2998 = ((~^forvar2978) ?
                  $unsigned((&$signed(reg2962[(3'h4):(2'h2)]))) : ($unsigned((8'h9f)) ?
                      $unsigned({$unsigned(reg2954)}) : $signed($unsigned((&reg2977)))));
            end
          reg2999 <= {($signed($signed(reg2982)) ?
                  ({(reg2971 * reg2998), reg2974} - $signed((reg2958 ?
                      reg2986 : reg2975))) : wire1688[(4'he):(4'hb)])};
          for (forvar3000 = (1'h0); (forvar3000 < (3'h6)); forvar3000 = (forvar3000 + (1'h1)))
            begin
              reg3001 <= (^reg2989[(3'h7):(3'h5)]);
              reg3002 <= $signed((reg2995 - (($signed(reg2959) || wire1687) ?
                  reg2989[(1'h0):(1'h0)] : (|(forvar2994 ?
                      reg2995 : (7'h47))))));
              reg3003 <= $signed({reg2981,
                  ((|$signed(reg2966)) ?
                      {wire2946[(3'h6):(2'h3)]} : ($unsigned(reg2951) ?
                          $signed(reg2974) : $signed(reg2975)))});
              reg3004 <= (7'h4c);
              reg3005 <= {(&forvar3000), wire1694, $unsigned((~(8'hb7)))};
              reg3006 = $unsigned((~|(((reg2972 ? reg3001 : reg2996) ?
                  (reg2985 ? (7'h40) : (7'h55)) : {wire2948,
                      (7'h4f),
                      (7'h50)}) + forvar2968)));
              reg3007 = $signed((reg2973[(3'h5):(1'h1)] > {{(wire1689 != reg2988),
                      $signed(reg2998)}}));
            end
          reg3008 = $signed(reg3005[(1'h1):(1'h0)]);
        end
      reg3009 <= $signed(wire2946);
    end
  always
    @(posedge clk) begin
      for (forvar3010 = (1'h0); (forvar3010 < (3'h6)); forvar3010 = (forvar3010 + (1'h1)))
        begin
          reg3011 <= reg2954;
          if (wire1689)
            begin
              reg3012 <= $signed(reg2974[(4'hc):(2'h2)]);
              reg3013 = (|$signed({{(reg2962 ? (8'hab) : wire1691),
                      (reg2951 > wire1692),
                      $unsigned(reg2993)}}));
            end
          else
            begin
              reg3013 = $signed((~reg2993));
            end
          if ($unsigned($unsigned(((reg2955 ^~ $signed(reg3013)) <<< $unsigned(reg3013)))))
            begin
              reg3014 = reg3009;
              reg3015 <= reg3009;
              reg3016 = $signed({$signed(reg3001[(1'h1):(1'h1)])});
              reg3017 = (8'hba);
              reg3018 <= $unsigned(wire1687);
              reg3019 = (((&(reg3011 ?
                          $unsigned(reg2962) : $unsigned(reg2952))) ?
                      wire1688[(4'hd):(3'h5)] : (reg2954[(4'h8):(3'h5)] ^~ ($signed(reg2997) ?
                          (|reg2954) : $unsigned(reg2999)))) ?
                  ($signed(reg3009[(5'h10):(4'hf)]) != (((!reg2967) << wire1691[(3'h4):(1'h0)]) ~^ {reg2969[(3'h4):(2'h3)]})) : $signed((7'h51)));
            end
          else
            begin
              reg3014 = $signed(($signed($signed($signed(reg3017))) ?
                  reg3003[(5'h1b):(3'h7)] : wire1694[(3'h7):(3'h7)]));
              reg3015 <= (~$signed($unsigned(reg3001)));
              reg3016 = (forvar3010[(2'h3):(1'h1)] ?
                  reg3009[(4'hb):(4'h8)] : ($unsigned($unsigned($unsigned(wire1690))) ?
                      $unsigned({$unsigned(wire1687)}) : $signed($unsigned((wire2948 ?
                          reg3019 : wire1690)))));
              reg3017 = wire1692[(4'hc):(4'hc)];
              reg3019 = $signed(reg2967[(5'h1d):(4'he)]);
              reg3020 <= reg3014[(3'h4):(2'h2)];
            end
          for (forvar3021 = (1'h0); (forvar3021 < (1'h1)); forvar3021 = (forvar3021 + (1'h1)))
            begin
              reg3022 <= reg3016[(5'h16):(4'hb)];
            end
          reg3023 <= reg2975;
        end
      reg3024 <= ($unsigned((({wire1693} ?
          wire1689[(4'hf):(3'h7)] : $signed(reg2955)) >> $unsigned($unsigned((8'hbc))))) >>> (~($unsigned((reg2972 ?
          (7'h40) : reg2999)) & $signed((reg2975 ? reg2997 : reg3009)))));
    end
  always
    @(posedge clk) begin
      reg3025 = reg2969;
    end
  always
    @(posedge clk) begin
      reg3026 <= (({($signed(reg3009) ?
                      (reg2991 - reg2954) : $unsigned(reg3001)),
                  ((reg2972 <= reg2980) == reg2965[(3'h5):(3'h4)])} ?
              $unsigned((((7'h51) ?
                  reg2960 : reg3023) > (~reg2983))) : (reg2949[(4'h8):(4'h8)] >>> $signed(reg2954[(4'h9):(1'h1)]))) ?
          (reg2972 << $unsigned({$unsigned((7'h57)),
              wire1689})) : $signed(((reg2962 ^ (wire2946 ?
              reg2980 : reg3022)) << reg2969[(4'hc):(3'h4)])));
      if ((|reg3011))
        begin
          reg3027 <= ((~|$unsigned($unsigned({(8'ha3),
              wire1687}))) * reg2969[(3'h5):(2'h3)]);
          reg3028 = ((reg2997 ?
              wire1692[(1'h1):(1'h1)] : (((reg3005 ?
                      reg3004 : reg2952) | (wire2948 ? reg2972 : reg2983)) ?
                  $signed((wire1691 ?
                      reg3012 : wire1688)) : (|$signed(wire2948)))) * reg3022[(2'h2):(1'h0)]);
          reg3029 = reg3011;
        end
      else
        begin
          reg3027 <= $unsigned($signed($signed(wire1691)));
          for (forvar3028 = (1'h0); (forvar3028 < (1'h1)); forvar3028 = (forvar3028 + (1'h1)))
            begin
              reg3029 = (-reg3001);
              reg3030 <= $unsigned($unsigned(wire2948));
              reg3031 <= (7'h4a);
            end
          reg3032 <= reg2997[(5'h19):(5'h14)];
        end
      reg3033 <= ((~|(|$signed(wire2948[(2'h2):(2'h2)]))) ?
          $unsigned((~^reg2955)) : $signed(($unsigned(reg3026) ?
              ($unsigned(reg2951) ?
                  (reg3032 ?
                      reg2980 : wire1689) : ((8'hb6) >>> reg2967)) : reg3028)));
      reg3034 = reg2975;
      reg3035 <= (!reg3028);
    end
  assign wire3036 = ($signed($unsigned((~{reg3003}))) ?
                        $unsigned(reg3015[(3'h4):(2'h3)]) : (&$unsigned(((reg2983 ~^ wire2946) > reg3027[(1'h0):(1'h0)]))));
  always
    @(posedge clk) begin
      if ({wire1688[(1'h0):(1'h0)],
          {({reg3027[(1'h1):(1'h1)]} && {wire2946[(1'h1):(1'h1)],
                  $unsigned(reg3032)}),
              (+($signed(reg2962) ? $signed((7'h40)) : reg2980)),
              ({{reg2965}} ?
                  ((8'haf) * reg2975[(1'h0):(1'h0)]) : $unsigned($unsigned(wire1687)))},
          ((reg3032 ?
                  $signed((!reg2981)) : ((~^reg2954) ?
                      ((8'hb7) ? wire1691 : reg3023) : (reg3018 >>> reg3026))) ?
              (((reg3002 & reg2949) ? wire1690 : $signed((7'h56))) ?
                  $signed((reg3009 == wire1690)) : $unsigned(((7'h53) ?
                      reg3035 : wire1694))) : {reg2983[(4'hc):(4'ha)],
                  (reg3023[(3'h6):(3'h4)] ~^ {reg3027}),
                  (-reg2951)})})
        begin
          reg3037 = reg2987[(1'h1):(1'h0)];
          for (forvar3038 = (1'h0); (forvar3038 < (3'h6)); forvar3038 = (forvar3038 + (1'h1)))
            begin
              reg3039 <= reg2962;
              reg3040 = (reg3020 == (wire1690[(4'h8):(4'h8)] ^ ((8'hb0) * {(reg2975 || reg2993),
                  $unsigned(wire2948),
                  {reg2950}})));
              reg3041 <= reg2983[(4'hf):(4'hd)];
              reg3042 = wire1694[(5'h12):(4'hc)];
              reg3043 <= {((|$unsigned((wire1694 ?
                      reg3004 : wire1690))) - $unsigned(((wire2946 ~^ reg2997) ?
                      (reg2991 ? reg2954 : reg2981) : (~|wire1688))))};
              reg3044 = $unsigned(reg2983);
              reg3045 = reg3009;
            end
          reg3046 <= ((~^$signed(wire1691)) || reg3004);
          reg3047 <= (($signed(reg2967) >> (~&reg3033[(2'h2):(1'h1)])) * reg3004);
          for (forvar3048 = (1'h0); (forvar3048 < (1'h0)); forvar3048 = (forvar3048 + (1'h1)))
            begin
              reg3049 = ((^~$signed({reg2965[(2'h3):(2'h3)], {reg3020}})) ?
                  (wire1687 ?
                      (((reg2962 * reg2952) > $signed(reg2983)) < $unsigned($signed((8'hb8)))) : $unsigned(reg2987)) : {($unsigned(reg3026) ?
                          ((reg3035 ? (7'h43) : wire1688) ?
                              $unsigned(reg3035) : $signed(reg3037)) : {wire1693,
                              reg3009,
                              (reg2952 ? forvar3048 : reg3018)}),
                      (((reg3024 ? reg3002 : reg3022) ?
                          (~^reg2999) : reg3020[(4'hb):(4'h9)]) || reg3024)});
              reg3050 = (~&(~|($unsigned((reg2993 == reg2997)) ?
                  reg2949[(4'hb):(3'h6)] : (((8'haf) ?
                      reg2969 : reg3018) != (~^wire1687)))));
              reg3051 = reg3003[(5'h13):(4'hc)];
              reg3052 = $signed(reg3022[(4'ha):(4'ha)]);
              reg3053 = reg3003[(4'hf):(3'h7)];
              reg3054 = ((reg3035[(5'h13):(4'hd)] ?
                  {((reg3042 ~^ reg2991) ? (reg3022 || reg3051) : (|reg3032)),
                      wire1694[(3'h4):(2'h3)]} : wire2948[(1'h1):(1'h0)]) * ({reg2951[(2'h3):(1'h1)],
                      (7'h40),
                      $signed(reg2960)} ?
                  $signed(forvar3048[(1'h1):(1'h1)]) : {reg3040[(3'h4):(3'h4)],
                      (^~reg3012),
                      (wire1694[(4'hf):(3'h6)] ?
                          (reg3020 ? reg3042 : reg3041) : (!reg2955))}));
              reg3055 = (&reg2991[(4'ha):(3'h4)]);
            end
          reg3056 = reg3032;
          reg3057 = ({reg2969,
                  $unsigned({$unsigned(reg2975), $unsigned(reg3040)}),
                  reg2950} ?
              (reg3022 | reg3031) : reg3001[(1'h1):(1'h0)]);
        end
      else
        begin
          reg3038 <= $signed((+$signed($unsigned(wire1690[(4'hb):(1'h0)]))));
          for (forvar3039 = (1'h0); (forvar3039 < (3'h4)); forvar3039 = (forvar3039 + (1'h1)))
            begin
              reg3040 = $unsigned(($signed((~(reg2987 ?
                  reg3055 : (7'h52)))) ~^ reg3040[(4'h8):(3'h4)]));
              reg3041 <= $unsigned((reg2969 ?
                  $unsigned(reg3023[(3'h7):(3'h6)]) : reg2969[(4'h9):(1'h0)]));
              reg3043 <= (!$unsigned(({reg3023[(5'h13):(5'h12)],
                      (wire2946 <<< reg3051),
                      (reg3051 ? reg2993 : (8'hb2))} ?
                  {((7'h53) ? reg3033 : reg2991),
                      (~&reg2949)} : (reg3041[(5'h16):(3'h5)] ?
                      wire1689 : $signed((8'hba))))));
              reg3044 = (reg3027 ?
                  reg2980[(4'h9):(2'h2)] : ($signed((&(reg3024 | wire2946))) + (($signed(reg3039) ?
                      ((7'h54) && (8'hb3)) : (reg3002 ?
                          (8'hb8) : reg3031)) >>> $unsigned($signed(forvar3039)))));
            end
          reg3045 = ((|reg3027[(1'h0):(1'h0)]) || $unsigned(((!reg3023[(4'hb):(2'h2)]) ?
              wire1691[(3'h5):(1'h1)] : ($signed(forvar3039) == $unsigned(reg2999)))));
          for (forvar3046 = (1'h0); (forvar3046 < (2'h2)); forvar3046 = (forvar3046 + (1'h1)))
            begin
              reg3048 = $unsigned(((~^$unsigned(reg3018[(5'h1a):(5'h16)])) + (8'hb1)));
              reg3049 = $unsigned(reg3003[(4'h9):(2'h3)]);
              reg3058 <= {reg3048[(3'h6):(3'h5)]};
            end
        end
      reg3059 <= (&wire1691[(2'h2):(1'h0)]);
      for (forvar3060 = (1'h0); (forvar3060 < (2'h2)); forvar3060 = (forvar3060 + (1'h1)))
        begin
          for (forvar3061 = (1'h0); (forvar3061 < (3'h5)); forvar3061 = (forvar3061 + (1'h1)))
            begin
              reg3062 = (~&reg3057);
              reg3063 <= (($unsigned(reg2960[(4'ha):(3'h6)]) && reg2962) == reg3053[(4'ha):(1'h1)]);
              reg3064 = $signed((reg3018[(4'hc):(4'ha)] > $unsigned($unsigned(reg3009))));
            end
          reg3065 <= ((~$unsigned(reg3002[(4'h8):(3'h5)])) ?
              $signed((reg3011 ?
                  reg3033[(1'h1):(1'h0)] : (^~$unsigned(reg2955)))) : forvar3060[(5'h11):(4'h9)]);
          reg3066 = {wire1694[(3'h6):(3'h6)], reg2980};
          reg3067 <= ((+(7'h49)) ?
              $signed(reg2993[(1'h0):(1'h0)]) : ((^(|((7'h48) ?
                  reg2962 : reg3001))) * reg3048));
          for (forvar3068 = (1'h0); (forvar3068 < (3'h4)); forvar3068 = (forvar3068 + (1'h1)))
            begin
              reg3069 = ($unsigned(reg3042) ?
                  {(^((-reg3020) & reg3002)), reg3059} : $unsigned((reg3049 ?
                      (reg3024[(3'h4):(2'h3)] - (&(8'ha8))) : $signed($signed(reg3035)))));
            end
        end
    end
  assign wire3070 = ({reg3032, (-(reg3063 ? $unsigned(reg3038) : wire3036))} ?
                        {reg3043,
                            (~|((!(8'hac)) ?
                                {reg3027} : $signed(wire1687)))} : $unsigned(reg3032[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      reg3071 <= $unsigned(reg3033);
      if (wire1694)
        begin
          if ($unsigned({((reg3026[(1'h0):(1'h0)] ?
                      (reg3002 >= wire3036) : reg3003) ?
                  ((|reg3063) && reg3043[(1'h0):(1'h0)]) : reg3043)}))
            begin
              reg3072 = $unsigned($signed($unsigned((|(~&reg3041)))));
              reg3073 <= (7'h49);
              reg3074 = (&(($signed($signed(reg3033)) - ($signed(wire1693) ?
                      (8'haa) : $unsigned(reg3067))) ?
                  $unsigned(reg2983[(4'hc):(4'hc)]) : ($signed((~reg2993)) > reg2954[(2'h3):(1'h0)])));
              reg3075 <= reg2993[(2'h3):(2'h3)];
              reg3076 = ((((8'hb1) && (|$unsigned(reg3073))) ?
                      (((reg3022 ? (8'h9d) : reg3024) ?
                              $unsigned(reg3001) : (wire1690 <= wire1688)) ?
                          wire1693 : reg3003[(4'hb):(2'h2)]) : reg2993[(3'h5):(3'h5)]) ?
                  $unsigned(reg3047[(4'h8):(1'h1)]) : (~^{(reg3003 >> $unsigned(reg2993))}));
              reg3077 <= $unsigned($unsigned((($unsigned(reg3032) || reg2969[(1'h1):(1'h1)]) >= ({reg2962,
                  reg3015} <<< (-reg3072)))));
              reg3078 = ({(wire3036[(4'h9):(2'h2)] ?
                          reg3043 : (|wire2946[(3'h5):(1'h0)])),
                      reg3072} ?
                  $unsigned(wire1692[(4'ha):(4'h9)]) : (&$unsigned((~^((8'hb9) ?
                      wire1688 : reg3077)))));
            end
          else
            begin
              reg3073 <= reg2965[(3'h4):(1'h1)];
              reg3074 = reg2955;
              reg3075 <= ($signed((&{$signed(reg3041)})) ?
                  reg2967[(5'h13):(5'h13)] : (7'h41));
              reg3077 <= $unsigned($signed((^reg3004[(1'h0):(1'h0)])));
              reg3079 <= wire1692[(4'hb):(3'h6)];
              reg3080 <= {((reg3058[(3'h7):(3'h6)] - (reg3076[(5'h11):(4'h9)] ?
                          ((7'h56) ? reg2983 : (7'h4a)) : {reg3059, (8'hab)})) ?
                      $unsigned($signed((reg3058 ?
                          reg2983 : reg2991))) : (($signed(reg2960) + (reg3026 * reg3046)) * (~&reg3026[(3'h4):(2'h3)]))),
                  reg3033,
                  ($signed($unsigned((reg3073 <<< reg3074))) ?
                      (~($unsigned((8'hbd)) ?
                          {wire1692,
                              reg3046} : reg3074[(3'h7):(1'h0)])) : $unsigned((|reg3001[(1'h0):(1'h0)])))};
              reg3081 <= (reg3015[(3'h5):(3'h5)] ?
                  (~&({(reg2993 ? reg3003 : reg2983),
                          (reg2981 ? reg3067 : wire1689)} ?
                      {(reg3073 ?
                              reg3079 : reg3039)} : $signed($unsigned(reg3032)))) : wire1693[(4'hc):(2'h2)]);
            end
          if ($unsigned(reg2951))
            begin
              reg3082 = reg3078;
              reg3083 = $unsigned(reg2993[(4'hf):(3'h6)]);
              reg3084 = ($unsigned($signed($signed(reg3078))) ?
                  (^~wire1690[(4'h8):(4'h8)]) : (^$unsigned(reg3027[(1'h0):(1'h0)])));
              reg3085 <= (reg2967 <<< $signed((((~|reg2960) ?
                      reg3011[(4'ha):(3'h5)] : $unsigned(reg2974)) ?
                  (reg3081[(3'h6):(3'h6)] & $unsigned((8'ha5))) : (8'ha0))));
              reg3086 = (reg3074 ?
                  $unsigned(($unsigned(reg2987) ?
                      ($unsigned((8'hb6)) ?
                          $unsigned(reg3009) : (~|reg3067)) : ({reg3081,
                          reg2987} + (8'ha6)))) : reg3082);
              reg3087 = $unsigned(reg3027);
              reg3088 = (+reg2999);
            end
          else
            begin
              reg3082 = wire1688[(2'h2):(2'h2)];
              reg3085 <= ((reg2960[(3'h6):(1'h0)] ?
                  (~&(reg3063 <<< (reg3031 >>> reg2962))) : $unsigned(((reg2980 ?
                          reg2967 : (8'hb9)) ?
                      reg3065 : (reg2999 | reg3011)))) * (-((+reg3058) <= {{reg3081,
                      reg3076,
                      (8'hab)},
                  (-reg3041),
                  reg3086})));
            end
        end
      else
        begin
          if ($unsigned((^($unsigned($signed(reg3022)) << $unsigned($unsigned(reg3004))))))
            begin
              reg3072 = $signed($unsigned($signed(reg2975[(2'h3):(2'h2)])));
            end
          else
            begin
              reg3073 <= reg2972[(1'h0):(1'h0)];
              reg3075 <= $unsigned((reg2987[(3'h5):(1'h0)] ?
                  ({reg3030[(5'h12):(3'h5)]} * ($signed(reg3082) ?
                      (reg2965 < wire3036) : $signed(reg3078))) : (wire1689 == wire1689[(5'h1a):(4'he)])));
            end
          reg3077 <= (+reg3001);
          if ($unsigned(reg3032[(1'h0):(1'h0)]))
            begin
              reg3078 = {(reg2987[(3'h4):(2'h2)] == $signed($signed(reg3020[(2'h3):(1'h1)]))),
                  $unsigned({((+reg2983) || reg2993[(2'h2):(1'h0)]),
                      reg2967[(5'h1c):(3'h4)],
                      $signed((!reg2981))}),
                  $signed({wire1692, reg3023, reg3038[(3'h4):(3'h4)]})};
              reg3082 = (~|(~|((reg2952 ?
                  (reg3086 >= reg2969) : reg3011) ^ ((reg3022 - reg3039) && $signed(reg2997)))));
              reg3083 = $unsigned(reg3079[(3'h6):(3'h5)]);
            end
          else
            begin
              reg3078 = $signed($unsigned((reg3027 ?
                  $signed(((7'h4d) ~^ reg3088)) : {(!reg3041), (^~reg3038)})));
              reg3082 = (~^$unsigned($unsigned((&(reg3085 < reg2954)))));
              reg3083 = ($unsigned((((~^reg2997) ?
                  (reg3030 ?
                      reg3027 : wire3036) : ((8'hb4) >> (8'hbf))) | $unsigned((reg3059 > reg3073)))) * (|$unsigned($unsigned((reg3023 > reg3087)))));
              reg3085 <= $signed(wire3070[(2'h2):(1'h0)]);
              reg3089 <= $signed(reg3009[(5'h11):(2'h2)]);
              reg3090 = ((-((~(reg2981 ?
                  (7'h48) : reg2972)) ^~ $unsigned($signed(wire2948)))) ~^ ($unsigned(reg2955[(3'h7):(2'h3)]) ?
                  $signed($unsigned((~&wire3036))) : (|$signed((reg3033 << reg2975)))));
            end
          reg3091 = $unsigned(reg3015[(3'h4):(2'h2)]);
          for (forvar3092 = (1'h0); (forvar3092 < (2'h2)); forvar3092 = (forvar3092 + (1'h1)))
            begin
              reg3093 <= {(wire2948 ?
                      reg3012[(1'h0):(1'h0)] : {reg2955,
                          {reg2974,
                              (wire2946 ? reg3046 : reg2969),
                              (~wire2948)}})};
              reg3094 <= ($unsigned((forvar3092[(3'h7):(3'h7)] < ($unsigned(reg3030) & {(8'ha1),
                      wire1694}))) ?
                  $signed((reg2949[(5'h18):(4'hf)] ^~ reg3038[(2'h2):(2'h2)])) : {{$signed({reg3038}),
                          ((reg3033 ? reg3071 : wire2946) ?
                              reg3087[(4'hd):(4'h8)] : (~&(8'h9f)))}});
            end
        end
      reg3095 <= reg3085;
    end
  assign wire3096 = (~($unsigned($signed(reg3063[(5'h13):(4'h8)])) ?
                        reg3081 : ($unsigned((8'hb6)) ?
                            $unsigned({reg2999, (8'haa)}) : (^{reg3059,
                                reg2952}))));
  always
    @(posedge clk) begin
      for (forvar3097 = (1'h0); (forvar3097 < (2'h2)); forvar3097 = (forvar3097 + (1'h1)))
        begin
          reg3098 <= (+(^$unsigned(((!reg2983) | reg2955[(4'ha):(4'h8)]))));
          if ($unsigned(((8'hb7) ?
              (~^reg2974) : $signed(reg2999[(1'h1):(1'h0)]))))
            begin
              reg3099 <= ($signed((($unsigned(reg2960) | $signed(reg2954)) ?
                      {((8'haa) ? reg3095 : reg3023),
                          $unsigned((8'haa))} : $unsigned((~reg3095)))) ?
                  ((reg2993[(4'hd):(3'h6)] + ((~reg3046) >>> $signed(reg2993))) - $signed(((reg3047 == reg3022) || (reg2969 | reg2952)))) : {(8'had),
                      {((reg2974 ? reg3063 : reg2950) ?
                              ((7'h43) ? reg2972 : reg3080) : (reg3032 ?
                                  reg2980 : wire1690)),
                          wire1691[(3'h6):(1'h0)]}});
              reg3100 = (^~(~&$unsigned(wire1694)));
              reg3101 <= (+($unsigned((7'h51)) | $signed({wire1691[(1'h1):(1'h1)],
                  (~|reg3059),
                  (reg3032 ? reg3002 : reg3003)})));
              reg3102 <= (reg2954 ?
                  ($unsigned(reg3039[(1'h1):(1'h0)]) ?
                      (&(7'h4d)) : ($signed((reg3039 ?
                          reg3073 : (8'ha0))) - (wire1693[(2'h3):(1'h0)] ?
                          (!reg3071) : $signed(reg3094)))) : $signed((^reg3080)));
              reg3103 = (+$signed(reg3065));
              reg3104 = (~&(reg3095[(2'h2):(2'h2)] * reg3094[(2'h3):(1'h1)]));
              reg3105 = $signed($unsigned((~&$signed(reg3079))));
            end
          else
            begin
              reg3099 <= (+$signed(wire1688[(4'h9):(4'h9)]));
              reg3101 <= $signed((~^(~&(!reg3020))));
              reg3103 = ({(^$unsigned(reg3038)),
                      (&$signed($signed(reg2969))),
                      $unsigned($signed(reg3035[(5'h10):(4'hc)]))} ?
                  $unsigned((^((reg3081 >> (8'hb2)) << $signed(reg2997)))) : $signed(((reg3077 ?
                          {reg3031, reg3081} : (~|reg3077)) ?
                      reg3063[(1'h1):(1'h1)] : (((8'ha8) >>> reg2975) ?
                          reg3094[(1'h0):(1'h0)] : $signed(reg3100)))));
              reg3106 <= {$unsigned($signed(reg3103[(4'h9):(3'h7)]))};
              reg3107 <= reg2955;
              reg3108 = $signed((^~$unsigned((|(reg2960 >>> reg3002)))));
            end
        end
      reg3109 <= (^~(^(reg3020 ? reg3035[(4'hc):(3'h6)] : (8'ha6))));
      reg3110 <= $signed(reg3015[(3'h4):(2'h3)]);
      for (forvar3111 = (1'h0); (forvar3111 < (3'h5)); forvar3111 = (forvar3111 + (1'h1)))
        begin
          if (reg3022[(4'ha):(3'h4)])
            begin
              reg3112 = {reg3024,
                  ((8'haa) >> ($signed(wire1688[(2'h3):(1'h0)]) ?
                      $signed($unsigned(forvar3097)) : ((reg3081 >> (7'h51)) ?
                          (8'hab) : (!reg3081)))),
                  (($signed({reg3110}) ?
                          (-wire1694) : {(reg3102 ? reg2974 : reg3079)}) ?
                      (+reg3073[(1'h1):(1'h1)]) : $unsigned({reg3046[(1'h1):(1'h0)],
                          {reg2987},
                          $signed(reg3023)}))};
            end
          else
            begin
              reg3112 = $signed($unsigned(reg2955));
            end
          if (wire1688[(5'h10):(3'h7)])
            begin
              reg3113 <= (reg3039 ~^ reg3030[(2'h2):(1'h1)]);
            end
          else
            begin
              reg3114 = wire1688[(2'h3):(1'h1)];
              reg3115 = ((^~reg3015[(2'h2):(1'h0)]) ?
                  $signed({(reg2962 ?
                          (reg3098 ? reg2980 : reg3023) : {reg3067,
                              reg2981,
                              reg3108}),
                      reg3103}) : (reg3039[(3'h5):(2'h3)] ?
                      reg3109 : (reg3015 > reg2987[(2'h2):(2'h2)])));
              reg3116 <= ({$signed((8'hbf))} <<< ($unsigned((8'ha0)) >>> (reg3058[(4'he):(3'h4)] < (wire3036 ?
                  (reg3027 ? reg3059 : reg2949) : $signed(reg3047)))));
              reg3117 = (+reg3022);
              reg3118 <= reg2950;
              reg3119 = $signed({forvar3111,
                  (^~(8'h9e)),
                  (~^($unsigned(reg3089) ?
                      (reg2954 ? (7'h4a) : reg3027) : $signed(reg3089)))});
            end
          for (forvar3120 = (1'h0); (forvar3120 < (1'h0)); forvar3120 = (forvar3120 + (1'h1)))
            begin
              reg3121 = $unsigned((|reg2983[(4'hd):(4'h8)]));
              reg3122 <= (-reg3089);
              reg3123 = $unsigned($signed(reg3003));
              reg3124 <= reg3105[(1'h1):(1'h1)];
              reg3125 = reg3012;
              reg3126 = {$signed($signed((reg2972[(1'h1):(1'h1)] >>> reg3058[(4'h9):(2'h3)])))};
            end
          for (forvar3127 = (1'h0); (forvar3127 < (3'h6)); forvar3127 = (forvar3127 + (1'h1)))
            begin
              reg3128 <= reg3115;
              reg3129 = $signed(reg3015);
              reg3130 = ((|$signed(reg2975[(3'h4):(1'h1)])) ?
                  (((7'h4b) ?
                          (~$unsigned(reg3030)) : ($unsigned(forvar3111) ^ (reg2993 ?
                              reg2972 : reg2950))) ?
                      ({(reg2967 && (7'h52)),
                          wire3036[(5'h18):(5'h12)]} >= ($signed(wire1692) ?
                          ((7'h57) != (8'hbe)) : (reg3119 ^ reg3023))) : $unsigned($signed((~reg3077)))) : reg2955[(5'h10):(4'h9)]);
              reg3131 <= (~|{((~reg3105[(1'h1):(1'h0)]) ?
                      {reg3105,
                          (~&(8'h9d)),
                          (reg3077 <= reg3041)} : $signed(reg3073)),
                  $unsigned(reg3065),
                  reg3123[(2'h3):(2'h2)]});
              reg3132 <= (reg2969 * ($signed((^~(~reg3030))) || (^$unsigned($signed((8'ha5))))));
              reg3133 = reg3099;
              reg3134 <= (reg3065[(3'h7):(2'h2)] ?
                  (~&reg3046[(5'h15):(5'h12)]) : (reg3033[(1'h0):(1'h0)] ?
                      $unsigned((~|{reg2997,
                          reg3035})) : $signed((^reg3027[(2'h2):(1'h0)]))));
            end
          reg3135 <= $signed((((^reg3114) == reg3024) * (+(reg3130[(4'ha):(4'ha)] | ((8'ha2) >>> reg3004)))));
          reg3136 = (($signed((reg3005[(5'h12):(1'h1)] ?
                      $signed(reg3129) : {reg3103})) ?
                  (reg2974 >= reg3075[(5'h13):(4'hd)]) : $signed(reg3129[(5'h10):(4'ha)])) ?
              forvar3120[(4'h8):(1'h0)] : reg3134[(4'hb):(1'h1)]);
          reg3137 = $unsigned(({($signed((8'h9f)) >> $signed((8'hb5))),
              $unsigned($signed(reg3101)),
              (-reg3109[(5'h10):(4'ha)])} < $signed($unsigned($signed(reg2962)))));
        end
      for (forvar3138 = (1'h0); (forvar3138 < (3'h5)); forvar3138 = (forvar3138 + (1'h1)))
        begin
          for (forvar3139 = (1'h0); (forvar3139 < (3'h5)); forvar3139 = (forvar3139 + (1'h1)))
            begin
              reg3140 = reg2980[(5'h12):(3'h6)];
              reg3141 = $unsigned((reg2960[(2'h3):(2'h2)] ?
                  (~((8'hb8) ?
                      (reg3131 ?
                          reg3089 : wire3070) : $signed(reg2950))) : (reg2999[(4'h8):(3'h4)] == (|$signed(reg2993)))));
            end
          if (wire1689[(5'h13):(4'h8)])
            begin
              reg3142 <= (!reg3075);
            end
          else
            begin
              reg3143 = ($signed(reg3128[(4'hc):(2'h2)]) == $signed(((reg3103[(4'ha):(3'h4)] ?
                      (reg3041 ? reg3041 : reg3142) : $signed(reg2991)) ?
                  {(~reg3102)} : (~&((8'h9c) < reg3027)))));
              reg3144 <= (~|(({(wire2948 < reg3023)} >= {(8'h9c)}) ?
                  ({{(8'ha0),
                          (8'hac)}} - reg3030) : $unsigned($signed($signed(reg2983)))));
              reg3145 = reg3031;
              reg3146 = {forvar3111[(5'h19):(5'h11)],
                  (|(reg3015[(3'h4):(2'h3)] | reg2960[(4'h8):(2'h3)])),
                  ({(reg3046 + $unsigned(reg2965))} ?
                      {reg3145, (-((7'h49) & reg3059))} : reg3100)};
            end
        end
    end
  assign wire3147 = (reg3015[(2'h2):(1'h0)] ?
                        ((~&reg2962[(2'h3):(2'h2)]) ?
                            $unsigned((!$signed(wire1687))) : $signed({$unsigned(reg3071),
                                ((8'ha8) ?
                                    reg3065 : reg3022)})) : $unsigned((7'h40)));
  assign wire3148 = (($signed(reg3067[(2'h3):(1'h0)]) ?
                            reg3109 : (reg2967 ?
                                reg3020[(2'h3):(2'h3)] : (|$signed(reg3001)))) ?
                        $signed((+{(!reg3059)})) : (reg3041[(5'h14):(4'hd)] ?
                            $unsigned($signed({reg3085})) : (!((~^(7'h50)) ^ (^wire1694)))));
  always
    @(posedge clk) begin
      for (forvar3149 = (1'h0); (forvar3149 < (3'h6)); forvar3149 = (forvar3149 + (1'h1)))
        begin
          reg3150 <= reg3079[(2'h2):(1'h0)];
          for (forvar3151 = (1'h0); (forvar3151 < (3'h4)); forvar3151 = (forvar3151 + (1'h1)))
            begin
              reg3152 <= (~(^$signed($signed(wire3070[(1'h1):(1'h0)]))));
              reg3153 = reg2965[(4'h8):(1'h0)];
              reg3154 <= reg3022;
              reg3155 <= (~$unsigned({(reg3043[(5'h11):(4'h9)] >= (+(7'h47)))}));
              reg3156 = $signed(($unsigned($unsigned((|wire3148))) != $unsigned(wire1692)));
              reg3157 = wire3070[(3'h5):(1'h1)];
            end
          reg3158 = {reg3085, reg2991[(4'h8):(1'h0)]};
          if ($signed(reg3128))
            begin
              reg3159 = reg3059;
              reg3160 = $signed($signed((reg3158[(1'h1):(1'h0)] ?
                  ((wire3148 ^~ (7'h4e)) + reg3124[(2'h2):(1'h0)]) : (reg3063 ?
                      (reg3011 ? reg3155 : (7'h4d)) : reg3153))));
            end
          else
            begin
              reg3161 <= wire1688;
              reg3162 = ((~|$unsigned($signed(((8'hb5) ? reg3099 : reg3011)))) ?
                  reg3128[(2'h3):(2'h2)] : (8'hb4));
              reg3163 <= reg2972[(1'h1):(1'h1)];
              reg3164 = (~&$unsigned((~&$unsigned((&(7'h45))))));
              reg3165 <= ({reg3035[(4'hf):(4'h9)],
                      (((&reg3071) | wire1689) - (reg3073 < (|reg3156)))} ?
                  (~&wire2946) : reg3128[(1'h1):(1'h1)]);
              reg3166 <= $unsigned(wire3036[(4'he):(4'h8)]);
              reg3167 = $signed(($signed(reg2974[(5'h12):(4'h9)]) ?
                  reg2999 : $unsigned(reg3142)));
            end
          reg3168 <= {(|reg3011)};
          if ((((8'hb3) + ((|(reg3109 ?
                  reg2954 : reg3124)) <<< (reg3107 <= reg2965[(2'h2):(1'h1)]))) ?
              {reg2952[(1'h1):(1'h0)], (8'ha9), $signed(reg2965)} : reg3156))
            begin
              reg3169 <= (!wire3096);
              reg3170 <= $unsigned(reg2952[(2'h2):(2'h2)]);
              reg3171 = (8'ha6);
              reg3172 <= reg3043[(4'ha):(3'h6)];
              reg3173 <= reg3012;
            end
          else
            begin
              reg3171 = reg3135[(5'h13):(4'h8)];
              reg3174 = (&{(!((^reg2954) == (wire3096 && (8'hb1))))});
              reg3175 = reg3159[(1'h1):(1'h0)];
              reg3176 <= $signed((!reg3018));
              reg3177 = (|$unsigned($signed((-$unsigned(reg3107)))));
              reg3178 = ($signed(forvar3151) | {(-$unsigned((7'h49))),
                  (reg2949 != $signed((reg2962 ~^ reg3024))),
                  {wire1692[(2'h3):(2'h3)], $signed(reg2950[(5'h15):(4'ha)])}});
            end
        end
      if ((~|$unsigned($unsigned({(reg3015 ? reg3067 : (7'h40)), (~reg3001)}))))
        begin
          for (forvar3179 = (1'h0); (forvar3179 < (2'h2)); forvar3179 = (forvar3179 + (1'h1)))
            begin
              reg3180 <= $signed(wire2946[(1'h0):(1'h0)]);
              reg3181 = {((wire1692[(4'hd):(4'ha)] >> ((~reg3118) - reg3161)) ?
                      reg3172 : ($signed(((7'h41) ~^ reg3063)) ?
                          (|$unsigned(reg3022)) : ({reg3089,
                              (8'ha0),
                              reg2972} - reg3174))),
                  $unsigned({reg3180[(5'h15):(3'h5)]}),
                  $signed((~&(!reg3174)))};
              reg3182 = ((7'h41) + (((reg2962 ?
                      (wire1688 ?
                          reg3157 : reg3152) : (reg3158 || reg3098)) >>> $signed((reg3071 ?
                      wire1692 : wire1688))) ?
                  {($signed(reg2950) ? reg2949 : $unsigned(wire3147)),
                      ((^reg3165) ?
                          ((7'h47) ?
                              (8'ha7) : (7'h57)) : reg3173[(3'h6):(1'h0)])} : reg3075));
              reg3183 <= reg3165;
              reg3184 <= $unsigned(reg3175);
            end
          if (reg2954)
            begin
              reg3185 = reg2972;
              reg3186 = (!(+($unsigned((^~reg3152)) ?
                  (reg3128[(5'h11):(4'hf)] ?
                      reg2991[(5'h14):(3'h7)] : $signed(reg3172)) : reg2987[(4'h8):(3'h5)])));
              reg3187 = reg2962;
            end
          else
            begin
              reg3188 <= $signed((((!(|reg3116)) ^ $signed($signed(reg3059))) <= wire1694));
            end
          for (forvar3189 = (1'h0); (forvar3189 < (2'h3)); forvar3189 = (forvar3189 + (1'h1)))
            begin
              reg3190 <= reg3172;
              reg3191 = (!{reg3089[(2'h3):(1'h0)],
                  (|reg3031),
                  reg3098[(3'h6):(3'h6)]});
            end
          for (forvar3192 = (1'h0); (forvar3192 < (3'h5)); forvar3192 = (forvar3192 + (1'h1)))
            begin
              reg3193 = reg3004;
              reg3194 <= wire3148[(3'h4):(1'h1)];
              reg3195 = $unsigned(($signed((8'ha3)) ?
                  ({(reg2975 ? reg2991 : (8'hac)), $unsigned(reg3177)} ?
                      reg3191 : (~&$unsigned(reg3067))) : $unsigned($unsigned($signed((8'hbb))))));
            end
          for (forvar3196 = (1'h0); (forvar3196 < (1'h1)); forvar3196 = (forvar3196 + (1'h1)))
            begin
              reg3197 = $unsigned(((~|reg2993[(5'h10):(3'h6)]) <= {(~&{reg3047,
                      (8'hb3),
                      forvar3189}),
                  (+reg3172[(2'h2):(2'h2)])}));
            end
          reg3198 <= ($unsigned(reg2983[(4'hb):(1'h0)]) ?
              wire1690 : $unsigned(wire1692));
          for (forvar3199 = (1'h0); (forvar3199 < (3'h6)); forvar3199 = (forvar3199 + (1'h1)))
            begin
              reg3200 <= $signed(reg3038);
              reg3201 = $unsigned($unsigned(reg2955[(5'h10):(3'h4)]));
              reg3202 = $signed((|(+{reg3190[(1'h0):(1'h0)],
                  (reg3002 >> reg3190),
                  $signed(reg3080)})));
            end
        end
      else
        begin
          for (forvar3179 = (1'h0); (forvar3179 < (1'h1)); forvar3179 = (forvar3179 + (1'h1)))
            begin
              reg3180 <= $signed($unsigned((((reg2981 ? (8'hbd) : forvar3189) ?
                      ((8'hb6) ? reg3059 : reg3009) : reg3156) ?
                  reg3046 : {(!reg3080)})));
              reg3181 = {$unsigned($signed((reg3158[(2'h3):(2'h2)] || $unsigned(reg3046))))};
              reg3182 = (wire3148 > reg3079[(4'hc):(4'ha)]);
              reg3185 = ((-($unsigned(reg3067) ?
                      ($signed(forvar3179) ?
                          $signed(reg3200) : forvar3192[(2'h2):(2'h2)]) : (+$unsigned(reg2960)))) ?
                  (($unsigned(wire3036) != {(-(8'hb5))}) ?
                      $signed((reg3132[(2'h2):(1'h0)] && (reg3059 != reg3065))) : $signed((^reg3020[(3'h5):(1'h1)]))) : wire1694[(5'h17):(5'h12)]);
            end
          reg3188 <= (~|(({(+reg3018), (~|reg3023)} ?
                  $signed(reg3011[(5'h11):(3'h4)]) : wire3147) ?
              reg3011 : reg3002));
          if ((&$signed(((^~reg2951[(3'h6):(3'h4)]) ?
              ((reg3024 ? reg3079 : wire1689) ?
                  reg3023 : ((8'h9e) ?
                      (8'hbf) : reg2999)) : reg3195[(1'h1):(1'h0)]))))
            begin
              reg3189 <= ($signed(($signed(reg3156[(4'hd):(2'h2)]) ?
                  $unsigned($unsigned(reg3182)) : $unsigned((7'h43)))) >> reg3015);
              reg3191 = ($unsigned(((~(reg3182 ? forvar3189 : (7'h4f))) ?
                      reg3165 : (((8'hb5) + wire1692) * $unsigned(reg3165)))) ?
                  reg3135 : $unsigned(wire3147[(2'h3):(2'h2)]));
              reg3192 <= (&reg2951);
              reg3193 = reg3027;
              reg3194 <= (8'ha7);
              reg3195 = (((~^$signed($unsigned(reg2997))) < ($unsigned($signed(reg3191)) ?
                  reg3162 : {(reg3122 | (8'ha6))})) - $unsigned(reg3003[(3'h5):(2'h3)]));
            end
          else
            begin
              reg3189 <= reg3172;
              reg3190 <= reg3156;
              reg3192 <= ((~|reg3032[(3'h4):(2'h2)]) ?
                  reg2969 : $signed(((-$signed(reg3178)) ?
                      $signed({reg2960, (7'h42), (7'h4f)}) : {reg3189})));
              reg3193 = {reg3193,
                  {wire1691[(1'h0):(1'h0)],
                      (~^reg3180),
                      ((|reg3198) ~^ $unsigned((reg3011 ?
                          wire3036 : (7'h57))))},
                  {reg3102,
                      (($signed(reg2955) ?
                          $unsigned(forvar3199) : (8'h9e)) <= $unsigned((reg3142 == reg3187)))}};
              reg3195 = $unsigned(reg3093);
              reg3196 = (($signed(forvar3189) ?
                  reg3164[(3'h4):(2'h3)] : $unsigned((!(^~reg3085)))) <<< ((~reg3181[(4'hd):(3'h7)]) ?
                  {forvar3199[(1'h0):(1'h0)],
                      $unsigned(((7'h42) ? reg3093 : (8'ha8))),
                      (reg2967 ?
                          $signed(reg3173) : $unsigned(reg2949))} : (^reg3020)));
              reg3198 <= forvar3192;
            end
          reg3199 = wire1694;
          reg3201 = {(reg3095[(1'h1):(1'h0)] ^ $unsigned({reg3002})),
              $unsigned((($signed(reg3009) && (reg3168 ? reg3201 : reg3041)) ?
                  wire1692 : $signed($signed(reg3131))))};
          reg3202 = (&{($signed($unsigned(reg3199)) >= {wire1693[(5'h12):(3'h7)],
                  reg3182,
                  (reg3075 ? wire2948 : (7'h48))}),
              {reg2969[(3'h5):(3'h5)], (^(~&reg3135))}});
        end
      reg3203 = $unsigned(reg3200[(5'h11):(4'hb)]);
      for (forvar3204 = (1'h0); (forvar3204 < (1'h0)); forvar3204 = (forvar3204 + (1'h1)))
        begin
          reg3205 <= reg3002;
          if ($signed({({(reg2991 ? wire3148 : (8'h9f))} & (~&(&reg3031))),
              (^({reg3099} ? reg2950[(4'hb):(3'h7)] : (~|forvar3204)))}))
            begin
              reg3206 <= (8'hb2);
              reg3207 = reg3132[(3'h5):(3'h5)];
            end
          else
            begin
              reg3206 <= $signed((reg3038 == ($signed((8'ha6)) <<< (^$signed(reg3063)))));
              reg3207 = $unsigned((($signed($unsigned((8'ha9))) ?
                  $unsigned($unsigned(reg3033)) : $unsigned($signed(reg3107))) << reg3173));
            end
        end
      if ($unsigned($unsigned($unsigned((~^reg3144[(5'h18):(4'ha)])))))
        begin
          if ({$signed($signed($unsigned($unsigned((8'hb0)))))})
            begin
              reg3208 <= (reg3015[(2'h3):(1'h1)] ?
                  $signed((^$signed((reg3079 ?
                      reg3135 : reg3207)))) : (reg2950[(2'h2):(1'h0)] | $signed(reg3106)));
            end
          else
            begin
              reg3209 = $unsigned($unsigned(reg3058));
              reg3210 = (~(|$signed({{reg3022, reg3144, reg3113},
                  $unsigned(reg3001)})));
            end
          reg3211 = $signed($signed((wire3147 ?
              $unsigned($signed((8'hbb))) : $signed(((8'haf) ?
                  reg3144 : reg3170)))));
          reg3212 <= $signed(((-(^$unsigned(reg3180))) ?
              ($unsigned({(8'haa),
                  reg3033,
                  reg2980}) != $unsigned((7'h58))) : reg3181[(3'h6):(2'h2)]));
          for (forvar3213 = (1'h0); (forvar3213 < (2'h3)); forvar3213 = (forvar3213 + (1'h1)))
            begin
              reg3214 = $signed(reg2950);
              reg3215 <= ((^~{((reg3165 ^ reg3089) >= $signed(reg3142)),
                  ((reg3101 + (7'h4a)) >> (-reg3063)),
                  $unsigned(reg3162[(4'h9):(2'h2)])}) || $signed((reg3198 ?
                  ({(8'ha8), reg2954} != (reg3189 || reg3185)) : reg3164)));
              reg3216 = reg3116[(4'hd):(4'h9)];
              reg3217 = (((reg3047 ?
                      reg3158 : ((&forvar3199) ^~ $unsigned(reg3172))) ?
                  $signed({(!reg3168),
                      reg3142[(3'h6):(1'h0)],
                      $unsigned(reg2993)}) : ($signed($unsigned((8'ha5))) ?
                      reg3003 : (reg2991[(4'hc):(1'h0)] ?
                          (reg3063 ^ (8'ha3)) : ((7'h44) != reg3012)))) ^~ {(~|(reg3164[(2'h2):(2'h2)] ?
                      wire1689 : reg3113)),
                  {{$unsigned(reg2952), (&reg3109)}, (^(|reg3020))},
                  $signed((^~reg3004))});
              reg3218 <= (reg3156 << ((reg3135 ?
                      reg2997[(4'h9):(3'h7)] : {(reg3172 ? reg3071 : reg2991),
                          (|reg3206)}) ?
                  $unsigned(($signed(reg3004) ?
                      {forvar3192,
                          reg3041} : $unsigned(reg3024))) : $signed(((!reg3027) ?
                      forvar3189 : (&reg2983)))));
              reg3219 = ((^$unsigned(((reg3198 ? forvar3179 : reg2962) ?
                      $signed(reg3185) : ((7'h54) ? (7'h57) : reg3031)))) ?
                  $unsigned((reg2991 + {reg3206})) : wire1689);
              reg3220 <= (reg3095 ?
                  (reg3003[(2'h2):(1'h0)] >= (8'had)) : reg3175);
            end
        end
      else
        begin
          if ((reg2993 ?
              (reg3018[(5'h1c):(4'h9)] * (((8'hb3) ?
                      reg3046[(5'h13):(1'h1)] : reg3218[(5'h1b):(5'h1a)]) ?
                  reg3031 : forvar3151[(4'hb):(4'h9)])) : $unsigned(reg3165)))
            begin
              reg3208 <= (((((reg3030 ?
                          reg3190 : (8'hb7)) < (reg3216 ~^ reg3005)) ^ ((reg2999 | (8'hab)) ?
                          $unsigned(reg3183) : $signed(reg3201))) ?
                      reg3164[(2'h2):(1'h1)] : (&{{forvar3213,
                              (7'h40),
                              reg3134},
                          reg3131,
                          $unsigned(reg3085)})) ?
                  reg3067[(2'h3):(2'h2)] : reg3189);
              reg3212 <= (reg3184 ?
                  ((~|(~|(reg3160 ?
                      reg3102 : reg2991))) * reg3164) : ($unsigned($unsigned(reg3032)) << (~^(reg3005[(3'h6):(1'h1)] || (reg3035 ^ reg3071)))));
              reg3213 = ((~$unsigned((~|(reg3144 ?
                  reg3219 : reg3220)))) ~^ (($signed((reg3098 ?
                          reg3041 : wire3148)) ?
                      ($signed(reg3197) << $signed(reg3197)) : reg3065) ?
                  reg2999 : {reg3026}));
              reg3214 = {(+({(wire1687 ? forvar3149 : (8'h9f)),
                          reg3177[(5'h1c):(5'h10)]} ?
                      (&{reg3184, reg3059, reg3003}) : (|((8'ha0) ?
                          reg2975 : reg3172)))),
                  reg3177[(5'h17):(4'hb)]};
              reg3215 <= reg3116;
            end
          else
            begin
              reg3209 = {((&reg3024) ?
                      reg3197 : ((|$unsigned(reg3214)) ?
                          ($signed(reg2950) ?
                              (reg3215 == reg3160) : (&forvar3189)) : $unsigned({reg3213,
                              reg3004}))),
                  $unsigned(reg3160[(2'h2):(1'h0)])};
              reg3212 <= $signed($unsigned(reg3023[(5'h13):(3'h6)]));
              reg3215 <= {((+$signed(reg2980)) ?
                      (^~reg3208[(1'h1):(1'h0)]) : reg3192),
                  ((-(reg3030 + $signed(wire1692))) ?
                      {((+reg2955) - $signed(reg3186)),
                          reg3162} : $signed(((reg2972 * reg3198) ~^ wire2948)))};
              reg3216 = (reg3003[(5'h11):(4'hd)] ?
                  $unsigned((&reg3206[(4'h9):(1'h1)])) : ((((reg3157 ?
                          reg3208 : reg3201) >= reg3093) - $signed(reg3154[(2'h3):(2'h3)])) ?
                      $unsigned((7'h54)) : $unsigned((&(|(7'h49))))));
              reg3218 <= (!$unsigned(reg3131));
              reg3220 <= $unsigned(($signed(reg3203) < reg3003));
              reg3221 = $unsigned(((~{reg2962, $unsigned(reg3073)}) ?
                  reg3113[(4'ha):(4'ha)] : (~$unsigned($signed(reg2969)))));
            end
          if (reg3116)
            begin
              reg3222 <= ($unsigned(((^(reg3153 || (8'ha1))) << ($unsigned(reg3192) ^ (reg3187 <= reg3173)))) ?
                  $signed($signed(($unsigned((8'h9e)) ?
                      $signed((8'hb2)) : (reg2991 <= (8'ha9))))) : {(reg3023 ?
                          (reg3063[(3'h7):(2'h2)] ?
                              $signed(wire1689) : $signed(reg2954)) : ((reg3102 || reg3176) ?
                              $signed(reg2972) : (reg3027 ?
                                  (8'ha6) : wire1692)))});
              reg3223 = (&(^reg3184[(1'h0):(1'h0)]));
              reg3224 = ({forvar3189[(1'h1):(1'h0)],
                      $unsigned($signed((~&reg3134))),
                      (reg2972[(2'h2):(1'h1)] ?
                          ($unsigned(reg3002) ?
                              $unsigned(reg3003) : (wire1687 && reg2991)) : ((reg3159 || reg3002) * $unsigned(reg3073)))} ?
                  (~|forvar3149) : reg3093[(2'h2):(2'h2)]);
              reg3225 = reg2960;
              reg3226 <= (reg3122 ?
                  ((~&(~(reg3188 ? reg3214 : (7'h55)))) ?
                      (^~reg3065[(3'h6):(3'h5)]) : reg3033) : wire3070[(3'h7):(3'h6)]);
              reg3227 = $unsigned((~($unsigned((reg2962 & reg3038)) >= (reg2981[(4'h9):(3'h7)] & (-reg3186)))));
            end
          else
            begin
              reg3223 = reg3075[(4'hb):(3'h7)];
              reg3224 = ($unsigned($unsigned(({reg3160} + ((8'h9f) ?
                      reg3170 : reg3043)))) ?
                  $signed((^~$signed(((7'h4f) << wire1689)))) : $unsigned(reg3039[(3'h4):(3'h4)]));
              reg3225 = (((({reg2991} == reg3196[(4'h8):(3'h5)]) ?
                      {(reg3221 != reg3203)} : (~|reg3196)) & (8'hbb)) ?
                  ($unsigned(reg3208) >>> reg3067) : wire2948);
              reg3227 = (~(!reg3154[(2'h3):(1'h0)]));
              reg3228 <= ((reg3223 >>> reg3046) >= reg2993[(3'h7):(1'h0)]);
              reg3229 = ((8'h9d) ?
                  reg3184[(1'h0):(1'h0)] : ({((reg3167 >> reg3075) | $signed(reg3215)),
                      reg3159,
                      reg3200[(5'h13):(3'h7)]} + $unsigned($signed($unsigned((7'h4e))))));
            end
          reg3230 <= $signed(reg3212[(4'h8):(2'h3)]);
          reg3231 = $unsigned((~|$unsigned(reg3093[(4'hb):(3'h5)])));
        end
      reg3232 <= reg3215;
      for (forvar3233 = (1'h0); (forvar3233 < (2'h3)); forvar3233 = (forvar3233 + (1'h1)))
        begin
          reg3234 <= reg3122;
          if (reg3043[(4'hb):(3'h5)])
            begin
              reg3235 <= reg3198[(4'hb):(4'h9)];
              reg3236 <= reg3218[(5'h1d):(4'ha)];
              reg3237 <= forvar3233[(4'hf):(1'h0)];
              reg3238 <= (+{(($unsigned(reg2987) ?
                          reg2960[(4'hc):(4'h9)] : $signed(reg3181)) ?
                      $unsigned((~|reg3227)) : $signed((reg3002 ?
                          (7'h40) : reg3109))),
                  (($unsigned(reg3026) ? (~&reg3187) : (reg3184 >>> (8'hb5))) ?
                      $unsigned($signed(reg3159)) : wire3147[(1'h1):(1'h0)]),
                  (~|(reg3193 >= reg3162[(1'h0):(1'h0)]))});
              reg3239 <= {(~&(-((reg3159 > reg3200) ^~ $unsigned(reg3039)))),
                  $signed(reg3116[(3'h6):(1'h1)])};
              reg3240 <= $signed($signed({reg2981[(1'h1):(1'h0)],
                  $signed((reg3107 + reg3199)),
                  wire3148}));
            end
          else
            begin
              reg3235 <= (!($unsigned($unsigned($unsigned(reg2981))) != reg3223));
              reg3241 = (^~((reg3178 ?
                      ({(8'haf),
                          (8'h9e),
                          reg3128} < (reg3195 >= reg3161)) : ($unsigned(reg3228) ?
                          $unsigned(reg2987) : ((8'hbf) <<< reg3236))) ?
                  reg3004 : {((reg3182 ? reg3109 : reg2967) ?
                          reg3218[(2'h2):(1'h0)] : reg3046[(4'he):(2'h3)]),
                      $unsigned((+reg3067))}));
              reg3242 = reg3116[(4'hb):(3'h5)];
              reg3243 <= reg2954;
              reg3244 <= reg3166;
            end
          if (forvar3151)
            begin
              reg3245 = $unsigned((-{(reg3167 >= $unsigned(reg3039)),
                  (~&$signed(reg3221)),
                  $signed((reg3031 ? reg3209 : reg3198))}));
              reg3246 <= $unsigned(((wire3070 * (-reg3226[(3'h4):(2'h3)])) ?
                  reg2950 : ($unsigned((reg3101 ?
                      forvar3199 : reg3046)) ~^ ($signed(reg3216) ?
                      (wire1694 >> reg3035) : ((8'hbb) | reg3101)))));
            end
          else
            begin
              reg3245 = $signed($signed(({(reg3169 ? reg3217 : reg3005)} ?
                  (reg3155 ? {reg3059} : reg2974) : ((reg2951 ?
                          reg3238 : reg3093) ?
                      (8'ha5) : (wire1692 >= reg3181)))));
              reg3247 = $signed($unsigned((7'h4e)));
              reg3248 <= $unsigned(reg3234[(2'h2):(1'h1)]);
              reg3249 <= reg3214[(2'h2):(2'h2)];
              reg3250 <= reg3131;
              reg3251 = $signed($unsigned($unsigned({(+(7'h49)),
                  wire1689[(5'h14):(4'hc)],
                  (reg3182 ? reg3217 : (8'hb3))})));
            end
          reg3252 = (!reg3144);
          if ((reg3210 ?
              $unsigned($unsigned((reg3176 ?
                  reg3160 : $signed(wire1693)))) : reg3131[(3'h5):(2'h3)]))
            begin
              reg3253 <= reg3209;
              reg3254 = (forvar3149[(4'hd):(4'hc)] ?
                  reg3032[(5'h16):(2'h2)] : ($unsigned($signed($unsigned(reg3018))) ?
                      ((-$signed(wire2946)) ^~ $unsigned(reg3225[(3'h4):(3'h4)])) : (($unsigned(reg3213) ?
                              ((7'h40) ? reg3122 : reg3032) : (^reg3022)) ?
                          reg3162 : $signed((reg3150 + reg2987)))));
              reg3255 = $signed($unsigned($signed({reg2952,
                  reg3165[(4'he):(3'h7)]})));
              reg3256 = {$signed(($unsigned(((8'hbf) ^ reg3073)) | $signed(forvar3192[(3'h7):(3'h4)]))),
                  $unsigned(reg2962[(4'hf):(3'h5)]),
                  forvar3179};
              reg3257 <= {(&$unsigned($unsigned(reg3256[(5'h17):(5'h15)])))};
              reg3258 <= (((reg3026[(1'h1):(1'h1)] ?
                      (~^(reg3065 ?
                          reg3203 : reg3196)) : $unsigned(reg3222[(4'hb):(4'ha)])) ?
                  (reg3221[(2'h3):(2'h3)] <= $unsigned($signed((8'hb1)))) : ((|reg3160[(2'h2):(1'h0)]) >> (7'h44))) == reg3213);
            end
          else
            begin
              reg3253 <= ((($signed(reg3217[(4'ha):(3'h4)]) ?
                          (reg3196[(4'he):(4'hc)] ~^ (forvar3213 != reg3217)) : $unsigned((reg3244 ?
                              reg3198 : reg3200))) ?
                      reg3164[(3'h7):(3'h7)] : $signed($signed($unsigned(reg3171)))) ?
                  (({(reg3094 - reg3248)} ?
                      reg3157[(3'h6):(3'h6)] : (~(reg2981 ?
                          reg3219 : reg3219))) >>> ($signed(reg3237) != ((reg3230 ?
                      (8'ha4) : reg3198) <<< reg3009))) : (reg3085 == $unsigned(((&(8'h9d)) < reg3230))));
              reg3254 = (~^(^$unsigned({reg3124[(3'h4):(2'h2)],
                  reg3038,
                  (8'hb4)})));
              reg3255 = (-((~|wire1692[(3'h6):(3'h6)]) | $signed($unsigned(reg3198[(4'h9):(1'h1)]))));
            end
          if ((~&((!$unsigned($unsigned((7'h42)))) != (^$unsigned($unsigned(reg3009))))))
            begin
              reg3259 = $unsigned(reg3124);
              reg3260 = (7'h4a);
              reg3261 <= reg3199;
              reg3262 <= reg3261[(3'h6):(2'h3)];
              reg3263 = (~reg3255[(1'h1):(1'h0)]);
              reg3264 = ($signed((((reg2999 && reg3190) ?
                      $unsigned(reg3099) : $signed(reg3154)) | reg2949[(4'he):(4'he)])) ?
                  (reg3033[(2'h2):(1'h0)] ?
                      $signed({$unsigned((8'hbc)),
                          (reg3181 * reg3124)}) : $unsigned(reg3003)) : wire3147);
              reg3265 <= $signed((~$unsigned(reg3180[(1'h1):(1'h1)])));
            end
          else
            begin
              reg3259 = {reg3213};
              reg3261 <= $signed((reg3232[(3'h5):(2'h2)] ?
                  (~^(8'h9f)) : reg2952[(3'h5):(1'h0)]));
              reg3263 = reg3187[(5'h14):(5'h10)];
              reg3265 <= ({$unsigned(({wire1691,
                      reg2987} ^ $unsigned(reg3160))),
                  ($unsigned((reg3095 ? reg3183 : reg3220)) ?
                      ((reg3158 ~^ reg2983) ?
                          reg2997[(5'h1a):(3'h6)] : (reg3206 | reg3228)) : reg3175[(4'h9):(2'h2)])} || (8'h9e));
              reg3266 <= ($signed({(((8'ha2) - reg2997) != (reg3187 ?
                          reg3134 : reg3099))}) ?
                  reg3099[(2'h2):(2'h2)] : wire3096[(1'h1):(1'h1)]);
              reg3267 <= (({reg3153} - (((reg3095 ? (7'h52) : reg3221) ?
                      $signed(reg3041) : (reg3202 >= reg3116)) ?
                  $signed($unsigned((7'h46))) : $signed(reg3207[(2'h3):(1'h0)]))) ~^ ($unsigned(reg3001[(1'h1):(1'h1)]) ?
                  ($signed($signed((7'h4a))) >= reg3047) : (8'h9f)));
            end
        end
    end
  assign wire3268 = (8'ha1);
  always
    @(posedge clk) begin
      for (forvar3269 = (1'h0); (forvar3269 < (1'h1)); forvar3269 = (forvar3269 + (1'h1)))
        begin
          reg3270 = wire2948;
        end
      for (forvar3271 = (1'h0); (forvar3271 < (1'h1)); forvar3271 = (forvar3271 + (1'h1)))
        begin
          for (forvar3272 = (1'h0); (forvar3272 < (2'h2)); forvar3272 = (forvar3272 + (1'h1)))
            begin
              reg3273 <= $unsigned({wire1689[(5'h12):(4'hf)],
                  ($signed($unsigned((7'h43))) ?
                      $unsigned($signed(reg3266)) : ($signed(reg3212) * {(8'ha6),
                          reg3063}))});
            end
          if (($unsigned($signed(reg3035[(4'h8):(3'h7)])) + (^reg3142[(4'h8):(3'h7)])))
            begin
              reg3274 = wire3070[(1'h0):(1'h0)];
              reg3275 = (7'h47);
              reg3276 = reg3107[(3'h4):(2'h3)];
              reg3277 <= wire1687;
              reg3278 = (((($unsigned(reg3027) ?
                  (&(8'h9c)) : reg3080[(1'h0):(1'h0)]) ~^ $signed(reg3094[(1'h1):(1'h1)])) > (-$signed(((8'hab) ?
                  reg3020 : wire1692)))) >= (|$unsigned((~^reg3270))));
              reg3279 = (reg3270[(4'hf):(4'h8)] ?
                  reg3277[(3'h6):(3'h5)] : $signed(({(reg3226 ?
                          reg3232 : wire1689),
                      reg3095[(3'h5):(1'h0)],
                      $unsigned(reg3190)} >>> (reg3173 ?
                      $unsigned(reg3165) : (reg3270 ? reg3237 : reg3081)))));
              reg3280 <= reg3085;
            end
          else
            begin
              reg3274 = $signed($unsigned(reg3215[(3'h6):(2'h2)]));
            end
        end
      for (forvar3281 = (1'h0); (forvar3281 < (2'h3)); forvar3281 = (forvar3281 + (1'h1)))
        begin
          for (forvar3282 = (1'h0); (forvar3282 < (2'h2)); forvar3282 = (forvar3282 + (1'h1)))
            begin
              reg3283 = $signed($unsigned($unsigned($unsigned((^~reg3101)))));
              reg3284 <= reg3230[(1'h0):(1'h0)];
              reg3285 = (7'h44);
            end
          if ((reg3058 ? reg3220[(1'h1):(1'h0)] : wire1688[(5'h18):(4'hb)]))
            begin
              reg3286 = reg3098[(3'h6):(3'h5)];
              reg3287 = {$signed(($signed($signed(reg3279)) <<< (+$signed(reg3237)))),
                  ($signed($unsigned($unsigned(reg3063))) ?
                      (~|(reg3238 ^~ (reg3113 ~^ reg3258))) : reg3170),
                  {$unsigned((!{reg2974, reg3011}))}};
              reg3288 <= ($unsigned($unsigned((^(|reg3189)))) * (^(~reg3198[(4'hc):(4'hc)])));
              reg3289 = ({wire3148[(1'h1):(1'h1)]} << reg3169[(4'h9):(3'h6)]);
            end
          else
            begin
              reg3288 <= $unsigned(reg3155[(5'h1c):(5'h17)]);
            end
        end
      reg3290 = {($unsigned(($signed(reg3194) ?
                  reg3265 : (reg3024 && reg3059))) ?
              (reg3004 ?
                  $signed((~&reg3003)) : ($unsigned(wire1693) | {(7'h51),
                      (8'hbd)})) : $unsigned($unsigned(forvar3272[(2'h2):(2'h2)]))),
          (7'h47)};
      for (forvar3291 = (1'h0); (forvar3291 < (3'h6)); forvar3291 = (forvar3291 + (1'h1)))
        begin
          if ($signed((~|{($unsigned(reg3075) ?
                  $signed(reg3244) : {wire1690, reg2983}),
              ((7'h4a) < $signed(reg3258)),
              (reg3161[(5'h12):(4'he)] || (~&reg3243))})))
            begin
              reg3292 = ($signed((|($signed(reg3257) ?
                  (-reg2949) : (reg3089 ^ reg3023)))) <= reg3003);
              reg3293 <= reg3283[(4'h8):(2'h3)];
              reg3294 = reg2975[(2'h3):(1'h1)];
              reg3295 <= reg3262;
            end
          else
            begin
              reg3293 <= forvar3269;
              reg3295 <= (wire1689[(4'hf):(1'h1)] < (^~$unsigned((^~(reg2967 ?
                  (7'h41) : reg2974)))));
              reg3296 <= reg3235;
              reg3297 <= (reg3168 ?
                  reg3284[(3'h4):(3'h4)] : $unsigned({$signed((reg3188 * forvar3281)),
                      reg3079}));
              reg3298 <= reg3065[(3'h4):(2'h2)];
              reg3299 = {reg3198};
            end
          reg3300 <= reg3077[(1'h0):(1'h0)];
        end
      reg3301 = {reg3093,
          (+(((reg3118 < reg3297) * $signed(reg3228)) ?
              reg3011 : $unsigned({reg2987})))};
    end
  always
    @(posedge clk) begin
      if ((reg3253[(1'h1):(1'h1)] ?
          reg3266 : {$signed((+(reg3188 ? wire2948 : reg3102))), reg3189}))
        begin
          for (forvar3302 = (1'h0); (forvar3302 < (3'h4)); forvar3302 = (forvar3302 + (1'h1)))
            begin
              reg3303 = wire1692;
              reg3304 <= ($unsigned(($unsigned((&wire1694)) ?
                  ($signed(reg3002) ?
                      reg2981 : (^reg3220)) : {$unsigned(wire3096),
                      $signed((8'hac)),
                      (reg3190 ~^ reg3176)})) >= wire1693[(2'h2):(1'h0)]);
              reg3305 = {$unsigned((reg3248 >= $unsigned((reg2967 ^~ (7'h44)))))};
              reg3306 = $signed(reg3173[(5'h10):(4'hf)]);
            end
          reg3307 = reg3116[(4'h9):(1'h0)];
          reg3308 <= $unsigned(($unsigned(reg3011[(3'h7):(3'h6)]) >= ({{reg3295},
                  (reg3198 ^ reg2952),
                  (|(8'hbd))} ?
              reg2993 : reg3243[(4'h9):(1'h1)])));
        end
      else
        begin
          if ($signed(reg3305))
            begin
              reg3302 = (|reg2952);
              reg3303 = reg3089;
            end
          else
            begin
              reg3304 <= reg3298[(3'h7):(3'h4)];
              reg3305 = wire3147[(5'h10):(5'h10)];
              reg3308 <= $unsigned(($signed((~|$unsigned(reg3085))) ?
                  $unsigned($signed((reg3192 ^~ reg3297))) : (|(8'hb6))));
            end
          if ({(reg3306[(2'h2):(2'h2)] ^~ (reg3238[(3'h5):(3'h5)] == (|(+reg3261))))})
            begin
              reg3309 <= $signed($signed(($unsigned($signed((8'hbd))) ?
                  {reg3079[(4'ha):(3'h6)],
                      $signed(reg3009),
                      (reg3093 >> (7'h43))} : $unsigned((reg3183 || (7'h4d))))));
              reg3310 <= (+(~(-reg3257[(4'hd):(2'h3)])));
              reg3311 <= ($signed(reg3277) >= ((reg3298 || (!(&(8'hba)))) & $signed($unsigned($signed(wire2946)))));
              reg3312 <= reg3124[(3'h4):(1'h1)];
              reg3313 = reg3200[(3'h5):(3'h4)];
            end
          else
            begin
              reg3313 = {reg3080, reg3236[(4'h9):(1'h0)]};
              reg3314 = $unsigned(reg3168[(5'h14):(2'h3)]);
              reg3315 = $signed(reg3047);
              reg3316 <= reg3280;
              reg3317 = (+$unsigned(reg3023[(5'h12):(4'h9)]));
            end
        end
      for (forvar3318 = (1'h0); (forvar3318 < (2'h3)); forvar3318 = (forvar3318 + (1'h1)))
        begin
          reg3319 = {(reg3244 ?
                  (+(8'ha6)) : {$signed((reg3132 ? reg2991 : (8'ha8)))})};
          reg3320 = (-forvar3318);
          reg3321 = {reg3296[(4'h9):(4'h9)],
              (~|($unsigned((~&reg3059)) | ({reg3047, reg3073, reg3047} ?
                  (!forvar3318) : $signed((8'hab))))),
              reg3169};
          if ((reg3022 ? $unsigned($unsigned((~|(-reg3118)))) : reg3035))
            begin
              reg3322 <= (8'hbf);
              reg3323 <= $signed((reg3288[(5'h10):(1'h0)] + (8'hac)));
              reg3324 <= {(^wire1689[(4'h8):(3'h7)]),
                  (($signed((~wire1693)) ?
                      $unsigned(((8'hb2) & reg3128)) : reg3306[(1'h0):(1'h0)]) - reg3046[(3'h6):(3'h4)])};
              reg3325 = $unsigned(reg2952[(3'h5):(3'h5)]);
              reg3326 = $unsigned(reg2997);
              reg3327 = $signed(reg3300);
            end
          else
            begin
              reg3325 = reg3249[(4'hb):(3'h4)];
              reg3326 = (^reg3249);
            end
          reg3328 = reg3099[(5'h1f):(5'h1f)];
          reg3329 = reg2960[(3'h6):(2'h2)];
        end
      reg3330 = wire1693;
      if (((reg3168[(2'h3):(1'h0)] ?
              ((~&(reg3183 ^ reg3089)) ?
                  reg3200 : $unsigned((reg3001 ?
                      reg3041 : reg3248))) : reg3073) ?
          reg3327[(2'h2):(1'h1)] : reg3011))
        begin
          if ((({$unsigned(((8'ha0) ^~ (8'hb3))),
                  (!(reg3079 ? reg2997 : (8'hb0))),
                  reg2965} ?
              (~($signed(reg3093) ?
                  {wire1692} : (|reg3015))) : ($unsigned(reg3228[(5'h17):(4'h9)]) ?
                  reg3150 : ($signed(reg3297) ?
                      $signed(reg3304) : $unsigned(forvar3302)))) * reg3288[(1'h0):(1'h0)]))
            begin
              reg3331 = (({{(&reg3298),
                          (reg3128 ? reg3329 : reg3033),
                          ((8'ha0) && reg3063)}} ?
                  reg2975 : $unsigned(reg3226[(4'h9):(3'h7)])) || reg3240);
            end
          else
            begin
              reg3331 = $signed({reg3319});
              reg3332 <= $unsigned((reg3144[(5'h16):(5'h16)] << {((7'h4f) ?
                      (7'h48) : reg3110[(2'h2):(1'h0)]),
                  $unsigned($unsigned(reg3293))}));
              reg3333 <= ($unsigned($signed(((reg3107 ?
                  reg2949 : reg3280) && $signed(reg3026)))) && (&($signed((reg3208 - reg2950)) > reg3122[(3'h5):(3'h5)])));
              reg3334 <= {reg3004[(3'h4):(1'h0)]};
              reg3335 = (~^(7'h48));
              reg3336 = (&(^~($signed({reg3099, reg3326, (8'hbd)}) ?
                  $signed($signed(reg3150)) : reg3246[(1'h1):(1'h0)])));
              reg3337 <= $unsigned($unsigned(({(reg3331 + reg3208),
                  $unsigned((8'hb6))} && reg3192[(5'h1b):(5'h17)])));
            end
          reg3338 <= $unsigned($signed((8'hb4)));
          for (forvar3339 = (1'h0); (forvar3339 < (1'h1)); forvar3339 = (forvar3339 + (1'h1)))
            begin
              reg3340 <= (($signed(($unsigned((8'hbc)) ?
                          (reg3303 ? reg3047 : reg3063) : (7'h51))) ?
                      (({reg3240, reg2975} != ((8'ha1) ?
                          wire1690 : reg3277)) + $unsigned(wire1692)) : reg3331[(3'h4):(2'h2)]) ?
                  (&$unsigned(({wire3148} ^~ reg3122))) : $unsigned(($signed({reg3300,
                          reg3295,
                          reg3244}) ?
                      ($unsigned(reg3180) ?
                          {reg3089} : {reg3155,
                              reg2955,
                              reg3198}) : $unsigned((reg3321 != (8'ha3))))));
              reg3341 <= (((!(~&(~^(8'hac)))) ?
                  $signed((~|reg3280[(5'h19):(5'h16)])) : (~^reg3009)) < (+((+{reg3310,
                      reg3043,
                      reg3323}) ?
                  $unsigned(reg3314[(4'h8):(3'h4)]) : reg3218)));
              reg3342 = $unsigned($signed({(((8'hac) <= reg3020) ^ (~|forvar3302)),
                  ((8'hbf) ? (reg3266 * (7'h50)) : reg3324)}));
              reg3343 <= {(^~({(~&(8'hb4)), {reg3238}, $unsigned(reg3152)} ?
                      reg3020 : $signed((+reg3067)))),
                  {(^{$unsigned(reg3041), $signed((7'h47))})}};
              reg3344 <= reg3038;
              reg3345 <= (&{({(reg3032 && reg3165)} - reg3320),
                  $signed($signed($unsigned(reg3248))),
                  ($unsigned({reg3266}) < reg3184)});
              reg3346 <= reg3001[(1'h1):(1'h1)];
            end
          reg3347 = $unsigned(reg3095);
          reg3348 <= {(-(7'h58)), reg3188};
          if (reg2981)
            begin
              reg3349 <= (+reg3288);
              reg3350 = reg3116;
              reg3351 <= {(&$signed(({wire3268} != $unsigned(reg2965)))),
                  ($signed($signed(reg3319[(2'h2):(1'h0)])) ?
                      (reg3302[(2'h2):(1'h1)] >> ((reg3106 ?
                              reg3320 : reg2950) ?
                          reg2972[(1'h1):(1'h0)] : reg3273)) : $signed(reg3324[(5'h17):(2'h3)])),
                  (^reg3240)};
              reg3352 = $unsigned($unsigned((reg3067[(3'h5):(3'h5)] ?
                  $signed($unsigned(reg2983)) : reg2955)));
              reg3353 = reg3101[(2'h2):(1'h1)];
              reg3354 <= (-$signed((reg3030[(1'h0):(1'h0)] && (reg3198[(4'hc):(3'h5)] < $signed(reg3239)))));
              reg3355 = (&$unsigned(reg3348[(2'h3):(1'h1)]));
            end
          else
            begin
              reg3349 <= (reg3071 ?
                  $signed(($unsigned((reg3296 ?
                      reg3102 : reg3071)) >= reg3237)) : (8'ha7));
              reg3350 = reg3343;
              reg3351 <= (reg3333[(2'h2):(1'h1)] <= ($signed(reg3022) & $signed((~&reg3250))));
              reg3354 <= $unsigned((~^(-reg3184[(1'h0):(1'h0)])));
              reg3355 = reg3183;
              reg3356 = (reg3323[(1'h1):(1'h0)] >>> (reg3063 ?
                  ((reg3128[(4'ha):(1'h1)] || reg3170[(5'h16):(1'h0)]) <<< reg3352[(3'h7):(2'h3)]) : (reg3340[(5'h12):(5'h10)] ?
                      $unsigned(((7'h40) < reg3323)) : $unsigned(reg2987[(2'h2):(2'h2)]))));
              reg3357 = reg3304;
            end
          if ((-((8'ha3) && reg3150[(5'h19):(5'h10)])))
            begin
              reg3358 = reg3194;
              reg3359 <= (|(reg3063[(4'hb):(2'h2)] - (|($unsigned(reg3018) ^ (8'ha2)))));
              reg3360 = (((reg3332 - reg3333[(3'h7):(1'h0)]) - reg3314[(5'h16):(3'h7)]) * reg3262[(5'h13):(3'h5)]);
              reg3361 <= $unsigned((((7'h4a) >= ((reg3360 ?
                      reg3340 : reg2991) | {reg3313, reg3257, reg3011})) ?
                  (reg3314[(4'ha):(4'h8)] << (&$unsigned(reg2962))) : $unsigned((&$signed(reg3189)))));
              reg3362 <= (7'h4c);
            end
          else
            begin
              reg3358 = reg3063;
              reg3359 <= (|(reg3344 ?
                  ($unsigned({reg3340, reg3206}) ?
                      reg3304[(4'hc):(3'h4)] : reg3015) : ($unsigned($signed((7'h4b))) < ({reg3020} | (forvar3318 || wire1689)))));
              reg3361 <= (({((reg3035 ?
                      reg3180 : reg3335) ^~ (reg3152 >>> reg3302)),
                  reg3273[(5'h12):(1'h0)],
                  (reg3280[(5'h12):(4'h9)] ^ (reg3004 <= (7'h51)))} * {(|(^reg3355)),
                  (((8'hbf) ? reg2954 : reg3075) ? (!reg3244) : (-reg3307)),
                  $signed((reg3106 ?
                      reg3309 : reg3205))}) < ((~&reg3077) && ((reg2993 <<< wire1692[(3'h7):(3'h6)]) ?
                  reg2949[(5'h17):(4'h9)] : (~^(reg3258 ?
                      reg3284 : reg3011)))));
              reg3362 <= (!(+reg3340));
              reg3363 = $signed($signed((!reg2969[(4'ha):(1'h0)])));
            end
        end
      else
        begin
          reg3331 = reg3161;
          for (forvar3332 = (1'h0); (forvar3332 < (2'h2)); forvar3332 = (forvar3332 + (1'h1)))
            begin
              reg3333 <= $signed(reg3321);
              reg3335 = wire1689;
              reg3337 <= reg3303;
              reg3339 = reg3295;
            end
        end
    end
  assign wire3364 = $signed(reg2969);
  always
    @(posedge clk) begin
      for (forvar3365 = (1'h0); (forvar3365 < (1'h0)); forvar3365 = (forvar3365 + (1'h1)))
        begin
          reg3366 = (reg3258 == {$unsigned(reg3003[(5'h14):(4'hf)]), reg3026});
          if (reg3208[(1'h0):(1'h0)])
            begin
              reg3367 <= $unsigned($unsigned((7'h4c)));
              reg3368 = $unsigned((($signed((reg3349 ? reg3094 : reg3152)) ?
                      reg3172[(3'h7):(3'h4)] : (~|(reg3099 ?
                          reg3113 : forvar3365))) ?
                  (|(^~reg3235[(2'h2):(1'h0)])) : $unsigned((reg3124 ^ {reg2980}))));
              reg3369 = (8'hb0);
              reg3370 <= reg3134[(4'h8):(3'h4)];
              reg3371 = (reg3238[(3'h5):(2'h2)] ?
                  (~|$unsigned($signed({(8'haf)}))) : (^~reg3345[(2'h3):(1'h1)]));
            end
          else
            begin
              reg3368 = $unsigned((^~(((reg3345 ~^ (7'h47)) ?
                  reg3312[(3'h4):(3'h4)] : reg3362) > ((^reg3122) << wire1690[(4'he):(1'h0)]))));
              reg3369 = ($unsigned(reg3298) * $signed({{(|reg3334),
                      (reg2967 ? (7'h58) : reg3132),
                      (reg3332 && reg3230)},
                  (&$unsigned(reg3240)),
                  ({wire1687} <= reg3234)}));
              reg3370 <= reg3226[(3'h4):(1'h1)];
              reg3372 <= ((^~reg3172[(4'hc):(1'h0)]) ?
                  reg3176[(5'h1a):(5'h16)] : reg3237[(5'h10):(3'h4)]);
              reg3373 <= ({((~|((8'hb4) ? reg3226 : reg3361)) ?
                          ((^reg3113) > (+(8'ha0))) : reg3322),
                      $signed($signed((reg3192 ? (8'hbc) : reg3367)))} ?
                  reg3368[(4'he):(3'h7)] : {($unsigned($signed(reg3009)) ?
                          ($unsigned(reg3012) << (&wire3036)) : $unsigned((reg3124 ?
                              reg3065 : reg3020)))});
              reg3374 <= (&reg3080[(1'h0):(1'h0)]);
            end
        end
      if ($signed($signed({reg3085[(5'h10):(4'hb)],
          wire1687[(4'ha):(2'h2)],
          ((^reg3165) ~^ (reg2955 ? reg2983 : reg3004))})))
        begin
          reg3375 = reg3038;
          for (forvar3376 = (1'h0); (forvar3376 < (3'h4)); forvar3376 = (forvar3376 + (1'h1)))
            begin
              reg3377 = (wire3268 ?
                  ($unsigned({(-reg3310),
                      reg3189[(4'hc):(2'h2)],
                      reg3237[(3'h6):(2'h2)]}) == $signed(((!reg3001) ?
                      (-wire3036) : (reg2980 ?
                          reg3020 : reg2950)))) : (^~$signed($unsigned($unsigned((7'h51))))));
              reg3378 = {reg3265[(5'h1b):(1'h0)],
                  {reg2949},
                  reg3144[(4'hb):(3'h6)]};
              reg3379 = (^~wire1689);
            end
          reg3380 <= {(reg3212[(3'h5):(2'h3)] != (({reg3288,
                      reg2954,
                      reg3046} >>> (wire1688 ? reg2969 : (8'ha6))) ?
                  (reg3161 || reg3265[(5'h17):(2'h3)]) : (^~reg3371)))};
        end
      else
        begin
          if ((-(7'h45)))
            begin
              reg3376 <= $signed(reg3124);
              reg3380 <= (8'hae);
              reg3381 = ((|$signed($unsigned((reg3310 >>> wire1691)))) ?
                  reg3312[(4'h8):(3'h4)] : reg3106[(4'h8):(3'h6)]);
              reg3382 = {$signed(reg3135[(4'hb):(3'h4)])};
              reg3383 <= $signed((($signed(reg3131[(1'h0):(1'h0)]) <= (-$signed(reg3253))) >> (~&$unsigned((reg2975 >> (7'h55))))));
              reg3384 <= (((reg3058 ?
                      $unsigned((reg3118 && forvar3376)) : $unsigned(reg3020[(1'h0):(1'h0)])) ^~ reg3298[(3'h7):(3'h4)]) ?
                  ((~^(reg3226[(1'h1):(1'h1)] ^ $signed(reg3374))) ?
                      $unsigned((reg3206 + (reg3267 ^ reg2987))) : $signed(($signed(wire3147) ?
                          reg3033 : (reg3046 ?
                              wire1691 : reg3293)))) : ($signed(wire3148) ^ {$signed(reg3243[(4'hf):(3'h6)])}));
              reg3385 = ($signed(reg3073[(3'h4):(1'h1)]) ?
                  $signed((~&$signed((7'h40)))) : ((^~reg3035) ?
                      ($unsigned(((7'h4b) ? reg3155 : (7'h4f))) ?
                          (&$signed(reg3102)) : (reg2952[(3'h5):(1'h0)] ?
                              (&reg3030) : (+reg3374))) : ((!{reg3063,
                              reg3253}) ?
                          (+(~(8'hb7))) : (reg3375[(4'hc):(2'h3)] * $signed(reg3011)))));
            end
          else
            begin
              reg3376 <= reg3273;
              reg3380 <= {$unsigned({{$unsigned(reg3098),
                          $unsigned(reg3288),
                          $unsigned(reg3343)},
                      reg3215}),
                  (!$unsigned({(^reg3102), $unsigned(reg3262)})),
                  {$signed($signed((wire1688 <= reg3308))),
                      (((reg3205 ? reg3332 : reg3284) ?
                              reg3226[(3'h5):(3'h4)] : (+reg3310)) ?
                          reg3101 : reg3065)}};
              reg3381 = reg3322[(3'h5):(3'h5)];
              reg3382 = reg3323[(3'h6):(3'h5)];
              reg3383 <= wire1689[(3'h5):(3'h5)];
              reg3384 <= (reg3372[(3'h5):(2'h2)] ?
                  ((reg3142 <= (~(!reg3004))) ^~ reg3293) : (~^reg3109));
              reg3385 = reg3102[(4'he):(3'h6)];
            end
          if ($unsigned($unsigned(wire1687)))
            begin
              reg3386 = ((|($signed(reg2965) == $unsigned(reg3374))) ?
                  (&$unsigned((7'h54))) : $signed(reg3222));
              reg3387 = (7'h50);
            end
          else
            begin
              reg3386 = reg3161;
              reg3387 = (reg3277[(1'h0):(1'h0)] <<< ($signed((((7'h47) ^ (8'hac)) && (reg3039 << (8'hb6)))) ?
                  (wire1692 >> (-(reg3190 & reg3132))) : {reg3110[(2'h2):(2'h2)],
                      ((&reg3337) <<< $unsigned((8'hb0))),
                      $unsigned($signed(reg3189))}));
              reg3388 = ($unsigned((($unsigned(reg3208) ?
                  $signed(reg2962) : (reg3023 + reg3047)) | ((reg3154 - reg3152) ?
                  reg3311 : (reg2951 ?
                      reg3094 : reg2981)))) ~^ (!$unsigned((~reg3033))));
            end
        end
      if (($signed($signed(reg3022[(5'h12):(4'hb)])) >>> ((^~reg2960[(1'h1):(1'h1)]) ?
          ($unsigned((reg3333 ? reg3198 : (8'hbe))) ?
              reg3152[(4'h9):(3'h5)] : {(reg3198 <<< reg3253)}) : $signed((reg3385 ?
              (~^reg3344) : (reg3235 ? reg3077 : reg2955))))))
        begin
          reg3389 = (({$unsigned(reg3337[(3'h6):(3'h4)])} ?
              (reg3192 ^~ (reg3065 ?
                  $unsigned(reg3154) : reg3316)) : {((~|reg3150) != $unsigned(reg3354)),
                  reg3047}) > (7'h4d));
        end
      else
        begin
          for (forvar3389 = (1'h0); (forvar3389 < (3'h5)); forvar3389 = (forvar3389 + (1'h1)))
            begin
              reg3390 = $unsigned(({{$unsigned(reg3188), $signed(reg3337)},
                      (~|(~(8'hb9))),
                      $unsigned(reg3205)} ?
                  (reg2967 ?
                      $unsigned((reg2997 ^~ reg3002)) : reg3180[(5'h14):(4'hc)]) : (^~(-(7'h54)))));
              reg3391 = $unsigned(reg3183);
              reg3392 <= (reg3190 ?
                  $signed((&$unsigned(reg3205))) : $unsigned(reg3361));
              reg3393 = reg3288;
              reg3394 = ({$signed(reg3163),
                      $signed(((reg3102 + reg3310) ?
                          $signed(reg3253) : $signed(reg3047))),
                      (8'ha4)} ?
                  (~&reg3266) : (&reg3116[(5'h11):(4'hd)]));
              reg3395 <= reg3338[(1'h1):(1'h1)];
            end
          reg3396 <= (^~(~$signed(((|wire3036) ?
              (reg3253 ? reg3152 : reg3378) : (7'h45)))));
          reg3397 = ($signed($signed(reg3234)) ?
              $unsigned($signed(reg3280[(5'h18):(5'h16)])) : reg3059);
          for (forvar3398 = (1'h0); (forvar3398 < (3'h5)); forvar3398 = (forvar3398 + (1'h1)))
            begin
              reg3399 = {(&((7'h53) & {(reg3284 == (8'had)),
                      reg2983,
                      $unsigned(reg3012)}))};
              reg3400 <= (reg3024 >> reg3382[(4'ha):(1'h1)]);
              reg3401 = reg3031;
              reg3402 <= ({reg3370,
                  (($signed((7'h56)) >>> (reg3071 ? reg3349 : reg3236)) ?
                      (^~(reg3012 ?
                          forvar3376 : (8'hba))) : reg3089[(3'h4):(1'h0)]),
                  $unsigned({(!forvar3398),
                      (^(7'h4d)),
                      (&reg3396)})} + (reg3200[(2'h2):(2'h2)] & {$signed($signed(reg3338)),
                  $unsigned({reg3239, reg2999})}));
            end
        end
      reg3403 <= reg2949[(1'h0):(1'h0)];
      reg3404 <= {(&(reg3300[(2'h2):(2'h2)] ? (~|reg3184) : reg3081)),
          reg3396[(3'h7):(3'h5)]};
    end
  assign wire3405 = (^$signed(reg3361));
  assign wire3406 = {reg3324[(5'h16):(4'he)]};
  assign wire3407 = (^~reg3118);
  assign wire3408 = reg3004[(5'h13):(4'ha)];
  assign wire3409 = reg3122;
  assign wire3410 = reg3343;
  always
    @(posedge clk) begin
      if (({reg3284[(2'h3):(2'h2)],
          reg3124[(3'h4):(2'h3)],
          wire2946[(2'h2):(1'h0)]} * $unsigned(reg3173)))
        begin
          if (({((reg3077 || reg3261) >= reg3359),
              reg2972[(1'h0):(1'h0)]} <<< {reg3093, $signed(reg3246)}))
            begin
              reg3411 <= (|reg2965[(3'h6):(3'h5)]);
              reg3412 <= $signed(reg3018);
              reg3413 = (^~$unsigned((($signed((8'hae)) ?
                      (~^wire3070) : (reg3309 ~^ reg2974)) ?
                  ($unsigned(reg3183) ~^ $unsigned(reg3161)) : $signed((7'h4f)))));
              reg3414 <= (((reg3206[(1'h1):(1'h1)] <<< $unsigned(wire1692[(3'h6):(3'h5)])) ^ reg3065) <= ($signed($unsigned((+reg3172))) ?
                  {wire3364[(4'h9):(3'h4)],
                      (~&(reg3118 >>> reg3155)),
                      ($signed(reg3033) * $signed(reg3106))} : reg3308[(1'h1):(1'h0)]));
              reg3415 <= $signed($unsigned((!reg3220)));
              reg3416 <= reg3250;
              reg3417 <= (~^reg3238[(3'h4):(2'h3)]);
            end
          else
            begin
              reg3413 = (reg3416 + ((&reg3113) ?
                  reg3192 : ($signed((reg3236 | reg3058)) == reg3304[(4'h9):(4'h8)])));
              reg3414 <= reg3372;
              reg3418 = {(reg3094 ?
                      (^~({reg3280,
                          reg3198} < $unsigned((8'hb3)))) : reg3110[(3'h6):(2'h3)]),
                  reg2975};
              reg3419 <= reg3316;
              reg3420 <= ((!$signed(reg3341[(3'h4):(3'h4)])) ?
                  ({((-wire1693) ?
                          ((7'h44) ?
                              reg3009 : reg3230) : $signed(reg3400))} != ({(8'hb5),
                      $unsigned(reg3015)} > (reg2962 >= {reg3265,
                      reg3220}))) : reg3188[(1'h1):(1'h0)]);
            end
          reg3421 = $signed($signed(((((8'haa) ?
              reg3235 : reg3337) < reg3093) >= reg2967)));
        end
      else
        begin
          if (($signed(({{(8'hbd), wire3410}, (7'h47), $unsigned((8'h9c))} ?
              reg3343[(2'h3):(2'h2)] : {reg3009[(1'h0):(1'h0)],
                  $unsigned(reg3340)})) && reg3194[(4'hd):(2'h3)]))
            begin
              reg3411 <= $unsigned($signed($signed(reg2955[(4'hd):(4'hb)])));
              reg3413 = ((($unsigned((reg3001 == (7'h46))) ?
                      $signed((reg3230 ?
                          reg3163 : (7'h4a))) : $unsigned((reg3246 ^ reg3079))) ?
                  reg3124[(1'h1):(1'h1)] : (reg3001 ?
                      wire3408[(2'h2):(1'h0)] : ($unsigned(reg3396) >>> (&reg3400)))) - (((-reg3332[(5'h17):(4'h8)]) ?
                      $signed((reg3412 ?
                          (8'ha5) : reg3165)) : (reg2951[(5'h11):(1'h1)] < (~^wire1687))) ?
                  (8'ha9) : $signed($signed((reg3194 ? (8'ha9) : (8'hbe))))));
            end
          else
            begin
              reg3413 = reg3005;
              reg3418 = (({$signed((^~reg3011)),
                      ($signed((8'hbc)) >= reg3089[(2'h2):(1'h0)])} || $signed(reg3266)) ?
                  reg3027[(1'h1):(1'h0)] : reg3392);
              reg3421 = (((8'haf) ~^ $signed(reg2949[(4'hd):(4'hb)])) >>> reg3067[(3'h5):(3'h4)]);
              reg3422 = ({($unsigned($signed(reg2974)) ? reg3118 : reg3170),
                      (reg3004[(3'h4):(2'h2)] | $signed($signed((7'h57))))} ?
                  $signed($unsigned($signed($signed(reg3102)))) : reg3383[(3'h5):(1'h0)]);
              reg3423 = ((~|(!($signed(wire1689) >= {reg2980}))) == reg3094[(1'h0):(1'h0)]);
            end
          for (forvar3424 = (1'h0); (forvar3424 < (2'h3)); forvar3424 = (forvar3424 + (1'h1)))
            begin
              reg3425 = ((^~(~$signed($unsigned(reg3118)))) >>> $unsigned({$unsigned(reg3414)}));
            end
        end
      for (forvar3426 = (1'h0); (forvar3426 < (3'h6)); forvar3426 = (forvar3426 + (1'h1)))
        begin
          if (reg3190)
            begin
              reg3427 = {(|(|reg3422[(1'h0):(1'h0)]))};
              reg3428 <= $unsigned(({(&(8'had)),
                      ({reg2950} ? $unsigned(reg2969) : {wire3406, reg3001})} ?
                  (reg3043[(4'hb):(3'h5)] ?
                      reg3300[(3'h4):(3'h4)] : {$unsigned(reg3323),
                          {reg2997, reg3367, wire3407},
                          (reg3396 != reg3297)}) : reg3002));
              reg3429 = reg3218[(5'h1a):(5'h16)];
              reg3430 <= (({(&(8'hbd)),
                          reg2972,
                          (~^((8'ha8) ? reg3374 : reg2981))} ?
                      (reg3022 ?
                          reg3423[(2'h2):(1'h0)] : ((reg3248 || reg3414) == reg3337[(2'h3):(1'h1)])) : $signed(reg3402[(4'h8):(3'h5)])) ?
                  reg3128 : ((reg3058 >> ($signed((8'hb0)) ?
                      $unsigned(reg3341) : $unsigned(reg3248))) ^~ $signed(($unsigned(reg3346) ?
                      $unsigned(reg3422) : reg3059[(2'h3):(2'h3)]))));
              reg3431 <= ($signed(reg3131) ?
                  ({$signed(wire3410),
                      reg3246[(3'h4):(1'h1)]} != (($unsigned(reg2991) | (reg3173 ?
                          reg3080 : reg3373)) ?
                      ($unsigned(reg3194) | $unsigned(reg3194)) : $signed($unsigned(reg3009)))) : (|(!($unsigned(reg3296) | $unsigned(reg3022)))));
              reg3432 = reg3079[(4'hb):(3'h6)];
              reg3433 = (((|($signed(reg2952) && reg3234)) ?
                      {{(reg3280 && reg3332)}, reg3058} : reg3304) ?
                  $signed(reg3155[(5'h19):(4'hf)]) : $signed($unsigned((+reg3232))));
            end
          else
            begin
              reg3428 <= {$unsigned(reg3380),
                  $unsigned((((~|reg3093) ?
                          (reg3046 <= reg3373) : (&wire1692)) ?
                      (reg3235[(4'h8):(3'h5)] << reg2969[(1'h1):(1'h0)]) : $unsigned($unsigned(reg3026)))),
                  $unsigned((($unsigned(reg3258) >= $signed(reg3205)) ?
                      ((reg3295 ?
                          reg3173 : reg3230) >= (reg3166 > (7'h52))) : (~^reg3312[(4'ha):(1'h1)])))};
              reg3429 = $signed((-reg3404[(5'h1a):(4'hf)]));
              reg3430 <= $signed(wire1692[(1'h0):(1'h0)]);
              reg3432 = $unsigned($signed(reg3184[(3'h5):(3'h5)]));
              reg3434 <= reg3030[(5'h14):(4'h8)];
              reg3435 <= reg3311[(1'h0):(1'h0)];
            end
          if (reg3020)
            begin
              reg3436 <= ((-(((&reg3361) ?
                      $signed(reg3079) : (reg3428 ? reg3004 : reg3367)) ?
                  $signed((!reg3134)) : reg3380)) <= $unsigned($signed(reg3124[(1'h0):(1'h0)])));
              reg3437 <= ($unsigned(((^~reg3168[(5'h15):(4'h9)]) << {reg3354,
                      reg3106})) ?
                  $signed(({reg3228[(5'h1c):(4'h8)]} ?
                      reg3343[(1'h1):(1'h1)] : ((reg3273 ? reg3288 : (7'h41)) ?
                          $unsigned(reg3020) : (reg3230 ?
                              reg3266 : (8'h9d))))) : (&$signed(($unsigned(reg3071) ?
                      {(7'h46), reg3089} : reg3337))));
              reg3438 <= ((+((reg3238[(3'h6):(2'h3)] ?
                      (7'h46) : ((8'hb7) ?
                          reg3280 : reg3134)) >= (reg3428[(4'ha):(4'h8)] ?
                      ((8'ha8) ?
                          reg3228 : reg3432) : reg3240[(3'h5):(1'h1)]))) ?
                  ((reg3116[(5'h11):(4'h8)] ?
                          ((&reg3323) ^ $unsigned(reg3253)) : wire1694[(5'h13):(2'h3)]) ?
                      (~^$unsigned($unsigned(reg2991))) : reg3012) : reg2991);
              reg3439 <= $signed(reg3022[(2'h2):(1'h0)]);
              reg3440 = reg2997;
              reg3441 = ($unsigned($signed(reg3332)) >>> $unsigned($signed($signed($signed(wire3405)))));
              reg3442 = ($unsigned(reg3215) ^ (reg3380[(3'h5):(2'h2)] ?
                  $unsigned($signed($signed(reg3312))) : (reg3194[(5'h16):(3'h4)] ?
                      reg3429 : ($unsigned(reg3346) ?
                          (&(8'ha1)) : reg3380[(4'hc):(4'hc)]))));
            end
          else
            begin
              reg3436 <= ($unsigned(reg3041[(1'h0):(1'h0)]) >= reg3009);
              reg3440 = (reg3432 ?
                  (!($unsigned($signed(reg3427)) <= (reg3237[(4'he):(4'hb)] ?
                      $signed(reg3429) : reg3370))) : ($unsigned((^((7'h46) < reg3309))) ^~ reg3220[(5'h13):(4'h8)]));
              reg3441 = (((^~$signed($signed(reg3428))) != reg3176) ?
                  ({((~|reg2999) && (-reg3101)),
                          {$signed(reg3277), $signed(reg3367), wire1694},
                          $signed((~reg3312))} ?
                      reg3065 : $signed(wire3147[(5'h11):(3'h7)])) : (7'h44));
              reg3443 <= ((^~(($signed(reg3396) > $signed(reg3032)) ?
                  $signed((^~(7'h40))) : reg3131)) <<< $signed($signed(($signed(reg3415) - $unsigned(reg3311)))));
            end
          reg3444 = $unsigned(reg3144[(4'h9):(3'h6)]);
          for (forvar3445 = (1'h0); (forvar3445 < (3'h6)); forvar3445 = (forvar3445 + (1'h1)))
            begin
              reg3446 = $signed({{$unsigned($signed(reg3022))},
                  ($unsigned($unsigned(reg3228)) + $signed((reg3168 | reg3296))),
                  wire1691});
              reg3447 <= reg3166[(2'h3):(1'h0)];
              reg3448 <= (^~reg3142[(4'h9):(2'h2)]);
              reg3449 <= ((8'ha1) | $signed({$signed({reg3348}),
                  (~{wire3408}),
                  $unsigned(reg3099[(5'h19):(5'h18)])}));
              reg3450 = $unsigned(($unsigned(reg2981[(5'h14):(4'ha)]) ?
                  reg3033[(2'h3):(1'h1)] : reg3334[(2'h2):(1'h1)]));
            end
        end
      reg3451 = $signed(reg3059[(3'h6):(2'h3)]);
      for (forvar3452 = (1'h0); (forvar3452 < (2'h2)); forvar3452 = (forvar3452 + (1'h1)))
        begin
          reg3453 = $unsigned((($signed(reg3266[(2'h2):(1'h0)]) ^~ (~^(forvar3452 <= reg3226))) ?
              (~|{reg3267}) : ({(~^forvar3426),
                  reg3400,
                  {reg3340}} != {{reg3362, wire3410, reg3446},
                  (reg2997 ? (8'ha2) : wire3147)})));
          reg3454 <= (($unsigned($unsigned({reg3316, reg3244})) ?
              {((reg3404 + reg3032) || reg2999)} : {reg3169[(5'h15):(1'h0)]}) <= (8'h9f));
          reg3455 = {$unsigned($unsigned((reg3024[(3'h4):(3'h4)] <<< reg2987[(3'h7):(3'h7)]))),
              {(^~{reg3018, reg3035, (7'h4c)}),
                  (reg3079 << (reg3257 ? (^reg3033) : (reg3169 < reg3288))),
                  ((^~(reg3403 & (8'hbd))) ?
                      (!reg3200[(4'he):(3'h7)]) : reg3101)}};
          for (forvar3456 = (1'h0); (forvar3456 < (1'h0)); forvar3456 = (forvar3456 + (1'h1)))
            begin
              reg3457 <= (^~(8'hb2));
            end
          reg3458 = ($signed((reg3418[(2'h3):(2'h2)] <<< reg3059)) ?
              {(($unsigned(wire3036) ?
                          reg2965[(2'h3):(2'h2)] : reg3180[(4'h8):(2'h3)]) ?
                      $unsigned((reg3173 <= reg3094)) : ($signed((8'h9c)) ?
                          $unsigned(reg3280) : $unsigned(reg3412)))} : $signed(((^~$unsigned(reg3134)) ^~ $signed(reg3450[(3'h4):(1'h1)]))));
        end
      for (forvar3459 = (1'h0); (forvar3459 < (3'h5)); forvar3459 = (forvar3459 + (1'h1)))
        begin
          if ($signed($unsigned($unsigned(((-reg3288) ?
              $signed(reg3176) : $signed((8'ha3)))))))
            begin
              reg3460 <= (wire3406 && reg3438[(3'h5):(3'h5)]);
              reg3461 <= $signed(((+$unsigned((-(7'h52)))) ?
                  (($signed(reg3296) ?
                          (^wire3096) : (reg3392 ? reg3374 : reg3206)) ?
                      reg3416[(1'h0):(1'h0)] : ($unsigned((8'haa)) ?
                          (reg3404 << reg3403) : (~^reg3015))) : (~reg3250[(5'h10):(2'h2)])));
              reg3462 <= ($signed($signed($unsigned((reg3416 | reg3372)))) ?
                  reg3396 : $signed((~^(~|reg3059[(3'h4):(2'h2)]))));
              reg3463 <= $unsigned(reg3206);
              reg3464 <= ((7'h58) ?
                  reg3135 : (($unsigned($signed(reg3102)) ?
                      ($signed(reg3250) ?
                          $unsigned(reg3443) : reg3176[(2'h3):(2'h3)]) : reg3277[(2'h2):(2'h2)]) & reg3198));
              reg3465 <= reg3026[(2'h2):(2'h2)];
              reg3466 <= ($unsigned({$unsigned(reg3012)}) << reg3421[(3'h4):(1'h0)]);
            end
          else
            begin
              reg3460 <= {reg2955};
              reg3461 <= reg3396;
              reg3467 = ({(8'hbb)} <<< reg3463);
              reg3468 = wire3364;
              reg3469 <= $unsigned(((reg2974 ?
                      ({reg3248, wire3147, reg2981} ?
                          $signed((7'h4d)) : forvar3445) : $signed((reg3168 == wire2946))) ?
                  $unsigned((reg3085[(4'hb):(2'h2)] ?
                      (reg3228 || reg3430) : reg2975[(1'h1):(1'h1)])) : $signed(reg3463[(3'h7):(3'h4)])));
              reg3470 = $signed(reg3128[(5'h10):(5'h10)]);
              reg3471 <= $signed(reg3033[(2'h3):(1'h0)]);
            end
          reg3472 = (^~reg3098[(3'h7):(2'h2)]);
          for (forvar3473 = (1'h0); (forvar3473 < (3'h6)); forvar3473 = (forvar3473 + (1'h1)))
            begin
              reg3474 = (~&{$signed((~$unsigned((7'h49)))),
                  {(8'hbd),
                      ($signed(reg3161) ? reg3429[(3'h6):(1'h0)] : reg3323),
                      (wire3364[(3'h4):(2'h2)] >= reg2967)},
                  $unsigned(((reg3165 ? reg2981 : reg3184) <<< {reg3419,
                      reg3412}))});
              reg3475 <= reg3421[(4'h9):(2'h2)];
              reg3476 <= (~&$signed(({{(8'ha9)}} <= (|(~&reg3165)))));
            end
        end
      reg3477 = reg3220;
    end
  always
    @(posedge clk) begin
      reg3478 <= reg3323;
    end
  module2644 #() modinst3480 (wire3479, clk, reg3436, reg3402, reg3152, reg3047);
  module2877 #() modinst3482 (.wire2878(reg3107), .wire2879(reg3122), .y(wire3481), .wire2882(reg3471), .clk(clk), .wire2881(reg2997), .wire2880(wire3409));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module92
#(parameter param1443 = ((^~((|((8'ha5) ? (8'ha7) : (8'h9e))) ? (((7'h4e) <= (8'hb1)) * (~&(8'ha5))) : ({(7'h51)} != ((7'h4a) ? (8'h9d) : (7'h52))))) * (!{((&(8'hb8)) ? ((7'h45) < (7'h40)) : ((7'h51) * (8'hb4))), ({(8'haf), (8'ha5)} == (+(7'h53)))})))
(y, clk, wire97, wire96, wire95, wire94, wire93);
  output wire [(32'h2507):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire97;
  input wire signed [(5'h15):(1'h0)] wire96;
  input wire signed [(4'hc):(1'h0)] wire95;
  input wire [(5'h13):(1'h0)] wire94;
  input wire [(5'h1e):(1'h0)] wire93;
  wire signed [(5'h1c):(1'h0)] wire1425;
  wire signed [(3'h4):(1'h0)] wire1367;
  wire signed [(5'h13):(1'h0)] wire1365;
  wire [(5'h13):(1'h0)] wire523;
  wire [(5'h1f):(1'h0)] wire435;
  wire signed [(5'h1d):(1'h0)] wire383;
  wire [(4'hc):(1'h0)] wire382;
  wire signed [(5'h18):(1'h0)] wire273;
  wire [(3'h7):(1'h0)] wire272;
  reg [(4'hc):(1'h0)] reg1441 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1439 = (1'h0);
  reg [(5'h13):(1'h0)] reg1437 = (1'h0);
  reg [(4'h9):(1'h0)] reg1435 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1434 = (1'h0);
  reg [(4'h9):(1'h0)] reg1433 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1431 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1430 = (1'h0);
  reg [(4'h8):(1'h0)] reg1428 = (1'h0);
  reg [(4'h8):(1'h0)] reg1424 = (1'h0);
  reg [(5'h17):(1'h0)] reg1419 = (1'h0);
  reg [(5'h12):(1'h0)] reg1418 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1414 = (1'h0);
  reg [(4'h8):(1'h0)] reg1412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1411 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1409 = (1'h0);
  reg [(3'h4):(1'h0)] reg1407 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1403 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1401 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1398 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1397 = (1'h0);
  reg [(3'h5):(1'h0)] reg1395 = (1'h0);
  reg [(4'ha):(1'h0)] reg1393 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1391 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1388 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1386 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1385 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1382 = (1'h0);
  reg [(3'h6):(1'h0)] reg1381 = (1'h0);
  reg [(5'h19):(1'h0)] reg1379 = (1'h0);
  reg [(5'h16):(1'h0)] reg1378 = (1'h0);
  reg [(5'h18):(1'h0)] reg1377 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1375 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1374 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1371 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1370 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg558 = (1'h0);
  reg [(5'h15):(1'h0)] reg557 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg555 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg553 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg551 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg550 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg544 = (1'h0);
  reg [(3'h4):(1'h0)] reg543 = (1'h0);
  reg signed [(4'he):(1'h0)] reg542 = (1'h0);
  reg [(5'h17):(1'h0)] reg540 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg539 = (1'h0);
  reg [(5'h1e):(1'h0)] reg535 = (1'h0);
  reg [(4'hb):(1'h0)] reg530 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg527 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg525 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg524 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg522 = (1'h0);
  reg [(3'h6):(1'h0)] reg521 = (1'h0);
  reg [(5'h15):(1'h0)] reg520 = (1'h0);
  reg [(4'he):(1'h0)] reg519 = (1'h0);
  reg [(5'h16):(1'h0)] reg518 = (1'h0);
  reg [(3'h7):(1'h0)] reg517 = (1'h0);
  reg [(5'h15):(1'h0)] reg514 = (1'h0);
  reg [(4'hd):(1'h0)] reg512 = (1'h0);
  reg [(5'h1a):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg508 = (1'h0);
  reg [(5'h16):(1'h0)] reg507 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg506 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg505 = (1'h0);
  reg [(5'h12):(1'h0)] reg504 = (1'h0);
  reg [(5'h15):(1'h0)] reg503 = (1'h0);
  reg [(5'h18):(1'h0)] reg501 = (1'h0);
  reg [(2'h2):(1'h0)] reg500 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg498 = (1'h0);
  reg [(5'h1d):(1'h0)] reg496 = (1'h0);
  reg [(4'hc):(1'h0)] reg491 = (1'h0);
  reg [(3'h7):(1'h0)] reg490 = (1'h0);
  reg [(2'h2):(1'h0)] reg482 = (1'h0);
  reg [(5'h16):(1'h0)] reg481 = (1'h0);
  reg [(3'h6):(1'h0)] reg479 = (1'h0);
  reg [(4'h8):(1'h0)] reg470 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg468 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg467 = (1'h0);
  reg [(5'h13):(1'h0)] reg466 = (1'h0);
  reg [(4'h9):(1'h0)] reg465 = (1'h0);
  reg [(4'hb):(1'h0)] reg463 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg461 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg460 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg457 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg456 = (1'h0);
  reg [(5'h10):(1'h0)] reg454 = (1'h0);
  reg [(2'h2):(1'h0)] reg453 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg452 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg450 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg445 = (1'h0);
  reg [(5'h10):(1'h0)] reg443 = (1'h0);
  reg [(5'h1f):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg440 = (1'h0);
  reg [(5'h16):(1'h0)] reg439 = (1'h0);
  reg [(5'h1a):(1'h0)] reg437 = (1'h0);
  reg [(5'h16):(1'h0)] reg434 = (1'h0);
  reg [(5'h19):(1'h0)] reg432 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg428 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg426 = (1'h0);
  reg [(5'h14):(1'h0)] reg420 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg419 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg418 = (1'h0);
  reg [(5'h18):(1'h0)] reg417 = (1'h0);
  reg [(5'h1b):(1'h0)] reg413 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg411 = (1'h0);
  reg [(5'h1d):(1'h0)] reg410 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg407 = (1'h0);
  reg [(4'h8):(1'h0)] reg403 = (1'h0);
  reg [(4'ha):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg391 = (1'h0);
  reg [(5'h12):(1'h0)] reg390 = (1'h0);
  reg [(3'h5):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg384 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg381 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg373 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg371 = (1'h0);
  reg [(3'h6):(1'h0)] reg370 = (1'h0);
  reg [(5'h17):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg366 = (1'h0);
  reg [(4'hc):(1'h0)] reg364 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg362 = (1'h0);
  reg [(4'hd):(1'h0)] reg360 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg358 = (1'h0);
  reg [(5'h1c):(1'h0)] reg357 = (1'h0);
  reg [(5'h19):(1'h0)] reg354 = (1'h0);
  reg [(4'hc):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg352 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg349 = (1'h0);
  reg [(4'h8):(1'h0)] reg347 = (1'h0);
  reg [(5'h13):(1'h0)] reg344 = (1'h0);
  reg [(5'h1f):(1'h0)] reg343 = (1'h0);
  reg [(4'hc):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg341 = (1'h0);
  reg [(2'h2):(1'h0)] reg340 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg337 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg336 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg335 = (1'h0);
  reg [(3'h6):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg329 = (1'h0);
  reg [(3'h6):(1'h0)] reg325 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg310 = (1'h0);
  reg [(4'hf):(1'h0)] reg300 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg320 = (1'h0);
  reg [(5'h1d):(1'h0)] reg317 = (1'h0);
  reg [(5'h18):(1'h0)] reg316 = (1'h0);
  reg [(5'h13):(1'h0)] reg314 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg313 = (1'h0);
  reg [(5'h1f):(1'h0)] reg309 = (1'h0);
  reg [(5'h1e):(1'h0)] reg308 = (1'h0);
  reg [(4'he):(1'h0)] reg307 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg305 = (1'h0);
  reg [(5'h1e):(1'h0)] reg296 = (1'h0);
  reg [(5'h13):(1'h0)] reg295 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg293 = (1'h0);
  reg [(2'h2):(1'h0)] reg292 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg290 = (1'h0);
  reg [(5'h1d):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg286 = (1'h0);
  reg [(5'h1b):(1'h0)] reg283 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg277 = (1'h0);
  reg [(4'he):(1'h0)] reg270 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg268 = (1'h0);
  reg signed [(4'he):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg265 = (1'h0);
  reg [(4'hf):(1'h0)] reg264 = (1'h0);
  reg [(4'ha):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg262 = (1'h0);
  reg [(4'hd):(1'h0)] reg260 = (1'h0);
  reg [(4'ha):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg250 = (1'h0);
  reg [(5'h1d):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg246 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg243 = (1'h0);
  reg [(4'ha):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg239 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg236 = (1'h0);
  reg [(3'h7):(1'h0)] reg230 = (1'h0);
  reg [(3'h7):(1'h0)] reg229 = (1'h0);
  reg [(5'h19):(1'h0)] reg227 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg224 = (1'h0);
  reg [(5'h12):(1'h0)] reg223 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg221 = (1'h0);
  reg [(4'hb):(1'h0)] reg220 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg219 = (1'h0);
  reg [(5'h19):(1'h0)] reg216 = (1'h0);
  reg [(4'hf):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg214 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg210 = (1'h0);
  reg [(5'h18):(1'h0)] reg207 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg201 = (1'h0);
  reg [(3'h7):(1'h0)] reg196 = (1'h0);
  reg [(4'he):(1'h0)] reg172 = (1'h0);
  reg [(5'h10):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg189 = (1'h0);
  reg [(4'he):(1'h0)] reg185 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg181 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg179 = (1'h0);
  reg [(5'h19):(1'h0)] reg178 = (1'h0);
  reg signed [(4'he):(1'h0)] reg174 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg173 = (1'h0);
  reg [(4'ha):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg169 = (1'h0);
  reg [(2'h2):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg166 = (1'h0);
  reg [(5'h14):(1'h0)] reg165 = (1'h0);
  reg [(4'ha):(1'h0)] reg164 = (1'h0);
  reg [(5'h19):(1'h0)] reg161 = (1'h0);
  reg [(5'h15):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg156 = (1'h0);
  reg [(4'hb):(1'h0)] reg153 = (1'h0);
  reg [(4'he):(1'h0)] reg152 = (1'h0);
  reg [(4'he):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg150 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg147 = (1'h0);
  reg [(5'h10):(1'h0)] reg145 = (1'h0);
  reg [(5'h14):(1'h0)] reg142 = (1'h0);
  reg [(5'h14):(1'h0)] reg141 = (1'h0);
  reg signed [(4'he):(1'h0)] reg138 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg137 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg135 = (1'h0);
  reg [(2'h2):(1'h0)] reg133 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg132 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg131 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg128 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg127 = (1'h0);
  reg [(5'h16):(1'h0)] reg123 = (1'h0);
  reg [(5'h1f):(1'h0)] reg122 = (1'h0);
  reg [(4'h9):(1'h0)] reg121 = (1'h0);
  reg [(5'h1f):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg117 = (1'h0);
  reg [(5'h11):(1'h0)] reg116 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg113 = (1'h0);
  reg [(4'hb):(1'h0)] reg112 = (1'h0);
  reg [(4'hc):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg109 = (1'h0);
  reg [(5'h1e):(1'h0)] reg105 = (1'h0);
  reg [(5'h10):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg98 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1442 = (1'h0);
  reg [(3'h4):(1'h0)] reg1440 = (1'h0);
  reg [(5'h12):(1'h0)] reg1438 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1436 = (1'h0);
  reg [(4'ha):(1'h0)] reg1432 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1429 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1427 = (1'h0);
  reg [(3'h7):(1'h0)] reg1426 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1423 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1422 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1421 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1420 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1417 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1416 = (1'h0);
  reg [(3'h7):(1'h0)] reg1415 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1413 = (1'h0);
  reg [(5'h19):(1'h0)] reg1410 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1406 = (1'h0);
  reg [(5'h10):(1'h0)] reg1405 = (1'h0);
  reg [(5'h19):(1'h0)] reg1404 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1402 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1400 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1399 = (1'h0);
  reg [(5'h11):(1'h0)] reg1396 = (1'h0);
  reg [(5'h12):(1'h0)] reg1394 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1392 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1390 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1389 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1387 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1384 = (1'h0);
  reg [(2'h3):(1'h0)] reg1383 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1380 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1376 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1373 = (1'h0);
  reg [(5'h17):(1'h0)] reg1372 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1369 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1368 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg560 = (1'h0);
  reg [(5'h12):(1'h0)] reg559 = (1'h0);
  reg [(5'h1a):(1'h0)] reg556 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg554 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar549 = (1'h0);
  reg [(3'h6):(1'h0)] reg548 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar547 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg545 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar541 = (1'h0);
  reg [(4'hf):(1'h0)] forvar538 = (1'h0);
  reg [(2'h2):(1'h0)] reg537 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg536 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg534 = (1'h0);
  reg [(4'hb):(1'h0)] reg533 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg531 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar528 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg516 = (1'h0);
  reg [(5'h17):(1'h0)] forvar515 = (1'h0);
  reg [(5'h16):(1'h0)] forvar513 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar511 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar504 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg515 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar514 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar512 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg511 = (1'h0);
  reg [(5'h19):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg502 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg497 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar495 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg494 = (1'h0);
  reg [(2'h2):(1'h0)] reg493 = (1'h0);
  reg [(2'h2):(1'h0)] reg492 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg489 = (1'h0);
  reg [(3'h7):(1'h0)] reg488 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg486 = (1'h0);
  reg [(5'h18):(1'h0)] reg485 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg484 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg483 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg478 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar476 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg475 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg474 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar473 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar471 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg469 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg464 = (1'h0);
  reg [(5'h1b):(1'h0)] reg462 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar436 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg451 = (1'h0);
  reg [(4'hf):(1'h0)] reg449 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg447 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg446 = (1'h0);
  reg [(4'h8):(1'h0)] reg444 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg442 = (1'h0);
  reg [(5'h14):(1'h0)] reg438 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg436 = (1'h0);
  reg [(5'h10):(1'h0)] reg433 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar431 = (1'h0);
  reg [(5'h1f):(1'h0)] reg430 = (1'h0);
  reg [(5'h1a):(1'h0)] reg429 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg427 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg425 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar424 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg422 = (1'h0);
  reg [(3'h6):(1'h0)] reg421 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg416 = (1'h0);
  reg [(5'h12):(1'h0)] reg415 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg414 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg412 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg406 = (1'h0);
  reg [(4'h8):(1'h0)] forvar405 = (1'h0);
  reg [(5'h1d):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg401 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar397 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg396 = (1'h0);
  reg [(5'h19):(1'h0)] forvar394 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg392 = (1'h0);
  reg [(4'h9):(1'h0)] reg389 = (1'h0);
  reg [(4'he):(1'h0)] forvar387 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg386 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg385 = (1'h0);
  reg [(5'h16):(1'h0)] reg380 = (1'h0);
  reg [(5'h19):(1'h0)] reg378 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar377 = (1'h0);
  reg [(5'h16):(1'h0)] reg376 = (1'h0);
  reg [(5'h1a):(1'h0)] reg372 = (1'h0);
  reg [(5'h16):(1'h0)] reg369 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg367 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar365 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar363 = (1'h0);
  reg [(4'h8):(1'h0)] forvar361 = (1'h0);
  reg signed [(4'he):(1'h0)] reg356 = (1'h0);
  reg [(4'hb):(1'h0)] reg355 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg350 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg348 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar345 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar339 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg338 = (1'h0);
  reg [(4'h9):(1'h0)] reg333 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg332 = (1'h0);
  reg [(5'h1c):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar330 = (1'h0);
  reg [(3'h7):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg326 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar314 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar307 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg324 = (1'h0);
  reg [(4'h8):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg321 = (1'h0);
  reg [(4'hd):(1'h0)] reg319 = (1'h0);
  reg [(4'ha):(1'h0)] reg318 = (1'h0);
  reg [(3'h7):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg312 = (1'h0);
  reg [(5'h1b):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar310 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg306 = (1'h0);
  reg [(5'h1e):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg303 = (1'h0);
  reg [(5'h14):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg301 = (1'h0);
  reg [(4'hf):(1'h0)] forvar300 = (1'h0);
  reg [(5'h17):(1'h0)] forvar296 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar293 = (1'h0);
  reg [(5'h10):(1'h0)] reg299 = (1'h0);
  reg [(5'h1e):(1'h0)] reg298 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg297 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg291 = (1'h0);
  reg [(5'h11):(1'h0)] reg288 = (1'h0);
  reg [(3'h5):(1'h0)] reg287 = (1'h0);
  reg [(2'h3):(1'h0)] reg285 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg284 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg282 = (1'h0);
  reg [(5'h18):(1'h0)] reg281 = (1'h0);
  reg [(5'h1f):(1'h0)] forvar280 = (1'h0);
  reg [(5'h1a):(1'h0)] reg279 = (1'h0);
  reg [(5'h11):(1'h0)] reg278 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg276 = (1'h0);
  reg [(2'h3):(1'h0)] forvar275 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar274 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar269 = (1'h0);
  reg signed [(4'he):(1'h0)] reg267 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg261 = (1'h0);
  reg [(5'h19):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg258 = (1'h0);
  reg [(3'h5):(1'h0)] reg256 = (1'h0);
  reg [(3'h6):(1'h0)] forvar255 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg254 = (1'h0);
  reg [(5'h14):(1'h0)] reg253 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar252 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg251 = (1'h0);
  reg [(4'he):(1'h0)] reg249 = (1'h0);
  reg [(4'h8):(1'h0)] forvar247 = (1'h0);
  reg [(5'h13):(1'h0)] reg245 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg242 = (1'h0);
  reg [(5'h1a):(1'h0)] reg240 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg235 = (1'h0);
  reg [(3'h4):(1'h0)] forvar234 = (1'h0);
  reg [(5'h1f):(1'h0)] reg233 = (1'h0);
  reg [(2'h2):(1'h0)] forvar232 = (1'h0);
  reg [(5'h1f):(1'h0)] reg231 = (1'h0);
  reg [(3'h7):(1'h0)] reg228 = (1'h0);
  reg [(5'h11):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg225 = (1'h0);
  reg [(5'h18):(1'h0)] reg209 = (1'h0);
  reg [(5'h19):(1'h0)] forvar204 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar218 = (1'h0);
  reg [(5'h12):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar212 = (1'h0);
  reg [(2'h3):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar209 = (1'h0);
  reg [(5'h10):(1'h0)] reg208 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg205 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg204 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg200 = (1'h0);
  reg [(5'h1b):(1'h0)] reg199 = (1'h0);
  reg [(5'h1d):(1'h0)] reg198 = (1'h0);
  reg [(5'h1f):(1'h0)] reg197 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar195 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg194 = (1'h0);
  reg [(4'hc):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar188 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg187 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg186 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar180 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg177 = (1'h0);
  reg [(5'h14):(1'h0)] reg176 = (1'h0);
  reg [(5'h1a):(1'h0)] reg175 = (1'h0);
  reg [(5'h10):(1'h0)] forvar172 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg170 = (1'h0);
  reg [(4'hc):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg163 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar162 = (1'h0);
  reg [(4'h8):(1'h0)] reg158 = (1'h0);
  reg [(4'ha):(1'h0)] reg157 = (1'h0);
  reg [(3'h4):(1'h0)] reg155 = (1'h0);
  reg [(5'h1b):(1'h0)] reg154 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg149 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar135 = (1'h0);
  reg [(4'h9):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg144 = (1'h0);
  reg [(5'h18):(1'h0)] reg143 = (1'h0);
  reg [(5'h11):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg139 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg136 = (1'h0);
  reg [(4'h9):(1'h0)] reg134 = (1'h0);
  reg [(4'ha):(1'h0)] forvar130 = (1'h0);
  reg [(5'h1f):(1'h0)] reg129 = (1'h0);
  reg [(5'h14):(1'h0)] reg126 = (1'h0);
  reg [(5'h14):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar118 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg114 = (1'h0);
  reg signed [(4'he):(1'h0)] reg110 = (1'h0);
  reg [(5'h15):(1'h0)] reg108 = (1'h0);
  reg [(3'h7):(1'h0)] reg107 = (1'h0);
  reg [(4'hd):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg103 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg102 = (1'h0);
  reg [(4'hd):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg100 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar99 = (1'h0);
  assign y = {wire1425,
                 wire1367,
                 wire1365,
                 wire523,
                 wire435,
                 wire383,
                 wire382,
                 wire273,
                 wire272,
                 reg1441,
                 reg1439,
                 reg1437,
                 reg1435,
                 reg1434,
                 reg1433,
                 reg1431,
                 reg1430,
                 reg1428,
                 reg1424,
                 reg1419,
                 reg1418,
                 reg1414,
                 reg1412,
                 reg1411,
                 reg1409,
                 reg1407,
                 reg1403,
                 reg1401,
                 reg1398,
                 reg1397,
                 reg1395,
                 reg1393,
                 reg1391,
                 reg1388,
                 reg1386,
                 reg1385,
                 reg1382,
                 reg1381,
                 reg1379,
                 reg1378,
                 reg1377,
                 reg1375,
                 reg1374,
                 reg1371,
                 reg1370,
                 reg558,
                 reg557,
                 reg555,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg544,
                 reg543,
                 reg542,
                 reg540,
                 reg539,
                 reg535,
                 reg530,
                 reg529,
                 reg527,
                 reg525,
                 reg524,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 reg514,
                 reg512,
                 reg510,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg501,
                 reg500,
                 reg498,
                 reg496,
                 reg491,
                 reg490,
                 reg482,
                 reg481,
                 reg479,
                 reg470,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg463,
                 reg461,
                 reg460,
                 reg457,
                 reg456,
                 reg454,
                 reg453,
                 reg452,
                 reg450,
                 reg448,
                 reg445,
                 reg443,
                 reg441,
                 reg440,
                 reg439,
                 reg437,
                 reg434,
                 reg432,
                 reg428,
                 reg426,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg413,
                 reg411,
                 reg410,
                 reg408,
                 reg407,
                 reg403,
                 reg395,
                 reg391,
                 reg390,
                 reg388,
                 reg384,
                 reg381,
                 reg379,
                 reg375,
                 reg374,
                 reg373,
                 reg371,
                 reg370,
                 reg368,
                 reg366,
                 reg364,
                 reg362,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg349,
                 reg347,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg329,
                 reg325,
                 reg310,
                 reg300,
                 reg323,
                 reg320,
                 reg317,
                 reg316,
                 reg314,
                 reg313,
                 reg309,
                 reg308,
                 reg307,
                 reg305,
                 reg296,
                 reg295,
                 reg293,
                 reg292,
                 reg290,
                 reg289,
                 reg286,
                 reg283,
                 reg277,
                 reg270,
                 reg268,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg260,
                 reg257,
                 reg250,
                 reg248,
                 reg246,
                 reg244,
                 reg243,
                 reg241,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg230,
                 reg229,
                 reg227,
                 reg212,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg216,
                 reg215,
                 reg214,
                 reg210,
                 reg207,
                 reg203,
                 reg201,
                 reg196,
                 reg172,
                 reg193,
                 reg192,
                 reg191,
                 reg189,
                 reg185,
                 reg181,
                 reg179,
                 reg178,
                 reg174,
                 reg173,
                 reg171,
                 reg169,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg161,
                 reg160,
                 reg159,
                 reg156,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg148,
                 reg147,
                 reg145,
                 reg142,
                 reg141,
                 reg138,
                 reg137,
                 reg135,
                 reg133,
                 reg132,
                 reg131,
                 reg128,
                 reg127,
                 reg123,
                 reg122,
                 reg121,
                 reg119,
                 reg117,
                 reg116,
                 reg115,
                 reg113,
                 reg112,
                 reg111,
                 reg109,
                 reg105,
                 reg104,
                 reg98,
                 reg1442,
                 reg1440,
                 reg1438,
                 forvar1436,
                 reg1432,
                 reg1429,
                 forvar1427,
                 reg1426,
                 reg1423,
                 reg1422,
                 reg1421,
                 reg1420,
                 reg1417,
                 reg1416,
                 reg1415,
                 forvar1413,
                 reg1410,
                 reg1408,
                 forvar1406,
                 reg1405,
                 reg1404,
                 reg1402,
                 reg1400,
                 reg1399,
                 reg1396,
                 reg1394,
                 reg1392,
                 forvar1390,
                 reg1389,
                 reg1387,
                 reg1384,
                 reg1383,
                 forvar1380,
                 forvar1376,
                 reg1373,
                 reg1372,
                 forvar1369,
                 forvar1368,
                 reg560,
                 reg559,
                 reg556,
                 reg554,
                 forvar549,
                 reg548,
                 forvar547,
                 reg546,
                 reg545,
                 forvar541,
                 forvar538,
                 reg537,
                 reg536,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 forvar528,
                 reg526,
                 reg516,
                 forvar515,
                 forvar513,
                 forvar511,
                 forvar504,
                 reg515,
                 forvar514,
                 reg513,
                 forvar512,
                 reg511,
                 reg509,
                 reg502,
                 reg499,
                 reg497,
                 forvar495,
                 reg494,
                 reg493,
                 reg492,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg480,
                 reg478,
                 reg477,
                 forvar476,
                 reg475,
                 reg474,
                 forvar473,
                 reg472,
                 forvar471,
                 reg469,
                 reg464,
                 reg462,
                 reg459,
                 reg458,
                 reg455,
                 forvar436,
                 reg451,
                 reg449,
                 reg447,
                 reg446,
                 reg444,
                 reg442,
                 reg438,
                 reg436,
                 reg433,
                 forvar431,
                 reg430,
                 reg429,
                 reg427,
                 reg425,
                 forvar424,
                 reg423,
                 reg422,
                 reg421,
                 reg416,
                 reg415,
                 reg414,
                 reg412,
                 reg409,
                 reg406,
                 forvar405,
                 reg404,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 forvar397,
                 reg396,
                 forvar394,
                 reg393,
                 reg392,
                 reg389,
                 forvar387,
                 reg386,
                 reg385,
                 reg380,
                 reg378,
                 forvar377,
                 reg376,
                 reg372,
                 reg369,
                 reg367,
                 forvar365,
                 forvar363,
                 forvar361,
                 reg356,
                 reg355,
                 reg350,
                 reg348,
                 reg346,
                 forvar345,
                 forvar339,
                 reg338,
                 reg333,
                 reg332,
                 reg331,
                 forvar330,
                 reg328,
                 reg327,
                 reg326,
                 forvar314,
                 forvar307,
                 reg324,
                 reg322,
                 reg321,
                 reg319,
                 reg318,
                 reg315,
                 reg312,
                 reg311,
                 forvar310,
                 reg306,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 forvar300,
                 forvar296,
                 forvar293,
                 reg299,
                 reg298,
                 reg297,
                 reg294,
                 reg291,
                 reg288,
                 reg287,
                 reg285,
                 reg284,
                 reg282,
                 reg281,
                 forvar280,
                 reg279,
                 reg278,
                 reg276,
                 forvar275,
                 forvar274,
                 reg271,
                 forvar269,
                 reg267,
                 reg261,
                 reg259,
                 reg258,
                 reg256,
                 forvar255,
                 reg254,
                 reg253,
                 forvar252,
                 reg251,
                 reg249,
                 forvar247,
                 reg245,
                 reg242,
                 reg240,
                 reg235,
                 forvar234,
                 reg233,
                 forvar232,
                 reg231,
                 reg228,
                 reg226,
                 reg225,
                 reg209,
                 forvar204,
                 forvar218,
                 reg217,
                 reg213,
                 forvar212,
                 reg211,
                 forvar209,
                 reg208,
                 reg206,
                 reg205,
                 reg204,
                 reg202,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 forvar195,
                 reg194,
                 reg190,
                 forvar188,
                 reg187,
                 reg186,
                 reg184,
                 reg183,
                 reg182,
                 forvar180,
                 reg177,
                 reg176,
                 reg175,
                 forvar172,
                 reg170,
                 reg162,
                 reg168,
                 reg163,
                 forvar162,
                 reg158,
                 reg157,
                 reg155,
                 reg154,
                 reg149,
                 reg146,
                 forvar135,
                 reg130,
                 reg144,
                 reg143,
                 reg140,
                 reg139,
                 reg136,
                 reg134,
                 forvar130,
                 reg129,
                 reg126,
                 reg125,
                 reg124,
                 reg120,
                 forvar118,
                 reg114,
                 reg110,
                 reg108,
                 reg107,
                 reg106,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 forvar99,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg98 <= ($unsigned(wire94) ?
          $unsigned($unsigned(wire97[(4'hd):(4'hd)])) : wire94[(2'h2):(2'h2)]);
      if ((~(^wire93)))
        begin
          for (forvar99 = (1'h0); (forvar99 < (1'h1)); forvar99 = (forvar99 + (1'h1)))
            begin
              reg100 = $unsigned($signed(forvar99));
              reg101 = reg100;
              reg102 = ((|$unsigned($unsigned($unsigned(wire96)))) ?
                  $signed(wire96) : wire96);
              reg103 = {(($signed((wire97 ? (8'ha6) : (8'had))) ?
                          ($unsigned((7'h51)) < (+wire94)) : $signed((reg101 && wire97))) ?
                      wire93[(3'h7):(3'h4)] : (~|(^~reg100[(3'h5):(2'h3)]))),
                  (^~(~^{wire97[(3'h7):(1'h0)], reg102[(4'hd):(4'h8)]})),
                  (reg102[(5'h14):(5'h12)] < $unsigned(reg100[(4'hb):(3'h7)]))};
              reg104 <= {($signed($signed(wire95[(1'h1):(1'h1)])) ?
                      (forvar99[(2'h3):(2'h3)] ?
                          (~^$unsigned(wire96)) : ($unsigned(reg103) ?
                              (wire97 * forvar99) : ((8'ha9) <<< wire93))) : (reg101[(4'h8):(3'h4)] * reg100)),
                  $signed($signed($unsigned($unsigned(wire96)))),
                  ({(forvar99[(3'h4):(2'h2)] && {wire96, wire95, reg102})} ?
                      (($unsigned(wire93) ? $unsigned((8'hb1)) : (+(8'ha0))) ?
                          $unsigned((wire97 <<< reg103)) : $unsigned($signed(wire96))) : forvar99)};
              reg105 <= {(((~|(forvar99 >= (8'hbf))) ?
                          reg103[(5'h14):(5'h12)] : $signed((wire93 << reg102))) ?
                      (reg100 ?
                          ((reg104 == wire97) ?
                              (reg98 ? reg102 : wire93) : {(7'h4a),
                                  wire97}) : (8'ha4)) : wire97)};
            end
        end
      else
        begin
          for (forvar99 = (1'h0); (forvar99 < (3'h5)); forvar99 = (forvar99 + (1'h1)))
            begin
              reg100 = ({wire94, reg103, wire94[(5'h12):(3'h4)]} ?
                  reg102 : reg100);
            end
          reg104 <= $signed(((((forvar99 ? reg102 : wire96) ?
                  reg105 : $unsigned(reg102)) ?
              (wire94[(4'hb):(3'h4)] >= {wire94,
                  (8'hb8)}) : (-$signed((8'hab)))) <= wire94[(5'h12):(4'he)]));
          if (wire97)
            begin
              reg105 <= wire94;
            end
          else
            begin
              reg106 = reg103[(4'h8):(1'h1)];
              reg107 = (({(~^(+reg100)), reg105[(4'hf):(3'h7)]} ?
                      ($signed($unsigned(reg102)) < (+reg105)) : (^reg102[(5'h11):(1'h0)])) ?
                  $signed((~|(~|$signed(reg101)))) : (~{(+$signed(reg106))}));
              reg108 = $signed($unsigned((reg98[(5'h13):(3'h6)] ~^ ((8'ha1) ^ {wire93,
                  wire96,
                  wire95}))));
              reg109 <= reg98[(5'h1d):(4'he)];
              reg110 = ($unsigned($unsigned($unsigned($signed(reg98)))) ?
                  wire94[(1'h0):(1'h0)] : $signed(wire97[(4'ha):(4'h9)]));
            end
          if (wire96[(5'h14):(1'h0)])
            begin
              reg111 <= (8'hb5);
            end
          else
            begin
              reg111 <= ($signed(reg103) ?
                  $signed((~((reg101 ? reg111 : reg98) | (wire93 ?
                      reg103 : wire93)))) : $unsigned(reg111));
              reg112 <= (({$signed((reg104 * wire95)),
                      reg101,
                      reg103[(5'h16):(5'h12)]} ?
                  $unsigned((reg98 <<< $unsigned(reg109))) : {($signed(wire95) ?
                          (forvar99 + wire93) : {(7'h40)}),
                      wire93,
                      reg101}) ^~ wire97);
              reg113 <= reg103[(5'h17):(4'hc)];
              reg114 = (+(-($unsigned((reg110 <<< (8'hba))) ?
                  (~(reg100 ?
                      (8'hbd) : reg109)) : ($unsigned(reg100) || {reg101,
                      reg105}))));
              reg115 <= (($unsigned((wire97[(5'h11):(4'h9)] ?
                      (^~reg104) : (~^reg98))) ?
                  {(reg110 < (reg112 ? (8'hb6) : reg107))} : (&{{reg110,
                          wire97,
                          reg111},
                      reg98,
                      (reg104 | reg106)})) == ({$unsigned(reg113[(5'h1a):(4'h8)]),
                      reg104[(4'h9):(1'h0)],
                      $signed($unsigned(reg114))} ?
                  reg101[(4'hc):(2'h2)] : ($signed($unsigned(wire94)) ?
                      ($unsigned(reg108) ?
                          ((7'h46) ?
                              reg101 : wire96) : reg112) : (&$signed(wire97)))));
              reg116 <= (&wire95[(4'ha):(3'h7)]);
            end
        end
      reg117 <= (!$signed($unsigned(reg113[(5'h1b):(5'h12)])));
      for (forvar118 = (1'h0); (forvar118 < (1'h1)); forvar118 = (forvar118 + (1'h1)))
        begin
          reg119 <= reg101[(3'h7):(3'h6)];
          reg120 = reg103;
          if ({(~&((((7'h58) >> wire95) ?
                      $unsigned(reg106) : (reg106 <<< reg105)) ?
                  ((reg116 <= reg101) ?
                      $unsigned(reg113) : $signed(wire94)) : wire94)),
              ((reg104[(1'h0):(1'h0)] - $signed((&wire95))) ^~ $unsigned(wire97[(4'hf):(4'hf)]))})
            begin
              reg121 <= wire93;
              reg122 <= ((($unsigned(reg113) > ((wire95 ?
                      wire96 : reg105) * $unsigned((7'h56)))) ?
                  ($signed((~(8'hb6))) ?
                      {wire97[(4'h8):(1'h0)]} : $signed(reg101[(4'ha):(1'h0)])) : $signed(reg119[(5'h19):(4'hf)])) <<< (reg101 ?
                  {$unsigned($unsigned(reg98))} : ((reg105[(4'he):(4'hd)] ~^ forvar99[(2'h3):(1'h1)]) <= $signed(forvar118))));
              reg123 <= $unsigned((reg115[(5'h18):(5'h15)] - (($signed(reg115) ?
                      reg119 : ((8'hb0) ? reg121 : reg105)) ?
                  reg110[(4'hd):(2'h2)] : $signed($signed(reg100)))));
            end
          else
            begin
              reg121 <= (reg113 & ((({reg119, reg113, reg103} ?
                      (~^reg110) : (reg119 ? wire96 : (7'h47))) ?
                  reg114[(4'h8):(3'h6)] : forvar118) != (~&($signed(wire94) ?
                  $signed(wire95) : reg113))));
              reg124 = $unsigned($unsigned((reg119 || reg102)));
              reg125 = (($signed((-{reg102, wire95})) | reg120) * (forvar118 ?
                  reg107[(2'h2):(1'h1)] : ($unsigned(reg101) ?
                      ($signed(reg104) || wire96) : (reg117 || $signed(forvar118)))));
            end
        end
      if ($signed((8'hb7)))
        begin
          if ((wire97 <<< $signed(reg111)))
            begin
              reg126 = (wire93 ? (&(~&reg104)) : $signed($unsigned(reg115)));
            end
          else
            begin
              reg127 <= $unsigned(($signed($unsigned($signed(reg104))) >= reg113));
              reg128 <= $unsigned(reg124);
              reg129 = ($unsigned(((-reg117[(2'h3):(2'h2)]) >>> (^(reg113 + reg121)))) ^~ $unsigned(reg116));
            end
          for (forvar130 = (1'h0); (forvar130 < (3'h6)); forvar130 = (forvar130 + (1'h1)))
            begin
              reg131 <= ((($signed((reg101 ? reg100 : wire96)) ?
                      reg101[(3'h5):(3'h5)] : $unsigned(reg102[(2'h2):(1'h1)])) ?
                  (~&$unsigned((forvar99 ?
                      reg117 : reg101))) : {forvar130[(2'h2):(1'h1)]}) && (+$signed(reg107[(1'h0):(1'h0)])));
              reg132 <= wire95;
              reg133 <= $signed(reg124);
              reg134 = (($unsigned((~&reg129)) ?
                  reg109[(2'h2):(1'h1)] : $unsigned((~&reg127[(2'h3):(1'h1)]))) != reg111[(4'h8):(2'h2)]);
              reg135 <= (($signed(reg107) & $signed({reg119[(5'h15):(1'h1)]})) ?
                  ($unsigned(reg125) ^ $signed(forvar118)) : reg132);
            end
          reg136 = wire93[(5'h12):(4'he)];
          if ($unsigned((^~({$unsigned((8'h9c)),
              $signed((8'ha4))} ^~ $unsigned((8'hab))))))
            begin
              reg137 <= $unsigned($unsigned($signed(((~reg124) ?
                  (reg122 ? wire97 : reg131) : $signed(reg135)))));
              reg138 <= reg133[(2'h2):(1'h1)];
              reg139 = reg117[(3'h5):(2'h2)];
              reg140 = (^~($signed((-(~^(7'h50)))) ^ (~&reg133)));
              reg141 <= reg135;
              reg142 <= $signed(forvar130[(3'h5):(1'h1)]);
            end
          else
            begin
              reg137 <= $signed(reg138);
              reg138 <= ({(&$unsigned((8'hbf)))} ?
                  {($signed(reg106[(4'hd):(3'h5)]) << (~^reg134))} : (&$unsigned(((reg126 | reg142) ?
                      {forvar130, reg104} : reg123))));
              reg141 <= (reg123 ?
                  reg98[(3'h5):(2'h3)] : (({(reg127 ? (8'hb5) : reg140),
                          (~^forvar118)} ?
                      (!{wire97}) : (^~(!reg102))) < (($signed((8'hb2)) ?
                      $signed(reg107) : $unsigned(forvar130)) << $unsigned((reg139 ?
                      reg125 : reg127)))));
              reg143 = reg102[(4'hf):(4'hd)];
              reg144 = (|(~(~$unsigned(reg142))));
            end
        end
      else
        begin
          if (((((reg105[(2'h3):(1'h1)] + reg119) & (8'hb7)) && (reg121[(2'h3):(2'h2)] ?
                  (7'h4e) : ({reg112, reg139, reg134} ^~ $unsigned(wire95)))) ?
              (reg109[(1'h1):(1'h1)] ?
                  wire97[(5'h12):(4'hc)] : $unsigned(((forvar99 ?
                          reg120 : (8'h9d)) ?
                      $unsigned(reg128) : reg110[(4'h8):(3'h5)]))) : (-($signed((^~reg100)) ?
                  ($signed(reg103) ?
                      $signed(reg116) : (reg138 ?
                          reg115 : reg132)) : reg107[(1'h1):(1'h1)]))))
            begin
              reg127 <= reg132[(3'h4):(2'h3)];
              reg129 = (^~reg123);
              reg130 = (~|(((7'h4e) ?
                      wire93[(5'h1c):(3'h6)] : (-(reg144 != wire93))) ?
                  $signed(reg124[(2'h2):(1'h1)]) : {(wire93[(4'ha):(3'h6)] >> (7'h52)),
                      $unsigned($unsigned(reg125))}));
              reg131 <= ((~&$signed({$unsigned(reg135)})) >>> ($unsigned((~&reg113[(2'h2):(2'h2)])) ?
                  ($unsigned((~(8'hbb))) ?
                      $unsigned((forvar118 & reg120)) : forvar99) : $unsigned((7'h4f))));
              reg134 = (^$unsigned((|(reg128 && (reg109 <= reg136)))));
            end
          else
            begin
              reg126 = (&$unsigned(({(wire95 ^ reg106)} ?
                  ($signed(reg124) ^ $unsigned((7'h4e))) : ((+reg138) == (reg114 - reg110)))));
              reg129 = reg114[(2'h2):(2'h2)];
              reg131 <= reg106;
            end
          for (forvar135 = (1'h0); (forvar135 < (3'h4)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg137 <= {$signed($unsigned($unsigned(reg117))),
                  {$signed(((reg114 ? reg116 : reg141) ?
                          $unsigned(reg112) : (reg143 == reg129)))},
                  {((reg122 == (reg113 <<< (8'hbc))) - {reg143[(1'h1):(1'h0)]}),
                      ($unsigned(reg117) == (^~(reg106 ? wire97 : reg132)))}};
              reg139 = (-reg133);
            end
          reg140 = (wire97[(4'hc):(4'hc)] ?
              (($signed((reg100 ? reg127 : reg119)) >> (reg109 <= (~&wire93))) ?
                  $signed((reg114[(2'h2):(1'h0)] ?
                      $unsigned(reg109) : reg123)) : (reg141 <<< $unsigned((reg123 ^ reg128)))) : reg121[(3'h6):(3'h6)]);
        end
    end
  always
    @(posedge clk) begin
      if (reg141[(2'h2):(1'h1)])
        begin
          if ($signed({$unsigned($unsigned((reg104 ? (8'hb0) : reg116)))}))
            begin
              reg145 <= {wire94[(5'h13):(4'hb)],
                  $unsigned(reg117[(2'h2):(1'h0)]),
                  reg98};
              reg146 = $unsigned((&$unsigned(reg104[(4'h8):(1'h0)])));
            end
          else
            begin
              reg145 <= reg119;
              reg146 = reg127[(3'h6):(3'h4)];
              reg147 <= $signed(((reg133[(1'h1):(1'h0)] >> ({reg128,
                  reg142,
                  reg138} && $signed(reg119))) < reg131));
              reg148 <= (8'hbd);
              reg149 = {(8'hb9), reg137[(3'h6):(3'h4)], reg148};
              reg150 <= reg109[(2'h2):(2'h2)];
            end
          if (reg149)
            begin
              reg151 <= reg116;
              reg152 <= reg145;
              reg153 <= $signed(((reg135 >= $unsigned({reg147,
                  (8'hbd),
                  wire94})) || $signed($unsigned((wire97 + reg147)))));
              reg154 = $signed($signed($unsigned(wire96)));
              reg155 = $signed({$unsigned(((reg141 ^ (7'h54)) ?
                      reg152[(4'ha):(4'h8)] : (!reg109)))});
            end
          else
            begin
              reg151 <= ($signed(reg109) >>> reg121);
              reg152 <= reg109;
            end
          if (wire96[(5'h11):(3'h6)])
            begin
              reg156 <= $unsigned(wire94[(3'h5):(1'h1)]);
              reg157 = reg137;
              reg158 = $unsigned($unsigned(((wire95[(4'hb):(4'h9)] - reg151) * reg154)));
            end
          else
            begin
              reg156 <= $unsigned(($unsigned(reg115) ?
                  (|((^~(8'hab)) > (^~(8'hac)))) : (-((~^reg128) < reg111))));
              reg159 <= $signed((reg157[(2'h3):(2'h2)] ?
                  reg115 : {$signed($unsigned(reg131))}));
              reg160 <= reg151;
              reg161 <= (+reg153[(4'hb):(1'h1)]);
            end
          for (forvar162 = (1'h0); (forvar162 < (2'h2)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg163 = $signed((reg115 ?
                  reg117 : {{$unsigned(reg152),
                          (reg159 && reg154),
                          wire96[(5'h14):(1'h0)]},
                      $unsigned({reg151, reg123}),
                      ($signed(reg117) - reg115[(5'h15):(5'h10)])}));
              reg164 <= (8'hb5);
              reg165 <= reg149[(4'h8):(1'h0)];
              reg166 <= (~^$unsigned(($unsigned($unsigned(wire95)) ?
                  (~$unsigned(reg98)) : reg149[(3'h6):(2'h2)])));
              reg167 <= (8'hb9);
              reg168 = (|$signed(reg157));
            end
        end
      else
        begin
          if ((+reg135[(5'h16):(5'h11)]))
            begin
              reg146 = reg161;
            end
          else
            begin
              reg145 <= reg117[(3'h4):(3'h4)];
            end
          reg149 = ((&$unsigned((^$signed(reg167)))) ?
              (reg146[(3'h5):(3'h4)] ?
                  reg121 : (reg155[(3'h4):(1'h0)] ?
                      reg113 : $unsigned(((8'ha1) ?
                          reg137 : (8'ha7))))) : (&(-($signed((8'hbe)) ^~ reg146))));
          if (((~($unsigned($signed((8'haa))) == ((|reg141) >>> (7'h52)))) && reg138))
            begin
              reg154 = reg151;
              reg156 <= $signed((&(~|$signed(reg147[(4'ha):(3'h7)]))));
              reg159 <= (reg115 ?
                  $unsigned(reg111) : (reg117[(3'h4):(1'h0)] ?
                      wire93 : (8'hb1)));
              reg162 = (({wire93[(4'he):(4'h9)], (-reg149[(3'h7):(3'h4)])} ?
                  (reg160[(5'h14):(4'hb)] >>> reg105[(3'h6):(3'h4)]) : (^(reg168[(3'h4):(2'h2)] > (reg113 > reg148)))) >>> $signed(reg166));
              reg164 <= (^($signed(reg117) ~^ {({reg121} & $unsigned(reg112))}));
              reg165 <= $unsigned({$unsigned($unsigned(reg113)),
                  $signed((8'hba)),
                  reg147[(4'hc):(4'hc)]});
            end
          else
            begin
              reg150 <= reg121;
            end
        end
      reg169 <= reg150[(5'h11):(4'hc)];
      reg170 = (&((((reg157 ? forvar162 : reg105) & (~^reg153)) ?
          (reg149 >= (reg154 ^~ reg117)) : $unsigned(((8'hbc) || reg128))) - $unsigned($signed((reg117 ?
          reg168 : reg98)))));
    end
  always
    @(posedge clk) begin
      if ({($signed($unsigned((reg165 && reg141))) ?
              $unsigned(reg111[(4'ha):(1'h0)]) : reg98),
          (reg164 ?
              $unsigned(reg160[(4'hc):(3'h5)]) : ($unsigned((wire96 ?
                      reg132 : reg142)) ?
                  ({wire96,
                      (8'ha2),
                      reg135} >>> $signed(reg151)) : reg111[(4'ha):(3'h5)]))})
        begin
          reg171 <= reg151;
          for (forvar172 = (1'h0); (forvar172 < (1'h0)); forvar172 = (forvar172 + (1'h1)))
            begin
              reg173 <= reg128;
              reg174 <= {reg131};
              reg175 = (+($signed(reg153[(1'h0):(1'h0)]) < reg145));
              reg176 = reg123[(4'h8):(3'h6)];
              reg177 = $unsigned($unsigned((|wire96[(2'h2):(2'h2)])));
              reg178 <= (&reg175[(5'h17):(4'hc)]);
            end
          reg179 <= ({reg167[(2'h2):(1'h1)]} ?
              ($signed((|(reg152 ? wire94 : wire96))) ?
                  $signed(reg135[(5'h14):(5'h14)]) : ($unsigned($unsigned(reg173)) << reg121)) : $unsigned($unsigned(wire97)));
          for (forvar180 = (1'h0); (forvar180 < (2'h3)); forvar180 = (forvar180 + (1'h1)))
            begin
              reg181 <= $unsigned($unsigned($unsigned($signed({(7'h58),
                  (7'h45)}))));
              reg182 = {reg167[(1'h1):(1'h1)],
                  (~&{(reg121 ? (~|(8'hbf)) : ((8'haf) ^ reg156))}),
                  reg105[(4'hb):(2'h3)]};
              reg183 = reg152;
              reg184 = (reg122[(5'h17):(1'h0)] ?
                  ((($signed(reg177) ? (reg152 | reg153) : $unsigned(reg98)) ?
                      reg178[(4'hc):(3'h4)] : (reg151[(4'ha):(1'h0)] * ((7'h47) ^~ reg165))) != reg164) : ($signed($signed((reg122 + reg111))) ?
                      (reg176 ?
                          forvar180 : {$unsigned(reg153)}) : $unsigned(($unsigned(reg128) * (~reg171)))));
              reg185 <= $unsigned(((!wire94) <= wire95[(3'h4):(2'h2)]));
              reg186 = reg148[(3'h4):(2'h2)];
              reg187 = reg115;
            end
          for (forvar188 = (1'h0); (forvar188 < (2'h3)); forvar188 = (forvar188 + (1'h1)))
            begin
              reg189 <= (((forvar172 - (reg156[(4'hf):(3'h4)] != (~|reg142))) >> reg184[(2'h3):(1'h0)]) ?
                  $signed({reg119, (^~((8'hac) ? (8'hbc) : reg119))}) : reg151);
              reg190 = $unsigned({reg112[(4'h8):(2'h2)],
                  $signed(((8'hb7) ?
                      reg165[(4'ha):(4'h9)] : wire93[(4'hc):(3'h5)])),
                  $unsigned(((reg131 << reg142) + (+(7'h4d))))});
              reg191 <= (reg128[(1'h1):(1'h0)] ?
                  $signed((|reg113[(3'h7):(1'h0)])) : reg177[(1'h0):(1'h0)]);
              reg192 <= (($unsigned((^~(&reg159))) != ((~reg111) ?
                  $unsigned($unsigned(reg159)) : reg148[(4'h8):(3'h7)])) != (reg123[(5'h14):(3'h5)] ?
                  (!(reg117 || reg116[(4'hd):(1'h1)])) : reg191[(3'h4):(2'h3)]));
              reg193 <= reg174[(4'hc):(2'h2)];
            end
        end
      else
        begin
          reg171 <= $unsigned($unsigned(($unsigned($signed((8'hb8))) ?
              reg179[(2'h2):(1'h1)] : {forvar172[(3'h4):(1'h1)],
                  {reg161, reg137}})));
          reg172 <= reg178[(4'he):(4'hc)];
        end
      reg194 = ($unsigned({$unsigned($signed(reg115))}) < $unsigned((^$unsigned((8'hbc)))));
      if ($signed(($signed(reg121) ?
          $unsigned(reg156) : (+({(8'haa)} != reg186[(1'h1):(1'h1)])))))
        begin
          for (forvar195 = (1'h0); (forvar195 < (1'h0)); forvar195 = (forvar195 + (1'h1)))
            begin
              reg196 <= reg178[(1'h0):(1'h0)];
              reg197 = $signed(reg152);
              reg198 = $signed($unsigned(($signed((~&(8'hb9))) ?
                  $signed((~&reg178)) : (!reg177))));
              reg199 = $unsigned(({$unsigned($signed((8'h9e))),
                      $unsigned({reg138})} ?
                  reg138[(4'ha):(2'h3)] : (^reg196)));
              reg200 = $unsigned(forvar180);
              reg201 <= reg174;
            end
          reg202 = ($signed($signed(((~|forvar180) ^ (reg186 * reg175)))) ?
              ({$unsigned((-forvar172)),
                  reg133,
                  (~&(wire97 != reg190))} >>> ({{reg200, reg183}} ?
                  (&(!reg121)) : $unsigned((wire95 || (8'hb4))))) : forvar180);
          if ($unsigned($unsigned(reg174)))
            begin
              reg203 <= $signed((&(($unsigned(reg197) < reg147) && (&reg178[(4'hf):(4'hb)]))));
            end
          else
            begin
              reg204 = reg192[(3'h5):(1'h1)];
              reg205 = (reg164 ^ (8'hb7));
              reg206 = $signed(reg189[(3'h4):(3'h4)]);
              reg207 <= (8'ha9);
              reg208 = $unsigned((7'h46));
            end
          for (forvar209 = (1'h0); (forvar209 < (3'h6)); forvar209 = (forvar209 + (1'h1)))
            begin
              reg210 <= ((($signed($signed(reg112)) ?
                      reg200[(4'ha):(3'h5)] : (8'ha5)) >= $unsigned(((~&reg119) ?
                      ((7'h51) + wire96) : (reg175 ? reg208 : reg202)))) ?
                  (!$unsigned((((7'h42) ?
                      reg174 : reg145) || reg179[(4'h9):(2'h3)]))) : (~^(reg172[(4'hc):(4'ha)] | reg182[(4'h8):(1'h1)])));
              reg211 = $signed({(~&(reg186[(1'h0):(1'h0)] >> (reg105 ?
                      reg182 : reg148)))});
            end
          for (forvar212 = (1'h0); (forvar212 < (3'h5)); forvar212 = (forvar212 + (1'h1)))
            begin
              reg213 = (reg204[(1'h0):(1'h0)] ? reg199 : {forvar212});
              reg214 <= {$unsigned(reg186)};
              reg215 <= reg185;
              reg216 <= {reg210,
                  ($unsigned({$signed((7'h52))}) ?
                      {$signed($signed(reg166))} : $signed((+reg207)))};
              reg217 = (reg204[(3'h7):(1'h1)] ?
                  $unsigned({{reg169[(1'h1):(1'h1)],
                          $unsigned((7'h54)),
                          $signed(reg187)},
                      ($signed((7'h50)) ?
                          wire95[(3'h7):(1'h0)] : {reg145, reg208})}) : reg159);
            end
          for (forvar218 = (1'h0); (forvar218 < (1'h0)); forvar218 = (forvar218 + (1'h1)))
            begin
              reg219 <= reg179[(4'h8):(2'h3)];
              reg220 <= $unsigned((reg185 ?
                  $unsigned(reg116) : {{$signed(reg175)},
                      ((reg113 <<< reg213) || {wire96})}));
              reg221 <= $unsigned(((reg115 ?
                  reg208[(3'h4):(1'h0)] : reg161[(5'h19):(3'h7)]) && $unsigned($unsigned((reg198 > reg184)))));
              reg222 <= (~$signed((^((reg187 ? reg127 : (7'h58)) || (reg182 ?
                  reg153 : reg220)))));
              reg223 <= reg142[(5'h13):(5'h11)];
              reg224 <= reg142[(4'hf):(4'hc)];
            end
        end
      else
        begin
          for (forvar195 = (1'h0); (forvar195 < (3'h5)); forvar195 = (forvar195 + (1'h1)))
            begin
              reg196 <= $signed((~|(~&$unsigned($unsigned(reg201)))));
              reg197 = reg115;
              reg198 = (7'h50);
              reg201 <= reg104;
              reg202 = $unsigned({((~&(-reg220)) ?
                      ((&reg206) && ((7'h46) ? wire96 : reg119)) : reg147)});
            end
          reg203 <= reg181[(2'h3):(1'h0)];
          for (forvar204 = (1'h0); (forvar204 < (2'h3)); forvar204 = (forvar204 + (1'h1)))
            begin
              reg207 <= {(((reg186[(2'h2):(1'h0)] ?
                          reg193[(4'hf):(2'h2)] : $unsigned(reg169)) ?
                      $signed(reg111[(3'h7):(3'h5)]) : {(reg112 ?
                              reg112 : reg217),
                          {reg204}}) >>> (((+(7'h40)) > $signed(reg197)) >= ($unsigned(reg145) == (~&reg206)))),
                  reg141[(3'h5):(3'h4)],
                  $unsigned(((|$signed(reg191)) ?
                      $signed((~reg216)) : ((reg119 ? reg173 : reg165) ?
                          $unsigned(reg133) : (~^forvar180))))};
              reg208 = $signed((~^(reg184[(4'h8):(1'h0)] < reg141)));
              reg209 = reg179;
              reg211 = (~|reg219[(1'h0):(1'h0)]);
              reg212 <= $signed(({$unsigned($signed(reg219)),
                  (~|$signed(reg105))} || $unsigned(({reg133, (8'hb7), reg133} ?
                  $signed(reg196) : (reg159 * wire96)))));
            end
          reg213 = forvar218[(4'h9):(3'h6)];
          reg214 <= (reg109 >>> (!$signed((reg177 ^~ (reg167 ?
              reg127 : reg122)))));
          reg217 = ($unsigned($signed($signed((reg221 && wire93)))) ?
              (($unsigned((reg105 ?
                      reg222 : reg179)) | (~&reg171[(3'h6):(1'h1)])) ?
                  ((reg148[(2'h3):(1'h1)] ?
                      $unsigned(forvar180) : reg207[(4'h8):(3'h6)]) >= reg141[(2'h2):(2'h2)]) : reg135[(3'h5):(2'h2)]) : $signed(($unsigned(forvar195) && $signed((reg194 && wire95)))));
          for (forvar218 = (1'h0); (forvar218 < (2'h3)); forvar218 = (forvar218 + (1'h1)))
            begin
              reg225 = $signed({{reg169}});
              reg226 = ((reg206[(1'h0):(1'h0)] ?
                      {reg117[(2'h2):(1'h1)]} : {{(reg181 | reg179)}}) ?
                  reg186 : $unsigned((^reg116[(1'h0):(1'h0)])));
              reg227 <= $unsigned($unsigned(reg197));
              reg228 = $unsigned({$signed($signed((reg216 ? reg104 : reg205))),
                  (|reg138)});
              reg229 <= ((~&$unsigned(reg169[(3'h7):(2'h2)])) ?
                  reg225[(3'h7):(2'h2)] : (reg159[(3'h6):(2'h3)] > (reg147 ?
                      $unsigned((forvar188 ?
                          reg172 : reg150)) : $signed($signed(reg161)))));
              reg230 <= {reg116, $unsigned(reg196), (-{reg177})};
              reg231 = {(($unsigned((8'had)) != ((|forvar209) - ((8'hac) || reg98))) ?
                      (reg173 ?
                          $signed(reg171[(3'h4):(1'h1)]) : $unsigned($signed(reg128))) : ((reg105[(1'h1):(1'h0)] <= (reg115 ?
                              reg196 : reg205)) ?
                          $unsigned(reg150[(3'h4):(3'h4)]) : (-reg192))),
                  ($signed(reg186) || (~reg148[(1'h1):(1'h1)])),
                  (reg189[(3'h7):(3'h4)] ?
                      reg156 : (!$signed($unsigned(reg224))))};
            end
        end
      for (forvar232 = (1'h0); (forvar232 < (2'h2)); forvar232 = (forvar232 + (1'h1)))
        begin
          reg233 = ($unsigned({reg191,
              $unsigned((reg217 ?
                  reg222 : reg123))}) & $unsigned($unsigned((reg226 | reg98[(5'h12):(3'h4)]))));
          for (forvar234 = (1'h0); (forvar234 < (1'h1)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 = (({(8'hb2)} ?
                  $unsigned({(~&wire97),
                      ((7'h4c) != reg109)}) : $signed($signed((forvar218 ?
                      wire94 : (8'had))))) | reg226);
              reg236 <= (reg233 ?
                  reg201 : ($signed(reg199) <= (((~reg231) ?
                      (forvar172 < (7'h54)) : (-forvar212)) & $signed((reg193 ?
                      reg174 : reg227)))));
            end
          if (reg183)
            begin
              reg237 <= forvar218;
              reg238 <= $signed(reg202[(4'h8):(2'h3)]);
              reg239 <= (-{reg169[(1'h0):(1'h0)]});
              reg240 = $unsigned((^(forvar195[(4'hf):(4'he)] ?
                  forvar204 : (reg123 ^~ (8'hac)))));
            end
          else
            begin
              reg240 = reg151[(3'h4):(1'h0)];
              reg241 <= reg229;
              reg242 = (($unsigned($signed($unsigned(reg220))) | $signed($unsigned(reg160))) ?
                  reg131[(3'h4):(2'h3)] : (~&reg116[(4'h8):(2'h2)]));
              reg243 <= ($unsigned(reg117) > $unsigned(reg189[(2'h2):(1'h0)]));
              reg244 <= $unsigned({{$signed($signed(forvar188)),
                      {(&reg225)},
                      reg231},
                  $signed(reg150[(5'h14):(4'h9)])});
              reg245 = $signed((reg237[(4'ha):(4'h9)] && ($unsigned($signed(reg183)) >> (+reg133))));
              reg246 <= wire93[(1'h0):(1'h0)];
            end
        end
      for (forvar247 = (1'h0); (forvar247 < (1'h1)); forvar247 = (forvar247 + (1'h1)))
        begin
          if ((^~((8'hbd) ?
              ((reg112 >>> {reg183,
                  reg202,
                  (8'hae)}) >= (~&forvar188[(3'h4):(2'h2)])) : (!((reg179 ?
                  reg117 : (7'h53)) && ((7'h40) ? reg128 : reg240))))))
            begin
              reg248 <= (~&$signed(($unsigned((-reg228)) && $signed((reg112 ?
                  (8'had) : (8'ha2))))));
            end
          else
            begin
              reg248 <= ((~^$unsigned(reg142)) * (7'h4b));
            end
        end
    end
  always
    @(posedge clk) begin
      reg249 = reg145;
      if ({$signed(wire97[(1'h0):(1'h0)]),
          (~&($signed((^reg238)) ? reg115 : (!(8'ha4)))),
          ($unsigned((^~reg246[(5'h11):(1'h1)])) ?
              reg115[(4'h9):(1'h0)] : reg172)})
        begin
          reg250 <= reg241;
        end
      else
        begin
          reg251 = reg237[(5'h13):(4'ha)];
          for (forvar252 = (1'h0); (forvar252 < (2'h2)); forvar252 = (forvar252 + (1'h1)))
            begin
              reg253 = {reg145[(3'h6):(3'h5)]};
            end
          reg254 = ({(wire95[(4'hb):(3'h5)] ?
                  $signed({reg161, reg237, reg111}) : ($signed(wire93) ?
                      $unsigned(reg248) : reg142[(1'h1):(1'h0)])),
              $signed(($signed(reg141) || (reg156 ? reg196 : reg250))),
              (reg185 ?
                  (~|(reg121 >>> reg241)) : $unsigned((reg229 >> reg253)))} <<< $unsigned($unsigned(((reg159 << wire97) ?
              (-reg238) : (!reg150)))));
          for (forvar255 = (1'h0); (forvar255 < (1'h0)); forvar255 = (forvar255 + (1'h1)))
            begin
              reg256 = $signed((-{reg248[(5'h17):(3'h6)]}));
              reg257 <= ((&{$signed($unsigned(reg164)),
                      $signed((reg138 ? reg201 : reg178))}) ?
                  ((((8'hbc) ? $signed(reg238) : $unsigned(reg251)) ?
                          reg238 : $signed($unsigned((7'h40)))) ?
                      reg253[(4'hc):(4'ha)] : $unsigned(reg221)) : {((reg116 - (~(7'h4e))) ?
                          (wire93[(2'h3):(1'h1)] ?
                              reg216[(5'h13):(1'h0)] : $unsigned(reg166)) : $signed(wire96[(4'hf):(2'h2)])),
                      $signed(reg156),
                      $signed({(|reg201),
                          ((7'h42) ? forvar255 : reg203),
                          reg181})});
            end
          if ({reg151})
            begin
              reg258 = reg236[(3'h5):(1'h1)];
              reg259 = {reg115, reg141[(5'h13):(3'h4)]};
              reg260 <= (~|(reg127[(1'h0):(1'h0)] ?
                  $signed(($signed(reg239) ?
                      reg222 : $signed(reg113))) : (~|reg229[(2'h3):(1'h1)])));
              reg261 = $unsigned($signed((((~|reg172) <<< (reg147 ^~ reg220)) ?
                  ((8'ha1) <= (|reg161)) : reg246[(3'h4):(1'h0)])));
              reg262 <= (reg250 == $signed(reg178));
              reg263 <= (^$unsigned((^(8'ha8))));
              reg264 <= (~((($signed(reg122) ?
                      (reg191 ? reg137 : reg251) : (~&reg156)) ?
                  $unsigned(reg224) : {$unsigned(wire97),
                      $unsigned(reg253),
                      $unsigned(reg171)}) >>> ($unsigned(reg166) == (reg193[(5'h10):(4'hf)] - reg237))));
            end
          else
            begin
              reg260 <= reg237;
              reg261 = reg248[(3'h5):(2'h3)];
              reg262 <= $unsigned(((!(8'hbb)) >> (reg127 ?
                  $signed((~|reg178)) : ((reg156 ? reg111 : reg122) ?
                      $unsigned(reg219) : reg236[(4'h9):(1'h0)]))));
              reg263 <= reg174[(4'h8):(3'h6)];
              reg264 <= (~|reg246[(5'h13):(2'h3)]);
              reg265 <= $unsigned($unsigned((reg196 != $signed($unsigned(reg115)))));
              reg266 <= reg203[(4'hb):(1'h1)];
            end
          reg267 = $signed((~reg254));
        end
      reg268 <= ($signed(reg259) ?
          reg267[(1'h1):(1'h1)] : (($signed(reg212) * {(reg241 <= (8'haf))}) >>> reg171));
      for (forvar269 = (1'h0); (forvar269 < (3'h5)); forvar269 = (forvar269 + (1'h1)))
        begin
          reg270 <= (((reg159 >= $signed((reg174 ?
                  (8'hbb) : (8'had)))) < $unsigned((!$unsigned(forvar255)))) ?
              (!$unsigned((reg239 ?
                  $unsigned(reg119) : ((7'h53) ?
                      (7'h47) : forvar269)))) : (~|reg241));
          reg271 = reg207;
        end
    end
  assign wire272 = $unsigned((($unsigned(reg109) ?
                       {$unsigned(reg265),
                           (reg131 ? reg138 : reg172),
                           $signed((8'hb4))} : reg137[(3'h7):(1'h1)]) ~^ (+$signed(reg222[(3'h4):(1'h1)]))));
  assign wire273 = reg222[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar274 = (1'h0); (forvar274 < (3'h4)); forvar274 = (forvar274 + (1'h1)))
        begin
          for (forvar275 = (1'h0); (forvar275 < (2'h2)); forvar275 = (forvar275 + (1'h1)))
            begin
              reg276 = reg141;
              reg277 <= (-reg179);
              reg278 = ($signed((~|(reg128[(1'h0):(1'h0)] >> (!reg246)))) ~^ (reg193 ?
                  $unsigned($unsigned({reg174,
                      reg150,
                      reg215})) : reg133[(2'h2):(1'h1)]));
              reg279 = (($unsigned(({reg196, reg220} ?
                          {reg201, reg191, reg178} : wire273[(3'h5):(1'h1)])) ?
                      ((reg105[(5'h17):(3'h6)] ?
                          reg115 : (^~reg128)) - {$signed(reg116),
                          reg191}) : $unsigned($unsigned((reg185 ~^ reg215)))) ?
                  reg137 : reg212[(2'h2):(1'h0)]);
            end
          for (forvar280 = (1'h0); (forvar280 < (2'h2)); forvar280 = (forvar280 + (1'h1)))
            begin
              reg281 = $signed((7'h4b));
              reg282 = ((^~reg123[(5'h14):(5'h13)]) >> $unsigned($unsigned((((8'hbc) ?
                  reg137 : reg266) ~^ {reg113}))));
              reg283 <= reg281;
              reg284 = ((^(~^wire95)) ?
                  {$unsigned(reg237[(3'h4):(2'h2)]),
                      $unsigned($unsigned($signed(reg165))),
                      $signed(($unsigned(reg203) ^~ $signed(reg133)))} : $signed(reg263));
              reg285 = (!$unsigned(($unsigned($unsigned((8'hb9))) || $signed((^~reg145)))));
            end
        end
      reg286 <= (reg214[(4'hd):(4'ha)] ?
          (((((8'hbe) ? reg172 : reg178) * {reg196, reg185}) ?
                  (7'h58) : reg105) ?
              reg284 : $signed((((7'h47) ? reg191 : reg138) ?
                  ((8'h9e) ?
                      reg238 : reg243) : {reg263}))) : reg116[(1'h0):(1'h0)]);
      reg287 = (7'h4c);
      reg288 = reg223[(4'he):(3'h4)];
    end
  always
    @(posedge clk) begin
      reg289 <= {reg262[(2'h2):(1'h0)]};
      reg290 <= reg220[(3'h4):(2'h2)];
      if ($unsigned($unsigned($unsigned($unsigned((reg104 ?
          reg230 : reg257))))))
        begin
          if ($signed(($signed($unsigned((wire97 || reg159))) ?
              reg174 : $unsigned($signed((reg270 < reg201))))))
            begin
              reg291 = (!reg244[(4'h8):(3'h4)]);
              reg292 <= ({$signed($signed((reg237 ? reg214 : reg174))),
                      $unsigned((reg115[(5'h17):(5'h12)] ?
                          (wire94 ? reg203 : (7'h45)) : $signed(reg171))),
                      ((^~(~&reg122)) ?
                          $unsigned($unsigned((7'h44))) : (reg135 * (8'hbe)))} ?
                  {(reg160[(1'h1):(1'h1)] ?
                          ((reg173 ? reg179 : (8'hb3)) ?
                              ((7'h41) == reg257) : (reg132 >>> (8'hab))) : $signed((reg160 ?
                              reg223 : (8'ha6))))} : reg167[(1'h1):(1'h0)]);
              reg293 <= (((~^((7'h50) <= $signed(wire273))) ?
                      (($unsigned(wire96) ? (~|reg212) : reg262) ?
                          (^$unsigned(reg112)) : reg137) : ({(~&reg147)} ?
                          reg104[(1'h1):(1'h0)] : (((7'h52) >> (8'ha7)) >> reg291[(4'hd):(2'h3)]))) ?
                  reg203[(5'h16):(5'h11)] : (wire95[(4'ha):(3'h6)] * reg98[(5'h16):(3'h7)]));
              reg294 = reg262[(4'hc):(1'h0)];
            end
          else
            begin
              reg292 <= $signed((~reg181));
              reg293 <= ((((~|(reg257 >> reg173)) * $unsigned((reg289 - (7'h4f)))) && {reg178}) >>> $unsigned($unsigned($signed((reg292 ?
                  reg105 : reg131)))));
              reg295 <= reg167;
              reg296 <= reg111;
              reg297 = reg227;
              reg298 = (~&$unsigned($signed((reg293 < {reg294}))));
              reg299 = (^((8'haa) == reg215[(4'hf):(4'ha)]));
            end
        end
      else
        begin
          reg291 = ($signed($signed((reg215[(2'h3):(2'h2)] ?
              reg192 : (reg270 ?
                  reg113 : reg248)))) > (reg298[(3'h6):(3'h4)] << (^~$unsigned(wire96[(1'h0):(1'h0)]))));
          reg292 <= reg227;
          for (forvar293 = (1'h0); (forvar293 < (1'h0)); forvar293 = (forvar293 + (1'h1)))
            begin
              reg295 <= (({{$unsigned(reg181), reg115}, reg220, reg222} ?
                  $unsigned($unsigned({reg283,
                      reg115})) : reg160) > $unsigned($unsigned(({reg257} ?
                  (reg221 ? reg191 : reg173) : $unsigned(reg145)))));
            end
          for (forvar296 = (1'h0); (forvar296 < (3'h5)); forvar296 = (forvar296 + (1'h1)))
            begin
              reg297 = {reg241,
                  (-reg236[(3'h4):(3'h4)]),
                  $unsigned((reg181[(2'h3):(2'h3)] ^ (|reg192[(4'he):(2'h3)])))};
            end
          reg298 = ((reg215[(4'hc):(3'h5)] < reg156) ?
              reg148 : reg297[(3'h4):(1'h1)]);
        end
      if (reg105[(5'h13):(4'hc)])
        begin
          for (forvar300 = (1'h0); (forvar300 < (1'h0)); forvar300 = (forvar300 + (1'h1)))
            begin
              reg301 = ($unsigned((reg164[(3'h5):(2'h2)] ?
                      ($signed(reg298) || reg277[(2'h2):(1'h1)]) : (^reg203[(3'h6):(3'h6)]))) ?
                  (({$signed(reg153), (reg98 <<< reg193)} ^~ $unsigned((reg131 ?
                          reg227 : reg164))) ?
                      reg164[(4'h9):(3'h6)] : ($signed((reg191 ^ (7'h40))) ?
                          $signed((8'hbe)) : reg201)) : (&(((reg224 < reg192) ?
                          (!reg161) : reg229) ?
                      (reg141 ?
                          ((8'ha0) ?
                              reg292 : reg263) : reg264[(3'h6):(3'h6)]) : $signed(reg296[(5'h14):(5'h11)]))));
              reg302 = reg227[(3'h5):(2'h3)];
              reg303 = ($unsigned((+(+(reg174 <= wire97)))) ?
                  reg291[(4'hb):(2'h2)] : {reg169,
                      {(~|(^~reg98)), reg133, $unsigned(reg216[(2'h3):(2'h2)])},
                      $signed(reg193)});
              reg304 = reg294[(2'h2):(1'h1)];
              reg305 <= $signed((reg161[(4'hc):(1'h1)] != (wire273 * (((7'h52) ?
                  reg173 : reg179) && $unsigned(reg189)))));
              reg306 = $unsigned($unsigned((8'ha9)));
              reg307 <= $unsigned($unsigned(wire273));
            end
          reg308 <= reg160;
          reg309 <= ($signed(reg250) << ($unsigned(reg257[(3'h4):(2'h2)]) ^ ((~|reg174) ?
              ((~&reg142) ?
                  $signed(reg266) : (reg196 <= reg263)) : (reg122[(3'h5):(1'h1)] ~^ reg263))));
          for (forvar310 = (1'h0); (forvar310 < (3'h4)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 = reg222[(1'h1):(1'h1)];
              reg312 = ($unsigned(reg178) ?
                  ((&(reg173[(1'h1):(1'h1)] ?
                      $signed(forvar296) : (^~reg294))) != (~^((^~reg112) <<< $signed(reg221)))) : {{$unsigned(reg268[(3'h7):(3'h6)]),
                          (reg290 ? $signed(reg215) : (reg265 >> reg193)),
                          reg117},
                      ({$signed(reg160),
                          {reg216, reg291, reg270},
                          $unsigned(reg123)} > reg215[(4'hd):(3'h6)])});
              reg313 <= reg161;
              reg314 <= $unsigned(wire96);
            end
          if (({$signed(($signed(reg308) ?
                  forvar300 : $signed(reg150)))} != reg151))
            begin
              reg315 = $unsigned($unsigned($signed($signed($unsigned((8'haa))))));
              reg316 <= reg306[(5'h16):(1'h1)];
            end
          else
            begin
              reg316 <= $signed($signed(({$unsigned(forvar310),
                      $signed(reg223)} ?
                  ({wire95} >> {reg116, reg312, reg161}) : ($unsigned(reg311) ?
                      {(8'hb1), reg115, reg122} : (+reg137)))));
              reg317 <= reg105[(5'h1c):(5'h1c)];
              reg318 = reg238[(4'h8):(3'h6)];
              reg319 = $unsigned(reg169);
            end
          if ((reg263[(3'h4):(1'h0)] ?
              reg174[(3'h4):(3'h4)] : $signed(forvar300[(3'h6):(2'h3)])))
            begin
              reg320 <= ((($signed(reg246[(5'h14):(1'h0)]) ?
                      ($unsigned(wire272) ?
                          (reg238 ?
                              reg222 : (8'ha2)) : reg141[(5'h11):(2'h2)]) : $signed(reg215[(1'h0):(1'h0)])) ?
                  ($unsigned($unsigned(reg312)) << (+$signed(reg189))) : reg203) << (~|reg297[(5'h12):(4'h9)]));
            end
          else
            begin
              reg321 = reg236[(4'he):(4'hd)];
              reg322 = reg210[(4'h8):(3'h7)];
              reg323 <= $unsigned(($unsigned($unsigned((reg166 ~^ (8'ha8)))) && $signed((~|(reg137 && reg304)))));
              reg324 = reg296[(4'hf):(3'h7)];
            end
        end
      else
        begin
          if ((-$signed((reg222[(1'h0):(1'h0)] >> $unsigned((reg207 && reg135))))))
            begin
              reg300 <= (|$unsigned(reg230[(3'h5):(3'h5)]));
              reg301 = wire273;
              reg302 = $unsigned($signed($unsigned(((~^reg161) == (^reg298)))));
              reg305 <= $unsigned((-$signed(reg117)));
            end
          else
            begin
              reg301 = (8'hbf);
            end
          reg306 = $unsigned($unsigned($signed($unsigned(reg138))));
          for (forvar307 = (1'h0); (forvar307 < (3'h5)); forvar307 = (forvar307 + (1'h1)))
            begin
              reg308 <= $signed(($signed(reg283) ?
                  {((~reg311) ?
                          reg244[(4'h8):(3'h4)] : $signed(reg166))} : (-wire95)));
              reg309 <= ($signed((~reg311[(4'hc):(4'ha)])) || $signed($signed($signed((reg105 >>> reg167)))));
              reg310 <= (!(~^reg159));
            end
          reg313 <= reg277[(2'h2):(1'h0)];
          for (forvar314 = (1'h0); (forvar314 < (3'h5)); forvar314 = (forvar314 + (1'h1)))
            begin
              reg316 <= reg302[(4'h8):(3'h5)];
              reg318 = reg294[(2'h3):(2'h3)];
            end
          if ($signed({(reg302 <<< ((reg201 ? reg296 : (8'hb6)) - wire97)),
              {$unsigned($signed(reg191))},
              (8'h9f)}))
            begin
              reg320 <= $unsigned(reg201[(2'h2):(2'h2)]);
              reg323 <= (^~$signed($signed((~|reg323[(1'h1):(1'h0)]))));
              reg325 <= (reg306 ?
                  reg246[(1'h1):(1'h0)] : reg227[(5'h18):(1'h0)]);
              reg326 = $signed((!(reg248 & (!(forvar293 < reg309)))));
              reg327 = (^(|$signed((~(~&reg111)))));
              reg328 = (reg132[(2'h2):(2'h2)] <= $signed((($unsigned(reg153) ?
                      ((8'ha4) ^~ (8'hbd)) : (reg246 < reg171)) ?
                  $unsigned($unsigned(reg270)) : (reg210 || forvar310[(4'hc):(3'h6)]))));
              reg329 <= reg320;
            end
          else
            begin
              reg319 = (~&(~((~|{reg243, reg329}) ^ $signed((reg223 ?
                  reg138 : reg221)))));
              reg320 <= {reg215};
              reg323 <= (^({($signed(reg322) - $unsigned((7'h55)))} >= $unsigned(reg250[(1'h0):(1'h0)])));
              reg324 = $signed($signed(reg152[(4'ha):(1'h1)]));
              reg326 = $signed({{({reg323} ? (~&reg167) : (7'h51))},
                  ({(|reg266), $signed(forvar307)} == reg238[(4'ha):(2'h3)])});
            end
        end
      for (forvar330 = (1'h0); (forvar330 < (3'h5)); forvar330 = (forvar330 + (1'h1)))
        begin
          if (reg238[(3'h5):(2'h3)])
            begin
              reg331 = (reg196 ?
                  (~&(-$unsigned(reg133))) : $unsigned((((~|(8'hb9)) ?
                          reg250[(4'hb):(2'h3)] : reg324) ?
                      reg166[(3'h4):(2'h2)] : ((+reg327) & $unsigned(reg298)))));
              reg332 = $signed($unsigned(($unsigned($unsigned(forvar307)) ?
                  reg127[(3'h7):(3'h4)] : (~|reg265))));
              reg333 = reg179;
            end
          else
            begin
              reg334 <= {(^~$signed($signed(reg310))),
                  (+(!({reg172, reg315, reg241} + (!reg323))))};
              reg335 <= $signed(((7'h4b) ?
                  reg260[(4'h9):(3'h5)] : reg135[(3'h4):(2'h3)]));
              reg336 <= {(~reg192),
                  ((reg305[(3'h5):(2'h3)] + $unsigned((+reg310))) ?
                      (8'ha6) : (reg98[(2'h3):(1'h1)] + ((wire273 == reg250) ?
                          reg291[(3'h5):(1'h0)] : (reg293 >= reg111)))),
                  reg291[(4'he):(4'h9)]};
              reg337 <= (+$unsigned((((reg248 >> (8'hb9)) ?
                  (forvar330 << reg224) : $unsigned(reg173)) && reg147)));
              reg338 = ($unsigned(((^{(8'haa), wire95, reg332}) ?
                      ($signed(reg171) <= (reg266 << wire272)) : (((8'h9c) ?
                          reg230 : reg167) & (reg151 ? reg127 : forvar330)))) ?
                  reg250 : $unsigned(reg201));
            end
          for (forvar339 = (1'h0); (forvar339 < (3'h5)); forvar339 = (forvar339 + (1'h1)))
            begin
              reg340 <= (7'h49);
              reg341 <= (^(-((reg223[(3'h7):(2'h2)] > (reg336 ?
                      reg295 : reg164)) ?
                  $signed({(7'h45), reg207}) : {$signed(reg214),
                      (reg236 ~^ reg141),
                      reg142[(4'h9):(3'h6)]})));
              reg342 <= reg301[(4'h8):(3'h7)];
              reg343 <= reg306[(3'h7):(3'h7)];
            end
          reg344 <= reg137;
          for (forvar345 = (1'h0); (forvar345 < (3'h5)); forvar345 = (forvar345 + (1'h1)))
            begin
              reg346 = reg98[(3'h6):(1'h0)];
              reg347 <= (&$unsigned($unsigned(reg210)));
              reg348 = $unsigned(forvar310);
              reg349 <= {(7'h40)};
              reg350 = $signed({(reg332 <= $unsigned(reg317[(3'h7):(2'h3)])),
                  $signed($signed($unsigned(reg227)))});
              reg351 <= reg342;
            end
          reg352 <= (8'h9f);
          if ((~^({$signed((forvar300 ? reg343 : (8'hab)))} ?
              {reg297, $unsigned((reg265 ? reg297 : reg325))} : (8'h9f))))
            begin
              reg353 <= reg323;
              reg354 <= $unsigned(reg349);
              reg355 = reg243;
              reg356 = wire94[(1'h0):(1'h0)];
              reg357 <= ((^reg277) + (^~reg295));
              reg358 <= ($unsigned($signed(({reg266} ?
                  reg221 : reg167))) <= $unsigned($unsigned(reg250[(4'hd):(1'h1)])));
              reg359 <= (~&$signed(reg295));
            end
          else
            begin
              reg353 <= (((~{(~reg128), (8'hbb), reg333}) ?
                  $signed((~^$signed(reg338))) : (reg142[(5'h10):(3'h6)] && ((reg151 ?
                          reg301 : reg196) ?
                      reg142 : (&reg223)))) < reg207[(4'he):(4'ha)]);
              reg355 = $signed($signed((7'h58)));
              reg356 = {((reg312[(3'h7):(2'h2)] < $signed(reg348[(1'h1):(1'h1)])) ?
                      reg178 : $signed((~(wire273 == (8'ha0))))),
                  (7'h51),
                  (reg328[(1'h0):(1'h0)] ?
                      (8'hb5) : (-{reg296[(5'h1b):(5'h1b)]}))};
              reg357 <= reg352[(4'hb):(4'hb)];
              reg358 <= {((|$unsigned(reg248[(2'h3):(1'h1)])) != (~|(&forvar296))),
                  ({reg248} ~^ ({{(8'hbc)}} ?
                      ({reg165, (7'h4f)} > reg313) : reg311))};
              reg359 <= reg326;
            end
        end
      reg360 <= forvar307;
      for (forvar361 = (1'h0); (forvar361 < (2'h3)); forvar361 = (forvar361 + (1'h1)))
        begin
          reg362 <= $unsigned(($unsigned($signed($unsigned(reg117))) ?
              reg112 : (~|{reg222[(3'h6):(1'h0)]})));
          for (forvar363 = (1'h0); (forvar363 < (2'h3)); forvar363 = (forvar363 + (1'h1)))
            begin
              reg364 <= (reg346 || (reg263[(2'h3):(1'h1)] ?
                  (((reg291 != reg250) == (reg309 ? reg133 : (8'hb5))) ?
                      reg329[(5'h19):(3'h5)] : ((~|reg222) <= $unsigned(reg178))) : reg305));
            end
          for (forvar365 = (1'h0); (forvar365 < (1'h0)); forvar365 = (forvar365 + (1'h1)))
            begin
              reg366 <= {(|((^~(reg323 - reg334)) ?
                      reg189 : (reg220 ~^ ((8'ha1) < (7'h43))))),
                  $unsigned(wire95[(2'h3):(1'h0)]),
                  reg219[(5'h1b):(5'h16)]};
              reg367 = (reg313[(3'h7):(1'h1)] ?
                  ((8'ha3) <<< $unsigned((~^reg141))) : (^~{(-$signed(reg181))}));
              reg368 <= $signed($unsigned((reg174 == (!(&reg304)))));
            end
          if ($unsigned((reg243 ?
              (((reg117 ? reg296 : reg178) || (reg332 << forvar293)) ?
                  $signed((~|reg216)) : reg270[(3'h6):(2'h2)]) : (8'hb8))))
            begin
              reg369 = reg354;
            end
          else
            begin
              reg370 <= wire95[(3'h6):(3'h4)];
              reg371 <= $signed($unsigned((((reg221 ? reg147 : (7'h54)) ?
                  (reg164 ?
                      reg171 : reg148) : reg229[(2'h2):(1'h1)]) > reg201)));
            end
          if ((reg227[(3'h5):(3'h4)] ?
              (~|(-($unsigned(reg152) >> $unsigned(reg343)))) : (^{(8'hb3),
                  reg159[(1'h1):(1'h0)]})))
            begin
              reg372 = (-{$signed(((reg243 ? (7'h44) : (7'h50)) > (reg135 ?
                      reg221 : reg246)))});
              reg373 <= (reg270[(4'he):(4'ha)] ?
                  $signed(reg227) : ({reg230[(2'h3):(1'h1)],
                          (reg150[(3'h7):(1'h0)] ?
                              (reg123 ? reg340 : reg270) : (|reg353)),
                          reg353} ?
                      (~|$signed(reg298[(4'hf):(3'h4)])) : $unsigned((reg127[(4'h8):(2'h3)] ?
                          (reg167 + wire96) : (~|(7'h49))))));
              reg374 <= $signed(({$signed(reg248[(4'h9):(2'h2)])} << ($unsigned(wire93) >>> (~&reg370))));
              reg375 <= $unsigned((&((8'ha7) >= reg223)));
              reg376 = reg257[(3'h5):(1'h1)];
            end
          else
            begin
              reg372 = $unsigned($unsigned($signed($signed((reg299 ?
                  reg257 : reg324)))));
            end
          for (forvar377 = (1'h0); (forvar377 < (3'h5)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg378 = reg289;
              reg379 <= reg324[(3'h6):(3'h6)];
              reg380 = (+$unsigned((((8'h9f) ?
                  (reg378 ? reg333 : reg379) : (wire96 ^~ (8'ha3))) > reg352)));
            end
          reg381 <= reg338[(1'h0):(1'h0)];
        end
    end
  assign wire382 = (-$signed(reg238[(1'h1):(1'h0)]));
  assign wire383 = (($signed($unsigned({reg137, reg210})) ?
                           (!$unsigned((!reg265))) : reg148[(3'h6):(3'h6)]) ?
                       reg127[(1'h0):(1'h0)] : $signed(reg374[(4'hd):(2'h3)]));
  always
    @(posedge clk) begin
      reg384 <= (8'hb4);
      reg385 = $signed(($signed(reg375) | $signed(reg214)));
      reg386 = {reg268[(2'h3):(1'h0)],
          ($signed(reg165) - (+$unsigned(reg173)))};
      for (forvar387 = (1'h0); (forvar387 < (2'h3)); forvar387 = (forvar387 + (1'h1)))
        begin
          reg388 <= reg121;
          if ($unsigned((|(((8'ha5) && ((8'hbd) || reg305)) ?
              $unsigned(((7'h50) ~^ reg123)) : (((7'h4b) ? reg142 : reg354) ?
                  {reg266} : reg127)))))
            begin
              reg389 = reg147;
              reg390 <= reg150;
              reg391 <= $signed((($unsigned(reg300[(3'h4):(1'h1)]) ?
                  $signed(reg308) : ((8'haf) ?
                      $unsigned(reg174) : (~|reg230))) >= {(&reg385[(3'h5):(1'h0)]),
                  reg359[(1'h0):(1'h0)]}));
            end
          else
            begin
              reg390 <= reg246;
              reg392 = ({(reg289[(5'h15):(2'h2)] * reg307[(3'h7):(3'h6)]),
                      wire94} ?
                  ($unsigned($signed($unsigned(reg374))) != reg334) : $signed((reg221 | reg210[(3'h5):(2'h2)])));
              reg393 = $signed($unsigned(($signed(reg156[(5'h13):(2'h2)]) * $unsigned(reg358[(4'hb):(4'ha)]))));
            end
          for (forvar394 = (1'h0); (forvar394 < (1'h0)); forvar394 = (forvar394 + (1'h1)))
            begin
              reg395 <= reg379;
              reg396 = reg353;
            end
          for (forvar397 = (1'h0); (forvar397 < (2'h2)); forvar397 = (forvar397 + (1'h1)))
            begin
              reg398 = $unsigned($signed(((~&(reg310 & reg214)) ?
                  ($signed(reg293) ? (7'h51) : $unsigned(reg309)) : (reg207 ?
                      (reg305 != reg366) : (8'ha2)))));
              reg399 = $unsigned(reg289[(4'hb):(3'h4)]);
              reg400 = reg148;
              reg401 = reg112;
              reg402 = reg364;
              reg403 <= reg265;
            end
          reg404 = reg223[(4'hf):(4'hc)];
          for (forvar405 = (1'h0); (forvar405 < (3'h4)); forvar405 = (forvar405 + (1'h1)))
            begin
              reg406 = $signed({($unsigned($signed(reg112)) ?
                      reg389 : ((reg185 >>> reg379) ?
                          $unsigned(reg398) : (reg340 ?
                              (7'h41) : forvar394)))});
            end
        end
      reg407 <= ($unsigned($signed((((8'hae) ? (7'h58) : (8'hbc)) ?
              reg229[(3'h5):(3'h4)] : $signed(reg112)))) ?
          {(^$signed(reg142)),
              ((7'h50) ?
                  $signed((~reg128)) : $signed($unsigned(reg239)))} : $unsigned(({(reg223 ^ reg309)} ?
              $unsigned($unsigned(reg404)) : $signed($signed(reg141)))));
      if (reg403)
        begin
          if (reg343[(3'h5):(3'h4)])
            begin
              reg408 <= $unsigned((-$unsigned((7'h4d))));
              reg409 = $signed((^reg222[(3'h6):(3'h4)]));
              reg410 <= ($signed((~&$unsigned((reg313 | reg156)))) > reg354);
            end
          else
            begin
              reg409 = $unsigned({reg185[(4'h9):(3'h5)],
                  (7'h55),
                  $unsigned(((-reg246) ?
                      (reg352 || (8'hae)) : {reg323, reg347, reg374}))});
              reg410 <= {$signed((-(((7'h48) ?
                      reg357 : reg128) ~^ reg308[(5'h10):(1'h1)]))),
                  reg263,
                  ($unsigned($signed($signed(reg229))) != {((reg203 ?
                              reg121 : reg395) ?
                          (7'h4c) : reg164[(4'h8):(4'h8)]),
                      (reg401 ? reg116 : (~&reg389))})};
              reg411 <= (7'h4d);
              reg412 = (|(((^(+reg373)) >> (reg381[(2'h2):(1'h0)] != $unsigned(reg189))) & $signed(((^~(7'h56)) ?
                  reg181[(5'h11):(4'hd)] : {(8'ha9)}))));
              reg413 <= $unsigned(wire273);
            end
          if ((reg406 | $signed(reg145)))
            begin
              reg414 = reg191;
              reg415 = reg219;
              reg416 = $signed(($unsigned($unsigned((reg151 | reg212))) | (reg98[(4'h8):(2'h2)] && ((reg224 && reg371) ?
                  $signed(reg352) : reg342))));
              reg417 <= $signed(reg263[(3'h7):(2'h2)]);
              reg418 <= ({reg305,
                  (~&reg370),
                  {($signed(reg150) ?
                          (reg179 ~^ reg358) : (reg395 * (8'hb1)))}} + ({($unsigned(wire94) & $signed(reg151)),
                      $signed($signed((7'h51))),
                      {reg353[(3'h4):(1'h0)]}} ?
                  $unsigned((8'hba)) : ($unsigned((reg147 ? reg214 : reg370)) ?
                      $signed((7'h49)) : ((reg171 ?
                          (7'h54) : wire97) == (~reg147)))));
              reg419 <= (reg290[(1'h0):(1'h0)] ?
                  (~|(~($unsigned(reg160) + $signed(reg121)))) : $unsigned(($unsigned((reg337 ?
                          reg238 : (8'hbe))) ?
                      (^~(reg210 ?
                          reg295 : reg244)) : $signed((wire96 > reg368)))));
              reg420 <= ((reg181[(2'h3):(2'h2)] ?
                  (reg398 >>> ($signed(reg359) ?
                      (reg257 ?
                          reg268 : reg223) : reg313)) : $signed(reg141)) >> $unsigned(reg408[(4'h9):(1'h1)]));
            end
          else
            begin
              reg414 = $unsigned(reg113);
              reg417 <= reg400[(4'hc):(3'h4)];
              reg421 = (reg174[(1'h1):(1'h1)] ? (!reg314) : reg296);
              reg422 = ({{reg227[(5'h14):(5'h11)]}} >= reg320[(4'hd):(3'h6)]);
            end
          reg423 = {(((~&$unsigned((8'hac))) | ($unsigned((8'hae)) ^~ $signed((8'haf)))) ?
                  (-$signed((~^reg116))) : ($signed($unsigned(reg196)) ?
                      reg402 : $signed($signed(reg215))))};
          for (forvar424 = (1'h0); (forvar424 < (2'h2)); forvar424 = (forvar424 + (1'h1)))
            begin
              reg425 = reg296;
              reg426 <= $unsigned((~{$unsigned(reg196),
                  reg395[(3'h4):(2'h3)],
                  (7'h54)}));
              reg427 = ($signed($unsigned((~|(7'h4a)))) > $signed((&wire273[(2'h3):(2'h2)])));
              reg428 <= $unsigned((&(((reg178 ?
                      reg347 : wire93) - $signed(reg277)) ?
                  (reg115[(5'h14):(3'h4)] ?
                      reg212 : (reg286 <<< wire94)) : reg219)));
              reg429 = ($signed(($signed({wire93,
                      reg402,
                      reg316}) == (!reg219))) ?
                  reg215 : $signed(reg373[(3'h6):(2'h3)]));
              reg430 = ((($unsigned($unsigned((8'hbb))) ?
                      reg429 : reg335) <<< {$unsigned($unsigned(reg138)),
                      $unsigned((~|forvar397))}) ?
                  $signed($signed($signed($signed(reg212)))) : (~(($unsigned(reg399) ~^ reg112) ?
                      (^(reg310 <= reg415)) : ((~^reg379) > (reg353 | reg401)))));
            end
          for (forvar431 = (1'h0); (forvar431 < (2'h2)); forvar431 = (forvar431 + (1'h1)))
            begin
              reg432 <= reg349[(3'h7):(2'h2)];
              reg433 = reg214;
              reg434 <= (($unsigned(reg409) <= (reg185[(3'h5):(3'h5)] ?
                      $signed((reg212 ?
                          wire383 : (8'hb7))) : $unsigned(reg351[(3'h5):(1'h0)]))) ?
                  {reg160,
                      reg317,
                      $unsigned(($signed(reg115) ?
                          reg308 : $unsigned(reg416)))} : $unsigned(wire96[(2'h2):(1'h0)]));
            end
        end
      else
        begin
          if ($signed(((8'ha3) ?
              ((-reg296[(3'h5):(2'h2)]) ?
                  $unsigned((^~reg224)) : (((8'ha5) << reg349) * $unsigned(forvar424))) : ($signed(((7'h43) ?
                  reg393 : reg412)) > $signed(reg193)))))
            begin
              reg409 = reg433[(4'h8):(2'h2)];
              reg412 = reg420[(1'h1):(1'h1)];
              reg413 <= $unsigned($unsigned(reg292[(2'h2):(1'h0)]));
            end
          else
            begin
              reg409 = $signed((~$unsigned($signed($unsigned(wire273)))));
              reg410 <= ((reg334 ?
                      (reg359[(1'h0):(1'h0)] << (8'ha2)) : $unsigned((~reg357))) ?
                  ($signed((^~$unsigned(reg237))) || (|reg357)) : (|{reg113[(5'h16):(3'h4)]}));
              reg412 = $unsigned($unsigned((8'ha2)));
            end
          if ({$signed($unsigned(reg386[(3'h7):(1'h1)])),
              (~|$unsigned((reg342[(3'h5):(2'h3)] ?
                  (^reg398) : ((8'ha1) ? reg392 : reg340)))),
              $signed($signed({(reg265 * reg153),
                  (reg270 << (8'ha5)),
                  $signed((7'h4b))}))})
            begin
              reg417 <= reg191[(2'h2):(1'h0)];
              reg418 <= (((((!reg428) >>> reg215[(2'h3):(2'h3)]) ?
                      $unsigned((reg221 < reg409)) : (7'h53)) ?
                  $signed(reg334) : ((|(reg229 ? reg433 : reg260)) ?
                      reg181 : {(|reg335)})) == reg227[(5'h16):(4'ha)]);
            end
          else
            begin
              reg414 = reg290[(2'h2):(1'h0)];
              reg415 = $signed((8'hb3));
            end
        end
    end
  assign wire435 = reg341[(4'he):(4'h9)];
  always
    @(posedge clk) begin
      if (((reg337 ?
              (($unsigned(wire97) ?
                  (-reg227) : {(8'hb9),
                      reg413,
                      (7'h4d)}) >> $signed($unsigned(reg224))) : reg264) ?
          $signed(($unsigned($unsigned((8'hb9))) & ((&reg133) >= (reg417 ?
              reg142 : reg368)))) : (7'h4d)))
        begin
          reg436 = $signed($signed((~|$signed((reg137 ? reg156 : reg98)))));
          reg437 <= (!(((reg334 >= reg109) ?
                  ({reg145,
                      reg221,
                      reg241} ^~ (~|reg374)) : $unsigned($signed(reg192))) ?
              reg374 : (!{$unsigned((8'ha8)), (reg122 ? reg270 : (7'h52))})));
          if ($unsigned((~(((8'ha9) <= reg109[(3'h4):(1'h1)]) || reg216[(2'h3):(2'h3)]))))
            begin
              reg438 = (~((reg105 == ((wire435 ? reg123 : reg207) ?
                  reg148 : reg381[(1'h0):(1'h0)])) != $signed(reg335)));
              reg439 <= ((~reg138) <= {(~^reg189)});
              reg440 <= $unsigned(reg104);
              reg441 <= (^(+reg207));
              reg442 = reg248;
              reg443 <= $signed($unsigned({reg300}));
              reg444 = (((8'hae) != $signed((~^{reg266, (8'h9c), reg357}))) ?
                  {reg334[(1'h0):(1'h0)],
                      (7'h4f),
                      ($signed((reg309 ^~ (7'h51))) < (~&(+reg268)))} : reg417);
            end
          else
            begin
              reg439 <= $signed((($unsigned(((8'ha9) != reg104)) << reg244[(3'h5):(3'h4)]) - reg174));
              reg442 = reg343;
            end
          if (reg196)
            begin
              reg445 <= ($unsigned($signed({(|reg243),
                  (~|reg212)})) ^~ ($unsigned($signed({reg296,
                  reg131,
                  reg353})) < reg133[(2'h2):(1'h1)]));
              reg446 = reg216;
              reg447 = $signed((($signed($unsigned(reg320)) << (^~(reg440 ?
                      reg98 : reg351))) ?
                  $unsigned(({reg141,
                      reg248,
                      (8'ha3)} + $unsigned(reg191))) : $signed({{reg250},
                      (+wire435)})));
            end
          else
            begin
              reg445 <= $signed($unsigned($signed(reg351)));
              reg446 = $signed(reg220[(2'h2):(1'h1)]);
              reg448 <= reg227;
              reg449 = ($signed(({$unsigned(reg289)} >= ((reg434 ?
                      reg411 : reg138) ~^ (|reg362)))) ?
                  (~&$signed(($signed(reg329) ?
                      reg413 : $unsigned(reg305)))) : reg147[(3'h5):(3'h4)]);
              reg450 <= (+(({reg116[(3'h5):(3'h4)]} ?
                      (((8'haa) ? reg384 : reg142) != (reg359 ?
                          (8'ha8) : reg309)) : {$signed(reg216)}) ?
                  {$unsigned($signed(wire96)),
                      $unsigned((-reg241))} : (+reg221)));
              reg451 = {$signed(wire272[(3'h4):(2'h3)])};
            end
        end
      else
        begin
          for (forvar436 = (1'h0); (forvar436 < (3'h5)); forvar436 = (forvar436 + (1'h1)))
            begin
              reg437 <= (|$signed(($unsigned((reg270 ?
                  reg260 : wire93)) << ((reg357 ? reg172 : reg153) ?
                  $signed(reg165) : reg352[(4'h8):(3'h4)]))));
              reg438 = reg127[(3'h5):(3'h5)];
              reg442 = (reg266 ?
                  (&(&$signed((reg216 | (8'hbf))))) : ((8'hb6) > reg260[(3'h4):(1'h1)]));
              reg444 = (^reg428);
              reg445 <= $unsigned(reg270[(1'h0):(1'h0)]);
              reg448 <= ($signed((~&$signed({reg128,
                  reg283}))) >>> (+$signed(reg413)));
            end
          reg449 = (($unsigned($signed((~|reg375))) ?
              $signed(wire435) : reg336[(5'h14):(5'h14)]) || reg283[(4'he):(2'h2)]);
          if (reg323[(4'hf):(4'hd)])
            begin
              reg451 = $unsigned((reg410 & $signed((reg407[(1'h1):(1'h0)] ?
                  $signed(reg191) : forvar436[(3'h6):(2'h2)]))));
            end
          else
            begin
              reg451 = $signed(wire272);
              reg452 <= ({reg265,
                  (({reg119} ?
                          reg169[(4'hd):(2'h2)] : ((8'ha0) ? reg428 : reg127)) ?
                      ((~|reg323) ?
                          $unsigned(reg142) : (reg381 < reg222)) : reg192[(4'h8):(3'h5)]),
                  $signed({(reg381 ? (7'h41) : reg207)})} << (({((7'h42) ?
                          wire95 : reg292),
                      $signed(reg128)} ?
                  $unsigned($signed((8'hbd))) : {{reg207,
                          reg159,
                          reg104}}) < ({(reg448 & reg105)} ?
                  $signed((reg268 >= reg309)) : (reg222 >> $signed((8'hbf))))));
              reg453 <= $unsigned((((reg104 ^~ reg384) >> reg354) ?
                  (8'hb5) : $unsigned((~&(8'hb8)))));
            end
          reg454 <= reg364;
          if (((-$signed({$unsigned(reg310),
              reg320[(3'h5):(1'h1)]})) ^~ $unsigned(((8'h9f) | (reg171 ?
              $signed(reg111) : $signed((8'ha8)))))))
            begin
              reg455 = reg153[(4'h9):(4'h9)];
              reg456 <= reg147[(4'h8):(3'h4)];
              reg457 <= (!({$signed({reg359, reg257})} ?
                  (&$unsigned($unsigned(reg449))) : ($signed($unsigned(reg344)) && $unsigned((wire95 == reg263)))));
              reg458 = $unsigned((&$unsigned($unsigned($signed(reg116)))));
              reg459 = (~^wire93);
              reg460 <= ({({(7'h4d)} != reg98[(5'h1e):(5'h19)])} > ((((reg220 ?
                          wire94 : (8'h9e)) ?
                      ((7'h49) ? reg212 : reg344) : (^~reg444)) ?
                  (reg434 ?
                      $unsigned(reg391) : (|reg420)) : $unsigned(reg128[(3'h4):(2'h3)])) * ({(^reg221),
                      $unsigned(wire435)} ?
                  (~|reg229) : ($unsigned(reg260) ?
                      (|reg215) : $signed(reg391)))));
            end
          else
            begin
              reg456 <= {reg138, reg349, reg289};
              reg458 = (~&reg283);
              reg460 <= (^~$unsigned(reg132));
              reg461 <= $unsigned((^reg224));
              reg462 = $unsigned(reg203[(3'h6):(3'h6)]);
            end
          if (reg381)
            begin
              reg463 <= (~|($unsigned($signed((reg147 > reg314))) ?
                  (^~($signed(reg250) ?
                      {reg417,
                          (7'h49)} : reg148[(2'h2):(2'h2)])) : (reg418 >> (reg220 ?
                      reg215[(3'h7):(3'h6)] : wire272[(3'h4):(1'h0)]))));
              reg464 = reg375[(3'h6):(3'h6)];
              reg465 <= (((reg262 ?
                          (&(reg122 ?
                              (8'ha9) : reg246)) : $signed((reg153 ^~ reg352))) ?
                      $unsigned(($signed(reg359) ?
                          (8'h9e) : (reg349 ?
                              reg189 : (7'h45)))) : reg239[(3'h5):(3'h4)]) ?
                  reg109[(1'h0):(1'h0)] : (wire93[(5'h15):(4'h8)] || reg439[(4'he):(3'h4)]));
              reg466 <= $signed(($unsigned({$unsigned(reg335),
                  $signed(reg403)}) || $signed({$unsigned(reg390),
                  {(8'hac), reg323, (7'h47)}})));
            end
          else
            begin
              reg463 <= ($signed((-(reg447[(2'h3):(2'h2)] ?
                      {reg262, reg445} : (8'hac)))) ?
                  (^{$signed((~^reg417)),
                      (-$unsigned(reg335))}) : (((~|(reg457 ?
                          reg354 : reg362)) ?
                      ((~reg236) ?
                          reg419 : reg260[(4'ha):(1'h0)]) : reg442[(4'hc):(3'h7)]) >> $signed($unsigned(reg391[(2'h2):(1'h0)]))));
              reg464 = $signed(reg173);
            end
          if (($signed($unsigned(((-reg413) ~^ $unsigned((8'hbc))))) ?
              ((8'ha0) ? reg248 : $signed((~{reg147}))) : reg308))
            begin
              reg467 <= reg152;
            end
          else
            begin
              reg467 <= ($unsigned((((reg132 ? (8'hae) : reg222) ?
                          (reg266 ? (8'ha0) : reg160) : (reg201 ^ reg219)) ?
                      (reg243 >= (^reg438)) : (reg413 <= (wire272 ?
                          (7'h53) : reg145)))) ?
                  reg119[(4'hf):(4'he)] : (~$unsigned((7'h47))));
              reg468 <= $signed(((($unsigned(wire97) <<< (8'ha5)) * (reg296[(4'hc):(4'ha)] ?
                  $signed(reg257) : reg244[(1'h1):(1'h1)])) + (~^reg354)));
              reg469 = reg466;
              reg470 <= $unsigned({$unsigned({$signed(reg207),
                      ((7'h48) ? reg138 : reg262)}),
                  {(-$signed(reg166)), reg161[(4'h9):(4'h9)]},
                  (-((~^reg212) ? (reg201 * reg456) : reg138))});
            end
        end
      for (forvar471 = (1'h0); (forvar471 < (3'h4)); forvar471 = (forvar471 + (1'h1)))
        begin
          reg472 = ((reg156 | $signed($signed(((8'hbf) ? reg131 : reg268)))) ?
              (~|(^($unsigned(reg457) ?
                  ((7'h43) ?
                      reg174 : reg323) : $unsigned(reg447)))) : (~^(!(reg364[(3'h5):(3'h4)] || (!reg119)))));
          for (forvar473 = (1'h0); (forvar473 < (2'h2)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 = ($unsigned($unsigned((~|(reg451 ^~ reg223)))) != (!{reg352,
                  wire383}));
            end
          reg475 = (-$unsigned((|$signed((^~reg352)))));
          for (forvar476 = (1'h0); (forvar476 < (3'h4)); forvar476 = (forvar476 + (1'h1)))
            begin
              reg477 = reg437;
              reg478 = reg359;
              reg479 <= reg460;
              reg480 = reg166[(3'h4):(1'h1)];
              reg481 <= $unsigned(reg453[(1'h1):(1'h0)]);
              reg482 <= ($signed($unsigned(($signed(reg353) > reg470))) ?
                  reg478[(4'h9):(3'h7)] : reg121);
              reg483 = {(!({(wire272 - reg371)} || $signed((reg137 ?
                      reg223 : wire272))))};
            end
          if ({{reg349[(4'h8):(3'h7)]}})
            begin
              reg484 = $unsigned((~^forvar473));
              reg485 = reg308;
              reg486 = $signed(($unsigned(((+reg478) ^ $unsigned(reg395))) >> ((|reg203) ?
                  reg325[(2'h2):(1'h1)] : reg461)));
              reg487 = $signed(reg354[(3'h4):(1'h0)]);
              reg488 = {(~reg482), $unsigned($signed(reg277[(3'h7):(3'h5)]))};
              reg489 = $unsigned((+{reg408,
                  (reg447 <<< $signed((7'h53))),
                  {$unsigned(reg454)}}));
            end
          else
            begin
              reg490 <= $signed(reg453[(2'h2):(1'h1)]);
              reg491 <= reg191[(3'h4):(3'h4)];
              reg492 = $unsigned(reg375);
              reg493 = $signed({(reg203 ? (-$signed(reg160)) : (8'hb4))});
              reg494 = ((8'ha0) <<< (&{(!{reg452, reg341})}));
            end
          for (forvar495 = (1'h0); (forvar495 < (1'h0)); forvar495 = (forvar495 + (1'h1)))
            begin
              reg496 <= $unsigned($unsigned(reg445));
              reg497 = $signed(reg165[(5'h11):(4'hd)]);
              reg498 <= (^reg323);
              reg499 = reg343[(5'h1b):(5'h14)];
              reg500 <= $signed($signed(($signed((reg466 || reg368)) ?
                  reg220[(3'h6):(2'h3)] : reg169)));
              reg501 <= reg371;
            end
        end
      if ($unsigned((7'h54)))
        begin
          if (((reg160[(5'h10):(4'he)] ?
              ($unsigned(reg239) != {$unsigned(reg354)}) : $unsigned($unsigned((reg467 ?
                  reg167 : reg458)))) == ((reg127[(3'h4):(1'h1)] ?
                  (~|$signed(wire94)) : reg289[(2'h3):(1'h1)]) ?
              (8'hb4) : (8'haa))))
            begin
              reg502 = $signed((~^reg496));
              reg503 <= $signed($unsigned((8'h9f)));
            end
          else
            begin
              reg503 <= reg181[(4'hf):(4'h8)];
              reg504 <= $signed(($signed(reg448[(1'h1):(1'h1)]) ?
                  ((reg295[(4'hf):(3'h5)] >>> (reg410 ? (8'hab) : (8'had))) ?
                      (reg133 == (reg354 && reg323)) : reg441) : ($signed((-wire272)) ?
                      ((reg496 ? (8'hb3) : (7'h49)) ^~ (&(8'hbd))) : ({reg171,
                          reg138,
                          reg475} && {reg448, reg478}))));
              reg505 <= reg178[(5'h11):(4'h8)];
              reg506 <= $unsigned((($signed((|reg418)) ^~ ($signed(reg418) || (&reg497))) & reg148));
              reg507 <= (({reg121[(2'h3):(1'h0)],
                      {{reg220, (8'hb6), reg459}, $signed(reg349), (|reg283)},
                      ($signed(reg483) ?
                          $signed((8'hbc)) : reg413[(4'h9):(3'h4)])} ?
                  {((reg266 ? reg167 : reg482) + reg239[(4'h9):(1'h0)]),
                      (reg448[(4'hc):(4'ha)] ?
                          {reg193} : (reg451 ? reg502 : reg224)),
                      $unsigned((&reg112))} : ((|$signed(reg390)) <<< (~|(reg475 <<< reg260)))) <<< $signed($signed(reg230)));
            end
          reg508 <= reg262[(4'h8):(2'h3)];
          reg509 = ((((^~{reg381, reg335}) ^ $signed(reg165)) >>> (7'h53)) ?
              (reg185[(3'h5):(3'h5)] >= (8'hac)) : (($signed((-wire97)) || $signed((&reg426))) != $signed($signed($signed(reg374)))));
          reg510 <= $signed(reg174);
          reg511 = (({$signed((reg152 == reg447)),
                  (~$unsigned(reg502)),
                  (7'h52)} ^~ $unsigned((~reg349[(5'h16):(3'h4)]))) ?
              reg265[(4'hd):(2'h2)] : (8'had));
          for (forvar512 = (1'h0); (forvar512 < (3'h6)); forvar512 = (forvar512 + (1'h1)))
            begin
              reg513 = {((|((reg336 ~^ (8'ha8)) * reg131)) - (reg469 * {(^reg160),
                      reg453[(1'h0):(1'h0)]})),
                  $signed((($unsigned((7'h4d)) ? (|(8'hb8)) : (7'h47)) ?
                      {((8'hb9) + (7'h40))} : (-reg354)))};
            end
          for (forvar514 = (1'h0); (forvar514 < (2'h2)); forvar514 = (forvar514 + (1'h1)))
            begin
              reg515 = (8'hab);
            end
        end
      else
        begin
          reg503 <= $signed((&(reg223[(3'h7):(3'h7)] & $signed((reg477 ?
              wire93 : reg440)))));
          for (forvar504 = (1'h0); (forvar504 < (3'h6)); forvar504 = (forvar504 + (1'h1)))
            begin
              reg505 <= (~^(($unsigned($signed((8'ha7))) ? reg156 : reg390) ?
                  wire272[(2'h2):(1'h0)] : $signed($signed((reg283 ?
                      (8'ha6) : reg411)))));
              reg506 <= ((&(7'h50)) ^ reg220);
              reg507 <= (-reg478);
              reg508 <= {(~^(^~(+reg229))),
                  ((|reg451[(3'h4):(2'h2)]) - $unsigned($signed(reg212[(3'h4):(2'h2)])))};
              reg510 <= (~|$unsigned((8'hba)));
            end
          for (forvar511 = (1'h0); (forvar511 < (3'h5)); forvar511 = (forvar511 + (1'h1)))
            begin
              reg512 <= ($unsigned(reg320[(3'h5):(2'h2)]) ?
                  (^~$signed(reg419[(1'h0):(1'h0)])) : $unsigned(reg434));
            end
          for (forvar513 = (1'h0); (forvar513 < (3'h5)); forvar513 = (forvar513 + (1'h1)))
            begin
              reg514 <= wire435;
            end
          for (forvar515 = (1'h0); (forvar515 < (2'h2)); forvar515 = (forvar515 + (1'h1)))
            begin
              reg516 = reg145;
            end
          if (reg491[(1'h1):(1'h0)])
            begin
              reg517 <= (reg512[(4'hb):(2'h2)] ?
                  reg456[(5'h12):(5'h12)] : (reg185 ?
                      {{$unsigned(reg467),
                              (reg483 >>> reg395),
                              (reg470 ? reg494 : reg145)},
                          reg469} : (&(reg444[(3'h7):(3'h5)] ?
                          reg368 : reg353[(4'h9):(2'h2)]))));
            end
          else
            begin
              reg517 <= ((reg470 ?
                  reg484[(3'h5):(3'h5)] : (((reg335 ? reg160 : (8'ha1)) ?
                          (reg458 ? reg145 : reg354) : (~|reg239)) ?
                      (^~$signed(reg309)) : reg492)) >= $unsigned((((reg133 | reg440) ?
                  $unsigned((7'h44)) : (^reg210)) || (-{wire95,
                  reg486,
                  reg507}))));
              reg518 <= reg121[(3'h5):(2'h3)];
              reg519 <= $unsigned($unsigned(reg357));
              reg520 <= $signed(($signed(reg469) > (reg469[(3'h4):(1'h0)] ?
                  ((-(7'h57)) >= $signed(reg366)) : forvar512[(1'h1):(1'h0)])));
              reg521 <= (~&{reg447});
            end
        end
      reg522 <= (forvar471 ? forvar473[(3'h7):(1'h0)] : $unsigned(reg434));
    end
  assign wire523 = $unsigned($unsigned(reg344));
  always
    @(posedge clk) begin
      reg524 <= reg189;
      reg525 <= $unsigned(((!reg147) ? reg263 : reg160[(5'h15):(5'h15)]));
      reg526 = $unsigned($unsigned((~^$signed(reg172))));
      reg527 <= reg500;
      for (forvar528 = (1'h0); (forvar528 < (3'h4)); forvar528 = (forvar528 + (1'h1)))
        begin
          if ($signed(reg482[(1'h0):(1'h0)]))
            begin
              reg529 <= reg347;
              reg530 <= (+(|(&reg526[(1'h0):(1'h0)])));
              reg531 = (^~$signed(($unsigned((reg437 ?
                  reg481 : reg290)) != {(reg248 ? (8'ha7) : reg224),
                  reg518[(5'h14):(3'h7)]})));
              reg532 = (~(7'h4e));
              reg533 = $signed((~^(reg532 << reg167)));
            end
          else
            begin
              reg531 = $unsigned({reg529[(2'h2):(1'h1)],
                  reg295[(4'he):(3'h6)]});
              reg532 = $signed((reg456 ?
                  (reg161 ?
                      {$unsigned(reg460)} : {wire382,
                          (reg407 ~^ (7'h45)),
                          (reg532 ? reg164 : reg313)}) : reg366));
              reg533 = (!$signed($signed(reg343[(1'h1):(1'h0)])));
              reg534 = reg265;
              reg535 <= reg104[(4'he):(2'h3)];
              reg536 = reg214[(4'hf):(2'h3)];
            end
          reg537 = ({(~&({reg224, (8'hbe), reg178} ?
                  reg320 : (|reg219)))} >> reg440[(5'h10):(4'hf)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar538 = (1'h0); (forvar538 < (3'h4)); forvar538 = (forvar538 + (1'h1)))
        begin
          reg539 <= reg334;
          reg540 <= (reg263[(2'h3):(2'h2)] & reg360[(4'hd):(2'h3)]);
          for (forvar541 = (1'h0); (forvar541 < (3'h6)); forvar541 = (forvar541 + (1'h1)))
            begin
              reg542 <= (-(!(^reg439)));
              reg543 <= reg344;
              reg544 <= reg277[(3'h7):(3'h6)];
              reg545 = {($signed(($signed(reg201) ?
                      {reg452, wire95} : (reg437 <= reg479))) + (8'hae))};
              reg546 = ($unsigned((|((wire273 ? (8'h9d) : (7'h50)) + ((7'h4c) ?
                      (7'h51) : reg500)))) ?
                  ({($signed(wire382) ?
                          (^(7'h44)) : wire435[(5'h1b):(5'h17)])} < ((reg236[(3'h7):(3'h6)] - ((7'h40) ?
                          reg545 : reg374)) ?
                      {((8'ha1) & reg353),
                          (~reg403),
                          (wire95 ? reg307 : reg119)} : (((8'ha2) ?
                          reg358 : reg395) + $unsigned(reg417)))) : (8'hb8));
            end
          for (forvar547 = (1'h0); (forvar547 < (3'h4)); forvar547 = (forvar547 + (1'h1)))
            begin
              reg548 = reg167[(1'h0):(1'h0)];
            end
          for (forvar549 = (1'h0); (forvar549 < (1'h0)); forvar549 = (forvar549 + (1'h1)))
            begin
              reg550 <= $signed($signed(reg178));
              reg551 <= ({$signed(((reg543 == reg465) ? (8'ha9) : (|reg390))),
                      $signed(((reg236 || reg481) != $signed(reg248))),
                      $unsigned((reg122 ? (&reg428) : ((8'hb1) >> reg379)))} ?
                  $unsigned({$signed(reg419),
                      $signed(reg548[(3'h5):(2'h2)]),
                      ((reg220 && reg481) ?
                          (reg142 ?
                              (8'ha1) : reg156) : $unsigned(reg147))}) : (8'ha8));
              reg552 <= (~|$signed((8'hb7)));
            end
          if ((reg552 ?
              wire97 : $signed((((reg105 <<< (7'h45)) >>> ((8'hbf) ?
                  reg305 : reg224)) == $unsigned(reg329)))))
            begin
              reg553 <= {reg352,
                  (+reg359[(1'h0):(1'h0)]),
                  reg241[(4'ha):(4'ha)]};
              reg554 = ($signed(reg336[(5'h13):(3'h4)]) && ($unsigned($unsigned((+reg374))) >>> $unsigned($signed(reg122))));
              reg555 <= $signed($signed({{$signed((7'h50)), reg518, {reg289}},
                  reg505[(2'h3):(1'h1)]}));
            end
          else
            begin
              reg553 <= ($signed(reg434[(3'h7):(1'h1)]) <= $signed($signed(reg535)));
              reg555 <= reg368;
              reg556 = $unsigned($signed((((~reg343) ?
                      reg290[(1'h1):(1'h1)] : ((7'h40) ? reg466 : reg344)) ?
                  {(^~reg408),
                      reg381[(1'h0):(1'h0)],
                      (~^reg334)} : (~^(reg313 ^ reg262)))));
              reg557 <= (-($signed((-reg290[(1'h0):(1'h0)])) ?
                  $unsigned((8'haa)) : reg141));
              reg558 <= ($signed($signed(reg496)) ?
                  $unsigned((^($unsigned(reg325) + ((8'hbc) ?
                      wire523 : (8'hb6))))) : ({(-$unsigned(reg98)),
                          $signed(reg314[(4'hb):(3'h6)]),
                          $unsigned($unsigned(reg445))} ?
                      $signed(((reg388 == reg503) ?
                          (reg192 ?
                              (7'h4b) : reg113) : $signed((8'hac)))) : reg212));
              reg559 = $unsigned((~^$unsigned($unsigned(reg552[(4'hb):(4'ha)]))));
              reg560 = $signed($unsigned((((+(8'h9c)) + (~|reg165)) < $unsigned($signed(reg111)))));
            end
        end
    end
  module561 #() modinst1366 (.wire563(reg189), .wire564(reg432), .clk(clk), .wire565(reg122), .y(wire1365), .wire562(reg250));
  assign wire1367 = $signed((reg123[(4'hd):(1'h1)] != reg362));
  always
    @(posedge clk) begin
      for (forvar1368 = (1'h0); (forvar1368 < (2'h3)); forvar1368 = (forvar1368 + (1'h1)))
        begin
          for (forvar1369 = (1'h0); (forvar1369 < (3'h5)); forvar1369 = (forvar1369 + (1'h1)))
            begin
              reg1370 <= (~^{(^(!{reg437}))});
              reg1371 <= $signed(($unsigned((^~reg408)) ^ $unsigned(($signed(reg164) || (reg185 ?
                  reg193 : reg104)))));
              reg1372 = (~|(reg407[(3'h4):(2'h2)] ?
                  (&(!reg426[(2'h3):(2'h3)])) : (reg505 ?
                      reg128 : (&(reg519 ~^ forvar1368)))));
              reg1373 = reg448[(5'h14):(4'hd)];
              reg1374 <= reg161[(5'h13):(5'h12)];
              reg1375 <= reg417[(5'h11):(4'hb)];
            end
          for (forvar1376 = (1'h0); (forvar1376 < (3'h5)); forvar1376 = (forvar1376 + (1'h1)))
            begin
              reg1377 <= ({(((7'h46) >> reg510[(5'h19):(4'ha)]) & reg490),
                      $unsigned(reg300[(4'h9):(1'h0)]),
                      reg504} ?
                  (~reg439) : reg456[(4'hc):(4'h9)]);
              reg1378 <= ((reg207[(5'h14):(2'h2)] ?
                      ($unsigned((reg113 + (8'hb3))) ?
                          $unsigned((reg530 ?
                              reg448 : reg417)) : reg132[(4'h8):(3'h4)]) : ($unsigned((wire435 ^~ wire273)) ^ (!$unsigned(reg293)))) ?
                  $signed((^reg192)) : $unsigned(reg391));
              reg1379 <= {(~((8'ha9) ?
                      (reg262[(1'h1):(1'h0)] <<< $signed((7'h52))) : reg152[(1'h0):(1'h0)]))};
            end
          for (forvar1380 = (1'h0); (forvar1380 < (1'h0)); forvar1380 = (forvar1380 + (1'h1)))
            begin
              reg1381 <= $signed($unsigned((-reg557[(4'hf):(1'h1)])));
              reg1382 <= reg207;
              reg1383 = reg522;
              reg1384 = $unsigned($signed((8'hbf)));
              reg1385 <= reg241[(2'h3):(2'h2)];
              reg1386 <= {(reg265 * (^~$unsigned(reg508[(5'h15):(5'h14)]))),
                  {reg317}};
            end
          reg1387 = $signed($signed((&$unsigned((reg527 ? reg1372 : reg104)))));
          reg1388 <= reg1372;
          reg1389 = {reg152[(3'h7):(1'h0)],
              ({((^reg138) * (reg243 ? reg352 : (7'h56))),
                  reg165,
                  (-$unsigned(reg320))} && $unsigned(reg115)),
              ($unsigned((8'hab)) - ($unsigned((reg336 ?
                  reg116 : reg467)) * {$signed(reg335), (~&reg542)}))};
        end
      for (forvar1390 = (1'h0); (forvar1390 < (1'h1)); forvar1390 = (forvar1390 + (1'h1)))
        begin
          reg1391 <= (reg366[(5'h12):(4'he)] ?
              $signed(((&(&reg535)) ^ reg292)) : reg268[(2'h3):(1'h1)]);
          if ((7'h51))
            begin
              reg1392 = $signed(((((reg230 ? reg224 : reg542) ?
                      {reg1379} : (^reg123)) - $unsigned(reg364)) ?
                  $unsigned(reg340[(1'h0):(1'h0)]) : $unsigned($unsigned(reg443))));
              reg1393 <= (8'hac);
              reg1394 = $unsigned((8'ha4));
              reg1395 <= ((((reg1386 ? reg371 : $unsigned((8'hae))) ?
                  {{(8'haa)}} : ($signed(reg325) && $unsigned(reg359))) >> (^$unsigned((~^reg524)))) & (|reg1378[(2'h2):(2'h2)]));
            end
          else
            begin
              reg1393 <= ((reg520[(4'hb):(4'ha)] ?
                      reg347 : ((7'h51) != (reg150 - reg411[(2'h2):(1'h0)]))) ?
                  (~^reg1378) : reg239[(3'h7):(3'h7)]);
              reg1394 = (^~(~|reg373[(4'ha):(2'h3)]));
              reg1395 <= ($unsigned(((!(reg535 > reg145)) <= {$signed(reg461)})) ?
                  $unsigned(reg347) : reg193[(3'h6):(3'h6)]);
              reg1396 = (reg123[(2'h2):(1'h1)] >= (^$unsigned((!{(8'h9e),
                  reg334}))));
              reg1397 <= (&((($signed(reg137) ?
                      ((8'ha6) > (7'h51)) : (reg340 ? reg310 : reg496)) ?
                  ((reg374 ? reg454 : reg260) + {reg504}) : ((~reg207) ?
                      (^~reg517) : (^reg465))) << $unsigned(reg395[(2'h3):(1'h1)])));
              reg1398 <= ((reg434 <<< $unsigned($unsigned($signed(reg525)))) || {(~&(reg1387 ?
                      $unsigned(reg1391) : (reg266 | reg142))),
                  (~|$unsigned($signed(reg552)))});
              reg1399 = ((($signed($unsigned(reg491)) ?
                      $signed(reg461) : (&(reg1382 ?
                          reg368 : reg388))) << (reg1375 ?
                      (((8'hbb) ? reg461 : reg359) ?
                          {reg230, (7'h4b), reg248} : {reg135,
                              reg557,
                              wire435}) : $signed((~|reg343)))) ?
                  ($unsigned((^$unsigned(forvar1376))) ?
                      $signed($signed(reg1395)) : reg286[(4'hd):(4'hd)]) : $signed(reg193[(4'hd):(4'hb)]));
            end
          if ({$unsigned($signed((|$signed(reg196))))})
            begin
              reg1400 = (~(|(^$signed((reg1385 != reg159)))));
              reg1401 <= ($unsigned($unsigned(reg344)) ?
                  (!((reg521[(2'h2):(1'h0)] == $unsigned(reg407)) + reg159)) : $unsigned($signed((+(|reg1377)))));
              reg1402 = $unsigned(((((reg196 ? reg510 : reg145) | {(8'hb2)}) ?
                  ($signed(reg171) != reg167[(1'h1):(1'h1)]) : {(reg368 >= reg555),
                      $unsigned(reg498),
                      {(8'hbb)}}) >>> (-reg201)));
              reg1403 <= ((|$unsigned($signed(((8'h9d) | (8'haf))))) ?
                  $signed($unsigned($signed((reg357 & reg116)))) : {(&(reg98[(4'ha):(1'h0)] ?
                          (wire97 ? reg296 : reg342) : wire435))});
              reg1404 = (($unsigned(((&(8'hb0)) ?
                      {reg270, reg342} : (&reg230))) ?
                  (reg510 + forvar1380[(1'h1):(1'h0)]) : {$unsigned(reg366[(5'h14):(3'h6)]),
                      ($signed(reg238) <<< $unsigned(reg116)),
                      $signed($signed(reg105))}) >= $signed($unsigned(($signed(reg445) ?
                  reg222 : {reg467}))));
            end
          else
            begin
              reg1400 = $signed($signed((~reg550[(2'h3):(1'h0)])));
              reg1401 <= (-$unsigned((~&$unsigned($unsigned((7'h4b))))));
              reg1402 = (8'ha4);
              reg1403 <= $signed($signed(reg450[(3'h5):(3'h5)]));
            end
          reg1405 = ((reg286[(4'h9):(1'h1)] ?
                  forvar1369 : ($signed($signed(reg357)) >>> (~^((8'hab) & (8'haa))))) ?
              (^(!(reg370 ?
                  (reg296 ?
                      reg529 : reg453) : reg192[(3'h5):(2'h3)]))) : (~|(reg524[(3'h4):(2'h3)] < wire1367)));
          for (forvar1406 = (1'h0); (forvar1406 < (3'h6)); forvar1406 = (forvar1406 + (1'h1)))
            begin
              reg1407 <= (8'hae);
              reg1408 = $unsigned(reg1396);
              reg1409 <= ((((&(reg357 ? reg1395 : reg133)) ?
                      (&(reg270 ? reg329 : (7'h48))) : (reg498 ?
                          (wire96 ? wire97 : reg127) : $unsigned((7'h51)))) ?
                  ({$signed(reg542), (~^reg1374)} ?
                      ((|reg504) < (reg524 ?
                          reg521 : reg329)) : reg440[(2'h2):(1'h1)]) : {reg105,
                      $signed({reg112}),
                      reg1399}) ^~ reg1385);
              reg1410 = $unsigned($unsigned((($unsigned(reg1386) >> reg434) * $signed($unsigned(reg132)))));
              reg1411 <= (!{(reg151[(3'h7):(2'h2)] == ((reg215 ~^ reg467) ?
                      (^~reg379) : reg142)),
                  {(!wire1367[(3'h4):(1'h1)]), reg428[(2'h3):(2'h2)]},
                  $unsigned((7'h58))});
              reg1412 <= ({reg373,
                  reg357[(4'hb):(4'h8)],
                  reg507[(3'h6):(3'h4)]} <= (reg450 < ((8'hae) ?
                  reg450[(3'h4):(3'h4)] : ($unsigned(reg390) ?
                      $unsigned(reg503) : reg308[(1'h0):(1'h0)]))));
            end
          for (forvar1413 = (1'h0); (forvar1413 < (3'h6)); forvar1413 = (forvar1413 + (1'h1)))
            begin
              reg1414 <= reg236[(4'he):(3'h5)];
              reg1415 = (!(({reg210, reg342[(3'h7):(1'h0)]} ?
                      $unsigned((reg229 >>> reg243)) : (!reg506[(4'h9):(3'h6)])) ?
                  reg219[(4'hc):(4'ha)] : $signed(((reg135 ? reg1384 : reg443) ?
                      (reg236 ? reg552 : reg1393) : reg379[(3'h7):(1'h0)]))));
            end
          if (reg456)
            begin
              reg1416 = reg432[(5'h19):(2'h2)];
              reg1417 = {reg467[(2'h2):(1'h0)],
                  ((($signed(reg1414) >>> (~&(7'h55))) ?
                          (reg542[(3'h5):(2'h3)] ?
                              $signed((8'ha3)) : $signed(reg1394)) : ((|forvar1390) >>> $signed((8'hb7)))) ?
                      reg551[(5'h17):(5'h13)] : $signed((-reg351[(2'h2):(1'h0)]))),
                  $unsigned(($signed($signed(reg1377)) ?
                      forvar1368 : $signed(reg535)))};
            end
          else
            begin
              reg1418 <= $signed((&reg1395[(3'h5):(3'h5)]));
              reg1419 <= (|((7'h4b) >>> (~$unsigned($signed(reg290)))));
              reg1420 = reg210[(2'h2):(2'h2)];
              reg1421 = ((7'h51) ~^ {reg165[(5'h14):(5'h10)]});
              reg1422 = (reg174 ?
                  ({((~|reg550) >> reg248[(5'h12):(4'ha)]),
                          ((reg173 >> reg453) ?
                              reg1407 : (reg179 ? reg1408 : reg434)),
                          {$unsigned(reg238), $unsigned(reg263)}} ?
                      $signed(reg461[(3'h6):(3'h6)]) : $unsigned(reg246[(4'hc):(2'h2)])) : reg135);
              reg1423 = reg368;
            end
        end
      reg1424 <= (|$unsigned((^(7'h54))));
    end
  assign wire1425 = {(-((~&(reg229 ?
                            reg164 : reg467)) < reg116[(3'h7):(2'h2)])),
                        reg150,
                        {$unsigned((+reg362[(4'hd):(4'hc)])),
                            $unsigned(($unsigned(reg131) || (~^(8'ha0))))}};
  always
    @(posedge clk) begin
      reg1426 = wire435[(3'h5):(2'h3)];
      for (forvar1427 = (1'h0); (forvar1427 < (2'h2)); forvar1427 = (forvar1427 + (1'h1)))
        begin
          reg1428 <= (reg360 ?
              $unsigned($signed(reg1397[(5'h18):(1'h1)])) : ($signed(reg137) ?
                  (7'h46) : $unsigned((^(reg257 ? (7'h4a) : reg463)))));
          reg1429 = ((reg520 ? (7'h49) : $unsigned(reg496[(5'h11):(3'h4)])) ?
              ((reg1378[(4'ha):(4'ha)] | {$signed((7'h4b)),
                  (~reg1370)}) << $signed($unsigned(reg426[(1'h0):(1'h0)]))) : reg491[(2'h3):(2'h3)]);
          reg1430 <= reg310[(3'h5):(3'h5)];
          reg1431 <= (-(^$unsigned(({reg289, reg257, reg467} ?
              (reg105 ? (7'h48) : reg1409) : reg542[(1'h0):(1'h0)]))));
          if ($unsigned(reg1393[(1'h1):(1'h0)]))
            begin
              reg1432 = ($unsigned((~|$signed($unsigned(reg262)))) == reg308);
            end
          else
            begin
              reg1432 = $signed(reg104[(2'h3):(1'h0)]);
              reg1433 <= $signed($unsigned(($signed((~|reg1401)) < reg270)));
              reg1434 <= (8'hb1);
              reg1435 <= wire1425[(4'h8):(1'h1)];
            end
          for (forvar1436 = (1'h0); (forvar1436 < (1'h1)); forvar1436 = (forvar1436 + (1'h1)))
            begin
              reg1437 <= (~(($signed($unsigned(reg239)) ?
                  ($signed(reg391) ?
                      (reg522 || reg181) : reg450[(3'h5):(1'h1)]) : ((reg374 ?
                          (7'h48) : wire96) ?
                      {(8'haa),
                          reg434,
                          (7'h48)} : $unsigned(reg500))) * reg153));
              reg1438 = ({$signed((&$unsigned(reg340))),
                  $signed(($unsigned(reg160) + (8'h9e)))} || ((^(reg169[(4'ha):(2'h3)] ?
                      (reg428 ^ reg467) : wire1425[(5'h1c):(4'ha)])) ?
                  $unsigned({$unsigned(reg128),
                      {reg347, reg390},
                      wire94}) : reg145[(2'h3):(2'h2)]));
              reg1439 <= (^~$signed((!$unsigned({(8'ha4), reg207, (8'hb0)}))));
              reg1440 = (reg116 >> $signed((($unsigned(reg337) <<< $unsigned(reg296)) >= ({reg454,
                      reg207,
                      reg104} ?
                  (^~reg1433) : $unsigned(reg215)))));
            end
        end
      reg1441 <= $signed((7'h45));
      reg1442 = (reg381[(1'h1):(1'h1)] ?
          {reg159[(3'h5):(2'h3)]} : reg481[(4'h9):(1'h0)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module561
#(parameter param1362 = {((~|(~^((8'ha6) ? (7'h44) : (8'hb5)))) ? (({(8'ha6)} ? (^(7'h57)) : ((7'h4b) >>> (8'h9f))) ? (~^{(7'h45)}) : (^((8'hbd) || (7'h55)))) : ((((8'hba) ? (8'h9d) : (8'ha7)) ? (7'h4c) : ((8'hb3) ? (7'h40) : (8'hbe))) > (8'hb1))), ((|{(-(8'ha2)), ((7'h46) * (8'hb6))}) ? {{((8'hb5) ? (7'h58) : (8'ha6)), ((7'h4d) | (7'h4e))}} : ((~|{(7'h58)}) == (((8'ha9) ? (8'hb6) : (7'h53)) ? ((8'ha7) ? (7'h4c) : (7'h4b)) : ((8'h9e) >>> (7'h55))))), (8'hbe)}, 
parameter param1363 = (!(param1362 ? {((param1362 ? param1362 : param1362) ^~ {param1362, (8'ha3), param1362}), ((param1362 ? param1362 : (7'h56)) ^~ (~&(8'h9e))), ({param1362, param1362} ? param1362 : param1362)} : (((+param1362) << ((7'h44) & param1362)) ? param1362 : (8'hab)))), 
parameter param1364 = param1363)
(y, clk, wire565, wire564, wire563, wire562);
  output wire [(32'h1cef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire565;
  input wire signed [(5'h19):(1'h0)] wire564;
  input wire signed [(2'h2):(1'h0)] wire563;
  input wire signed [(3'h6):(1'h0)] wire562;
  wire signed [(5'h1a):(1'h0)] wire1361;
  wire signed [(5'h12):(1'h0)] wire1359;
  wire signed [(2'h2):(1'h0)] wire1358;
  wire signed [(5'h19):(1'h0)] wire1357;
  wire signed [(2'h2):(1'h0)] wire1270;
  wire [(5'h1d):(1'h0)] wire1221;
  wire [(5'h12):(1'h0)] wire1220;
  wire signed [(4'h8):(1'h0)] wire1185;
  wire signed [(4'h9):(1'h0)] wire1110;
  wire signed [(5'h15):(1'h0)] wire1073;
  wire signed [(4'h9):(1'h0)] wire1072;
  wire [(5'h10):(1'h0)] wire1071;
  wire signed [(5'h1d):(1'h0)] wire1070;
  wire signed [(5'h15):(1'h0)] wire1068;
  wire signed [(5'h15):(1'h0)] wire615;
  wire signed [(5'h1e):(1'h0)] wire605;
  wire [(5'h13):(1'h0)] wire604;
  reg [(4'hf):(1'h0)] reg1356 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1355 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1353 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1352 = (1'h0);
  reg [(5'h11):(1'h0)] reg1351 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1347 = (1'h0);
  reg [(4'h8):(1'h0)] reg1345 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1343 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1342 = (1'h0);
  reg [(3'h7):(1'h0)] reg1340 = (1'h0);
  reg [(5'h10):(1'h0)] reg1339 = (1'h0);
  reg [(4'he):(1'h0)] reg1338 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1337 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1335 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1333 = (1'h0);
  reg [(4'hc):(1'h0)] reg1332 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1328 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1326 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1324 = (1'h0);
  reg [(3'h7):(1'h0)] reg1322 = (1'h0);
  reg [(5'h12):(1'h0)] reg1319 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1315 = (1'h0);
  reg [(5'h15):(1'h0)] reg1314 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1310 = (1'h0);
  reg [(4'h9):(1'h0)] reg1309 = (1'h0);
  reg [(4'h8):(1'h0)] reg1306 = (1'h0);
  reg [(4'hd):(1'h0)] reg1301 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1300 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1298 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1292 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1289 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1287 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1284 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1283 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1282 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1280 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1279 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1275 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1274 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1272 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1269 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1268 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1263 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1262 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1260 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1256 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1255 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1253 = (1'h0);
  reg [(5'h17):(1'h0)] reg1252 = (1'h0);
  reg [(5'h12):(1'h0)] reg1249 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1248 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1247 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1245 = (1'h0);
  reg [(5'h18):(1'h0)] reg1244 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1240 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1238 = (1'h0);
  reg [(2'h2):(1'h0)] reg1234 = (1'h0);
  reg [(2'h3):(1'h0)] reg1233 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1232 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1229 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1228 = (1'h0);
  reg [(5'h16):(1'h0)] reg1227 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1226 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1224 = (1'h0);
  reg [(5'h10):(1'h0)] reg1219 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1218 = (1'h0);
  reg [(4'he):(1'h0)] reg1217 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1216 = (1'h0);
  reg [(4'he):(1'h0)] reg1213 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1210 = (1'h0);
  reg [(3'h5):(1'h0)] reg1209 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1206 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1201 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1200 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1199 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1194 = (1'h0);
  reg [(5'h15):(1'h0)] reg1191 = (1'h0);
  reg [(5'h14):(1'h0)] reg1188 = (1'h0);
  reg [(5'h11):(1'h0)] reg1186 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1182 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1181 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1175 = (1'h0);
  reg [(4'hd):(1'h0)] reg1173 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1171 = (1'h0);
  reg [(5'h12):(1'h0)] reg1168 = (1'h0);
  reg [(5'h15):(1'h0)] reg1167 = (1'h0);
  reg [(5'h16):(1'h0)] reg1164 = (1'h0);
  reg [(5'h12):(1'h0)] reg1163 = (1'h0);
  reg [(4'ha):(1'h0)] reg1160 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1157 = (1'h0);
  reg [(4'hf):(1'h0)] reg1156 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1155 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1152 = (1'h0);
  reg [(4'ha):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1147 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1141 = (1'h0);
  reg [(3'h5):(1'h0)] reg1140 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1139 = (1'h0);
  reg [(5'h17):(1'h0)] reg1137 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1132 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1131 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1130 = (1'h0);
  reg [(5'h16):(1'h0)] reg1126 = (1'h0);
  reg [(5'h14):(1'h0)] reg1121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1118 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1113 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1108 = (1'h0);
  reg [(3'h5):(1'h0)] reg1106 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1105 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1104 = (1'h0);
  reg [(5'h13):(1'h0)] reg1102 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1100 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1098 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1097 = (1'h0);
  reg [(4'h8):(1'h0)] reg1095 = (1'h0);
  reg [(5'h14):(1'h0)] reg1094 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1093 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1092 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1090 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1089 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1086 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1083 = (1'h0);
  reg [(5'h16):(1'h0)] reg1081 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1077 = (1'h0);
  reg [(5'h11):(1'h0)] reg697 = (1'h0);
  reg [(4'hb):(1'h0)] reg696 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg695 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg693 = (1'h0);
  reg [(5'h10):(1'h0)] reg692 = (1'h0);
  reg [(4'hc):(1'h0)] reg691 = (1'h0);
  reg [(3'h6):(1'h0)] reg690 = (1'h0);
  reg [(5'h1f):(1'h0)] reg685 = (1'h0);
  reg [(4'h8):(1'h0)] reg674 = (1'h0);
  reg [(5'h18):(1'h0)] reg667 = (1'h0);
  reg [(4'h8):(1'h0)] reg680 = (1'h0);
  reg [(4'ha):(1'h0)] reg679 = (1'h0);
  reg [(5'h1a):(1'h0)] reg678 = (1'h0);
  reg [(5'h12):(1'h0)] reg677 = (1'h0);
  reg [(4'h8):(1'h0)] reg675 = (1'h0);
  reg [(3'h5):(1'h0)] reg670 = (1'h0);
  reg [(5'h1c):(1'h0)] reg669 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg663 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg658 = (1'h0);
  reg [(5'h11):(1'h0)] reg657 = (1'h0);
  reg [(4'he):(1'h0)] reg653 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg652 = (1'h0);
  reg [(3'h7):(1'h0)] reg650 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg649 = (1'h0);
  reg [(4'hc):(1'h0)] reg646 = (1'h0);
  reg [(5'h16):(1'h0)] reg630 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg644 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg643 = (1'h0);
  reg [(5'h1a):(1'h0)] reg642 = (1'h0);
  reg signed [(4'he):(1'h0)] reg641 = (1'h0);
  reg [(4'hf):(1'h0)] reg639 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg638 = (1'h0);
  reg signed [(4'he):(1'h0)] reg637 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg636 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg634 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg633 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg632 = (1'h0);
  reg [(3'h4):(1'h0)] reg631 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg625 = (1'h0);
  reg [(5'h10):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg621 = (1'h0);
  reg [(4'hd):(1'h0)] reg618 = (1'h0);
  reg [(5'h1a):(1'h0)] reg616 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg612 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg603 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg601 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg597 = (1'h0);
  reg [(4'hc):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg591 = (1'h0);
  reg [(5'h15):(1'h0)] reg590 = (1'h0);
  reg [(2'h2):(1'h0)] reg588 = (1'h0);
  reg [(4'hc):(1'h0)] reg582 = (1'h0);
  reg [(5'h1f):(1'h0)] reg581 = (1'h0);
  reg [(5'h18):(1'h0)] reg579 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg577 = (1'h0);
  reg [(5'h17):(1'h0)] reg576 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg573 = (1'h0);
  reg [(4'ha):(1'h0)] reg572 = (1'h0);
  reg [(2'h3):(1'h0)] reg571 = (1'h0);
  reg [(5'h1f):(1'h0)] reg570 = (1'h0);
  reg [(5'h19):(1'h0)] reg568 = (1'h0);
  reg [(5'h14):(1'h0)] reg567 = (1'h0);
  reg [(5'h15):(1'h0)] reg566 = (1'h0);
  reg [(5'h18):(1'h0)] reg1360 = (1'h0);
  reg [(4'hd):(1'h0)] reg1354 = (1'h0);
  reg [(5'h18):(1'h0)] reg1350 = (1'h0);
  reg [(4'ha):(1'h0)] reg1349 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar1348 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1346 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1344 = (1'h0);
  reg [(4'h8):(1'h0)] reg1341 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1336 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1334 = (1'h0);
  reg [(4'he):(1'h0)] reg1331 = (1'h0);
  reg [(5'h11):(1'h0)] reg1330 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1329 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1327 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1325 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1323 = (1'h0);
  reg [(3'h7):(1'h0)] reg1323 = (1'h0);
  reg [(5'h19):(1'h0)] reg1321 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1320 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar1311 = (1'h0);
  reg [(2'h3):(1'h0)] reg1318 = (1'h0);
  reg [(5'h17):(1'h0)] reg1317 = (1'h0);
  reg [(5'h13):(1'h0)] reg1316 = (1'h0);
  reg [(4'h9):(1'h0)] reg1313 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1312 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1311 = (1'h0);
  reg [(5'h13):(1'h0)] reg1308 = (1'h0);
  reg [(3'h6):(1'h0)] reg1307 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1305 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1304 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1303 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1302 = (1'h0);
  reg [(5'h17):(1'h0)] reg1299 = (1'h0);
  reg [(4'ha):(1'h0)] reg1297 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1296 = (1'h0);
  reg [(2'h3):(1'h0)] reg1295 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1294 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar1293 = (1'h0);
  reg [(4'h9):(1'h0)] reg1291 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1290 = (1'h0);
  reg [(5'h10):(1'h0)] reg1288 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1286 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1285 = (1'h0);
  reg [(4'h8):(1'h0)] reg1281 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1278 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1277 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1276 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1273 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1271 = (1'h0);
  reg [(2'h2):(1'h0)] reg1267 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1266 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1265 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1264 = (1'h0);
  reg [(4'he):(1'h0)] reg1261 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1250 = (1'h0);
  reg [(4'he):(1'h0)] reg1259 = (1'h0);
  reg [(2'h2):(1'h0)] reg1258 = (1'h0);
  reg [(5'h19):(1'h0)] reg1257 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1254 = (1'h0);
  reg [(5'h12):(1'h0)] reg1251 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1250 = (1'h0);
  reg [(4'hc):(1'h0)] reg1246 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1243 = (1'h0);
  reg [(4'hc):(1'h0)] reg1242 = (1'h0);
  reg [(5'h19):(1'h0)] reg1241 = (1'h0);
  reg [(5'h14):(1'h0)] reg1239 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1237 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1236 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1235 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1231 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1230 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1225 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1223 = (1'h0);
  reg [(5'h19):(1'h0)] reg1222 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1215 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1214 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1212 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1211 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1208 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1207 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1205 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1204 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1203 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1202 = (1'h0);
  reg [(5'h12):(1'h0)] reg1198 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1197 = (1'h0);
  reg [(5'h19):(1'h0)] reg1196 = (1'h0);
  reg [(2'h3):(1'h0)] reg1195 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1193 = (1'h0);
  reg [(4'h9):(1'h0)] reg1192 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1190 = (1'h0);
  reg [(5'h13):(1'h0)] reg1189 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1187 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1184 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1183 = (1'h0);
  reg [(5'h14):(1'h0)] reg1180 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1179 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1178 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1177 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1176 = (1'h0);
  reg [(5'h11):(1'h0)] reg1174 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1172 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1170 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1169 = (1'h0);
  reg [(5'h12):(1'h0)] reg1166 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1165 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1162 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1161 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1159 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1158 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1154 = (1'h0);
  reg [(4'he):(1'h0)] forvar1153 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1151 = (1'h0);
  reg [(5'h19):(1'h0)] reg1149 = (1'h0);
  reg [(5'h18):(1'h0)] reg1148 = (1'h0);
  reg [(4'he):(1'h0)] reg1146 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1145 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1144 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1143 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1142 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1139 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1133 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1129 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1138 = (1'h0);
  reg [(5'h13):(1'h0)] reg1136 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1135 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1134 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1133 = (1'h0);
  reg [(5'h12):(1'h0)] reg1129 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1128 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1127 = (1'h0);
  reg [(3'h4):(1'h0)] reg1125 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1124 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1123 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1122 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1120 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1119 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1117 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1116 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1115 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1114 = (1'h0);
  reg [(4'h8):(1'h0)] reg1112 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1111 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1109 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar1107 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1103 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1101 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar1099 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1091 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1096 = (1'h0);
  reg [(4'h8):(1'h0)] reg1091 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1085 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1088 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1087 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1085 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1082 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1074 = (1'h0);
  reg [(4'hb):(1'h0)] reg1080 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1079 = (1'h0);
  reg [(3'h4):(1'h0)] reg1078 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1076 = (1'h0);
  reg [(3'h7):(1'h0)] reg1075 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1074 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg701 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg700 = (1'h0);
  reg [(4'h9):(1'h0)] reg699 = (1'h0);
  reg [(2'h3):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg694 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg689 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg688 = (1'h0);
  reg [(5'h19):(1'h0)] reg687 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar684 = (1'h0);
  reg [(3'h4):(1'h0)] forvar683 = (1'h0);
  reg [(2'h3):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg682 = (1'h0);
  reg [(3'h4):(1'h0)] reg681 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg676 = (1'h0);
  reg [(5'h14):(1'h0)] forvar674 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg673 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg672 = (1'h0);
  reg [(5'h15):(1'h0)] reg671 = (1'h0);
  reg [(5'h16):(1'h0)] forvar667 = (1'h0);
  reg [(3'h7):(1'h0)] reg666 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar665 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg664 = (1'h0);
  reg [(4'h9):(1'h0)] reg662 = (1'h0);
  reg [(5'h1d):(1'h0)] reg661 = (1'h0);
  reg [(5'h13):(1'h0)] forvar660 = (1'h0);
  reg [(5'h13):(1'h0)] reg659 = (1'h0);
  reg [(5'h14):(1'h0)] reg656 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg655 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg654 = (1'h0);
  reg [(3'h6):(1'h0)] reg651 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar648 = (1'h0);
  reg [(4'hf):(1'h0)] forvar647 = (1'h0);
  reg [(5'h1b):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg640 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg635 = (1'h0);
  reg [(4'hd):(1'h0)] forvar630 = (1'h0);
  reg [(4'ha):(1'h0)] reg629 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg627 = (1'h0);
  reg [(2'h3):(1'h0)] reg626 = (1'h0);
  reg [(4'hb):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg622 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg620 = (1'h0);
  reg [(4'h9):(1'h0)] reg619 = (1'h0);
  reg [(4'he):(1'h0)] reg617 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg614 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg613 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg611 = (1'h0);
  reg [(5'h1c):(1'h0)] reg610 = (1'h0);
  reg signed [(4'he):(1'h0)] reg609 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar607 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg606 = (1'h0);
  reg [(5'h12):(1'h0)] reg602 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg599 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg598 = (1'h0);
  reg [(3'h5):(1'h0)] forvar596 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar594 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg593 = (1'h0);
  reg [(5'h13):(1'h0)] reg589 = (1'h0);
  reg [(4'hb):(1'h0)] reg587 = (1'h0);
  reg [(5'h15):(1'h0)] forvar586 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg585 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg584 = (1'h0);
  reg [(4'hb):(1'h0)] reg583 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar570 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg580 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg578 = (1'h0);
  reg [(5'h12):(1'h0)] reg575 = (1'h0);
  reg [(3'h7):(1'h0)] reg569 = (1'h0);
  assign y = {wire1361,
                 wire1359,
                 wire1358,
                 wire1357,
                 wire1270,
                 wire1221,
                 wire1220,
                 wire1185,
                 wire1110,
                 wire1073,
                 wire1072,
                 wire1071,
                 wire1070,
                 wire1068,
                 wire615,
                 wire605,
                 wire604,
                 reg1356,
                 reg1355,
                 reg1353,
                 reg1352,
                 reg1351,
                 reg1347,
                 reg1345,
                 reg1343,
                 reg1342,
                 reg1340,
                 reg1339,
                 reg1338,
                 reg1337,
                 reg1335,
                 reg1333,
                 reg1332,
                 reg1328,
                 reg1326,
                 reg1324,
                 reg1322,
                 reg1319,
                 reg1315,
                 reg1314,
                 reg1310,
                 reg1309,
                 reg1306,
                 reg1301,
                 reg1300,
                 reg1298,
                 reg1292,
                 reg1289,
                 reg1287,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1280,
                 reg1279,
                 reg1275,
                 reg1274,
                 reg1272,
                 reg1269,
                 reg1268,
                 reg1263,
                 reg1262,
                 reg1260,
                 reg1256,
                 reg1255,
                 reg1253,
                 reg1252,
                 reg1249,
                 reg1248,
                 reg1247,
                 reg1245,
                 reg1244,
                 reg1240,
                 reg1238,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1229,
                 reg1228,
                 reg1227,
                 reg1226,
                 reg1224,
                 reg1219,
                 reg1218,
                 reg1217,
                 reg1216,
                 reg1213,
                 reg1210,
                 reg1209,
                 reg1206,
                 reg1201,
                 reg1200,
                 reg1199,
                 reg1194,
                 reg1191,
                 reg1188,
                 reg1186,
                 reg1182,
                 reg1181,
                 reg1175,
                 reg1173,
                 reg1171,
                 reg1168,
                 reg1167,
                 reg1164,
                 reg1163,
                 reg1160,
                 reg1157,
                 reg1156,
                 reg1155,
                 reg1152,
                 reg1150,
                 reg1147,
                 reg1141,
                 reg1140,
                 reg1139,
                 reg1137,
                 reg1132,
                 reg1131,
                 reg1130,
                 reg1126,
                 reg1121,
                 reg1118,
                 reg1113,
                 reg1108,
                 reg1106,
                 reg1105,
                 reg1104,
                 reg1102,
                 reg1100,
                 reg1098,
                 reg1097,
                 reg1095,
                 reg1094,
                 reg1093,
                 reg1092,
                 reg1090,
                 reg1089,
                 reg1086,
                 reg1083,
                 reg1081,
                 reg1077,
                 reg697,
                 reg696,
                 reg695,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg685,
                 reg674,
                 reg667,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg675,
                 reg670,
                 reg669,
                 reg668,
                 reg663,
                 reg658,
                 reg657,
                 reg653,
                 reg652,
                 reg650,
                 reg649,
                 reg646,
                 reg630,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg628,
                 reg625,
                 reg623,
                 reg621,
                 reg618,
                 reg616,
                 reg612,
                 reg603,
                 reg601,
                 reg597,
                 reg595,
                 reg592,
                 reg591,
                 reg590,
                 reg588,
                 reg582,
                 reg581,
                 reg579,
                 reg577,
                 reg576,
                 reg574,
                 reg573,
                 reg572,
                 reg571,
                 reg570,
                 reg568,
                 reg567,
                 reg566,
                 reg1360,
                 reg1354,
                 reg1350,
                 reg1349,
                 forvar1348,
                 reg1346,
                 reg1344,
                 reg1341,
                 reg1336,
                 forvar1334,
                 reg1331,
                 reg1330,
                 reg1329,
                 reg1327,
                 reg1325,
                 forvar1323,
                 reg1323,
                 reg1321,
                 reg1320,
                 forvar1311,
                 reg1318,
                 reg1317,
                 reg1316,
                 reg1313,
                 reg1312,
                 reg1311,
                 reg1308,
                 reg1307,
                 reg1305,
                 reg1304,
                 reg1303,
                 reg1302,
                 reg1299,
                 reg1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 forvar1293,
                 reg1291,
                 reg1290,
                 reg1288,
                 reg1286,
                 forvar1285,
                 reg1281,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1273,
                 forvar1271,
                 reg1267,
                 reg1266,
                 reg1265,
                 reg1264,
                 reg1261,
                 reg1250,
                 reg1259,
                 reg1258,
                 reg1257,
                 reg1254,
                 reg1251,
                 forvar1250,
                 reg1246,
                 reg1243,
                 reg1242,
                 reg1241,
                 reg1239,
                 reg1237,
                 reg1236,
                 forvar1235,
                 reg1231,
                 forvar1230,
                 forvar1225,
                 forvar1223,
                 reg1222,
                 reg1215,
                 reg1214,
                 reg1212,
                 reg1211,
                 reg1208,
                 forvar1207,
                 forvar1205,
                 reg1204,
                 reg1203,
                 reg1202,
                 reg1198,
                 reg1197,
                 reg1196,
                 reg1195,
                 reg1193,
                 reg1192,
                 reg1190,
                 reg1189,
                 reg1187,
                 reg1184,
                 reg1183,
                 reg1180,
                 reg1179,
                 forvar1178,
                 reg1177,
                 reg1176,
                 reg1174,
                 reg1172,
                 reg1170,
                 reg1169,
                 reg1166,
                 reg1165,
                 forvar1162,
                 reg1161,
                 reg1159,
                 reg1158,
                 reg1154,
                 forvar1153,
                 reg1151,
                 reg1149,
                 reg1148,
                 reg1146,
                 reg1145,
                 forvar1144,
                 reg1143,
                 reg1142,
                 forvar1139,
                 reg1133,
                 forvar1129,
                 reg1138,
                 reg1136,
                 reg1135,
                 reg1134,
                 forvar1133,
                 reg1129,
                 reg1128,
                 reg1127,
                 reg1125,
                 reg1124,
                 reg1123,
                 forvar1122,
                 forvar1120,
                 reg1119,
                 reg1117,
                 reg1116,
                 forvar1115,
                 forvar1114,
                 reg1112,
                 reg1111,
                 reg1109,
                 forvar1107,
                 reg1103,
                 reg1101,
                 forvar1099,
                 forvar1091,
                 reg1096,
                 reg1091,
                 reg1085,
                 reg1088,
                 reg1087,
                 forvar1085,
                 reg1084,
                 forvar1082,
                 forvar1074,
                 reg1080,
                 reg1079,
                 reg1078,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg701,
                 reg700,
                 reg699,
                 reg698,
                 reg694,
                 reg689,
                 reg688,
                 reg687,
                 reg686,
                 forvar684,
                 forvar683,
                 reg665,
                 reg682,
                 reg681,
                 reg676,
                 forvar674,
                 reg673,
                 reg672,
                 reg671,
                 forvar667,
                 reg666,
                 forvar665,
                 reg664,
                 reg662,
                 reg661,
                 forvar660,
                 reg659,
                 reg656,
                 reg655,
                 reg654,
                 reg651,
                 forvar648,
                 forvar647,
                 reg645,
                 reg640,
                 reg635,
                 forvar630,
                 reg629,
                 reg627,
                 reg626,
                 reg624,
                 reg622,
                 reg620,
                 reg619,
                 reg617,
                 reg614,
                 reg613,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 forvar607,
                 reg606,
                 reg602,
                 reg600,
                 reg599,
                 reg598,
                 forvar596,
                 forvar594,
                 reg593,
                 reg589,
                 reg587,
                 forvar586,
                 reg585,
                 reg584,
                 reg583,
                 forvar570,
                 reg580,
                 reg578,
                 reg575,
                 reg569,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((&($unsigned((8'h9c)) && (~^(~(~&wire565))))))
        begin
          reg566 <= wire563;
          reg567 <= reg566[(4'h9):(1'h1)];
          if ((wire565 ?
              ($signed($signed(wire565)) | wire565[(3'h4):(1'h1)]) : {wire562[(1'h1):(1'h0)],
                  (({wire562} <= reg567) ?
                      ({wire563, reg566, wire563} && {reg566,
                          reg567}) : $unsigned((wire562 ? reg567 : wire562))),
                  (wire564 <= $signed((wire565 ? wire565 : wire565)))}))
            begin
              reg568 <= ((7'h58) ?
                  {(^$unsigned($unsigned(wire562)))} : $unsigned(wire563[(1'h0):(1'h0)]));
              reg569 = (^~(-reg566));
            end
          else
            begin
              reg569 = $signed(reg567);
              reg570 <= $signed((8'hb6));
              reg571 <= $signed(wire562[(2'h3):(1'h0)]);
              reg572 <= (&$signed((7'h46)));
              reg573 <= {((($unsigned(wire563) <<< wire565) ?
                          reg569[(1'h1):(1'h1)] : {$signed(reg570),
                              (reg569 & (8'haf)),
                              wire564[(1'h1):(1'h1)]}) ?
                      (~^($unsigned((7'h47)) ?
                          reg570[(3'h7):(1'h1)] : $unsigned(reg571))) : reg570)};
              reg574 <= (((($signed(reg573) ?
                      wire563[(1'h1):(1'h1)] : (reg566 ~^ reg572)) ^ (+(^~reg572))) >= $unsigned(({(8'ha8),
                      wire562} == (reg571 & reg572)))) ?
                  $unsigned(reg571[(2'h2):(1'h1)]) : (|((reg568[(5'h16):(4'h9)] ?
                          wire563[(2'h2):(2'h2)] : wire565[(3'h4):(1'h1)]) ?
                      $signed((7'h50)) : reg570[(5'h1e):(5'h12)])));
            end
          if (($unsigned((wire562 ?
              reg568 : reg573[(3'h5):(2'h2)])) > (({(reg567 >> reg567),
              (^~(8'ha9)),
              $signed(reg568)} <= reg573[(4'hf):(4'hb)]) < $signed($signed((~reg567))))))
            begin
              reg575 = ((($unsigned((reg567 ? wire563 : wire565)) ?
                          ((reg573 ? reg568 : reg568) << ((8'h9c) ?
                              wire563 : reg571)) : wire565) ?
                      {($unsigned(wire563) << $unsigned((8'hb9))),
                          ((wire565 ? reg566 : wire565) >> {reg571,
                              (8'hb5),
                              reg566}),
                          (7'h50)} : (~reg567[(5'h12):(4'ha)])) ?
                  (!reg570) : (^~$unsigned(wire563[(1'h0):(1'h0)])));
              reg576 <= $unsigned($unsigned($signed($signed($signed((8'h9d))))));
              reg577 <= reg571;
              reg578 = {wire563[(2'h2):(1'h1)],
                  reg568[(4'hd):(4'hc)],
                  reg568[(1'h0):(1'h0)]};
              reg579 <= (((($signed(wire565) || reg574[(3'h5):(3'h5)]) * {$signed(reg571),
                          (reg569 & reg567),
                          $signed(reg570)}) ?
                      $unsigned((-$unsigned((8'hbd)))) : $unsigned(reg568)) ?
                  $signed((reg569[(1'h0):(1'h0)] != ((wire564 ?
                      (7'h4c) : reg577) && reg569[(3'h6):(3'h6)]))) : {(($signed(reg567) >>> (~reg571)) >= (+((8'hb3) ?
                          reg574 : reg570)))});
            end
          else
            begin
              reg575 = $unsigned({$unsigned(($unsigned(reg566) & (&reg569)))});
              reg576 <= ($unsigned(reg569) ? wire565[(2'h3):(1'h0)] : reg571);
              reg578 = $unsigned((wire564 ~^ reg577));
              reg580 = $signed($unsigned(wire565));
              reg581 <= (~&((~&$signed($unsigned(reg567))) ?
                  $unsigned(($unsigned(reg578) < $signed(reg575))) : (^~{$signed((7'h57)),
                      reg579,
                      (reg575 ? (8'ha8) : wire564)})));
              reg582 <= $signed((^reg572));
            end
        end
      else
        begin
          reg569 = (!((((reg573 ? wire562 : (8'hb4)) ?
                  reg573[(5'h13):(2'h3)] : (~&reg573)) > $signed((8'ha3))) ?
              {wire562[(1'h0):(1'h0)],
                  ($signed(reg570) ?
                      $signed(reg579) : $signed(wire565))} : ((wire564 <= {reg576,
                      (7'h4d),
                      (8'hb7)}) ?
                  ((|reg569) << reg579) : reg580)));
          for (forvar570 = (1'h0); (forvar570 < (2'h3)); forvar570 = (forvar570 + (1'h1)))
            begin
              reg571 <= $signed(reg579[(1'h1):(1'h0)]);
              reg575 = ($signed(($unsigned(forvar570) ?
                  ($unsigned(reg582) ?
                      $signed(forvar570) : (reg567 ?
                          reg571 : reg568)) : ({reg577,
                      reg581,
                      reg575} && (8'ha9)))) <= reg578);
              reg578 = (^~((~reg575[(3'h4):(1'h1)]) ?
                  reg571[(1'h1):(1'h1)] : reg572));
              reg579 <= ($unsigned((!reg569[(1'h1):(1'h1)])) ?
                  $unsigned(reg566[(4'h9):(1'h1)]) : $unsigned({wire565[(1'h0):(1'h0)],
                      ((reg568 > reg574) ?
                          $unsigned((8'hb8)) : (reg570 ^ reg570))}));
              reg580 = {{(^~reg581), reg567},
                  $unsigned(wire562[(3'h5):(1'h0)])};
            end
          reg583 = $unsigned(((reg566[(5'h15):(3'h5)] ?
                  ((7'h4a) ?
                      ((7'h49) ?
                          reg575 : reg578) : (reg582 > reg575)) : $unsigned((reg574 ?
                      reg578 : reg575))) ?
              reg572 : (8'hbb)));
          reg584 = (reg578[(2'h2):(1'h1)] ?
              reg580[(4'hf):(1'h0)] : {$signed((~$unsigned(reg568)))});
          reg585 = $unsigned(reg583[(3'h5):(1'h0)]);
          for (forvar586 = (1'h0); (forvar586 < (2'h3)); forvar586 = (forvar586 + (1'h1)))
            begin
              reg587 = (7'h47);
              reg588 <= reg576[(4'hb):(3'h5)];
              reg589 = ((+(({reg581, reg584} >> $signed(reg588)) ?
                      ({forvar570} ~^ (forvar570 ?
                          reg581 : (7'h43))) : reg566[(4'hd):(4'hb)])) ?
                  reg581 : reg580[(4'hb):(1'h0)]);
              reg590 <= reg573;
              reg591 <= (^~reg589);
              reg592 <= ($unsigned($signed($unsigned((reg582 ?
                      wire562 : reg566)))) ?
                  reg580[(2'h3):(2'h2)] : {$signed((reg580[(4'hf):(3'h5)] ?
                          (wire563 ?
                              reg582 : (7'h41)) : (forvar570 << reg574))),
                      (-((reg582 ? reg587 : (7'h58)) ?
                          (reg566 ^ (7'h4f)) : $signed(wire565))),
                      $signed(reg579[(1'h1):(1'h0)])});
              reg593 = reg575;
            end
        end
      for (forvar594 = (1'h0); (forvar594 < (3'h6)); forvar594 = (forvar594 + (1'h1)))
        begin
          reg595 <= (7'h48);
          for (forvar596 = (1'h0); (forvar596 < (1'h0)); forvar596 = (forvar596 + (1'h1)))
            begin
              reg597 <= $unsigned((7'h58));
              reg598 = $signed(($unsigned((~&reg572)) ?
                  ((-{wire565, reg589, reg566}) ?
                      $signed((reg582 ?
                          reg567 : reg585)) : (~^(reg578 ^~ reg576))) : reg567));
              reg599 = reg588;
              reg600 = reg599;
              reg601 <= $unsigned(((!reg592[(1'h1):(1'h0)]) >>> (~reg583)));
              reg602 = (|(reg591[(5'h1b):(5'h15)] & reg591));
            end
          reg603 <= reg582[(2'h2):(1'h1)];
        end
    end
  assign wire604 = reg597[(4'h8):(3'h5)];
  assign wire605 = {reg572,
                       $signed(({{(7'h4c), reg571, wire564},
                           (|reg588)} >> (~reg595[(4'h8):(4'h8)]))),
                       $unsigned(reg573)};
  always
    @(posedge clk) begin
      reg606 = reg573[(5'h15):(4'ha)];
      for (forvar607 = (1'h0); (forvar607 < (2'h2)); forvar607 = (forvar607 + (1'h1)))
        begin
          if ((($signed(wire564) ?
                  {((reg574 >>> reg574) | $unsigned(wire562)),
                      {(forvar607 ? reg566 : reg572), (^reg579)}} : (8'hba)) ?
              ((((wire564 ?
                  (8'h9c) : reg590) ~^ $signed(wire562)) ^~ (~&((7'h53) ?
                  reg592 : reg597))) + $unsigned((&(&reg567)))) : reg572[(4'h9):(2'h3)]))
            begin
              reg608 = reg606;
              reg609 = reg590;
              reg610 = wire565[(2'h2):(1'h0)];
              reg611 = ($unsigned(reg579) << (~&(~|(~&$signed(reg576)))));
              reg612 <= (+(~^reg568));
              reg613 = reg609[(4'h9):(4'h9)];
              reg614 = $unsigned($signed($signed(($unsigned(reg613) * (reg606 ?
                  (8'hbc) : (7'h44))))));
            end
          else
            begin
              reg608 = {$unsigned(($unsigned((reg574 ? reg609 : reg568)) ?
                      {$unsigned(reg570)} : ((reg573 ?
                          reg603 : reg571) <= (reg591 ^~ (8'hbd)))))};
              reg609 = $unsigned(reg568[(4'hf):(4'hf)]);
              reg610 = reg613[(3'h5):(2'h2)];
            end
        end
    end
  assign wire615 = (-$unsigned(reg591));
  always
    @(posedge clk) begin
      reg616 <= reg582;
      reg617 = $unsigned(($signed((+reg597)) & (~^({(7'h45)} ?
          $signed((7'h4c)) : reg568))));
      if ($signed(((~$unsigned(wire565)) && (~|wire564))))
        begin
          if ($signed(reg573))
            begin
              reg618 <= reg570[(5'h10):(2'h2)];
              reg619 = reg616[(5'h10):(4'hc)];
              reg620 = (($unsigned((~|wire615[(4'hb):(3'h4)])) & wire604[(3'h7):(2'h3)]) << reg567);
            end
          else
            begin
              reg619 = (&{$signed(((~&reg570) == reg574)), reg595, (+reg591)});
              reg621 <= (-$unsigned(reg620));
            end
          if ((|reg592))
            begin
              reg622 = (wire562[(3'h5):(1'h1)] && ($unsigned(wire563[(1'h1):(1'h0)]) <<< (reg590[(4'hf):(1'h0)] << {reg568[(5'h19):(2'h2)],
                  $signed(reg612)})));
              reg623 <= (8'ha1);
              reg624 = ((reg588 | reg601) ?
                  (-$unsigned((wire562 < (reg620 >= reg617)))) : $signed(((reg619 >>> (7'h51)) ?
                      $unsigned($unsigned(wire565)) : (~|wire564))));
              reg625 <= (reg617 ?
                  reg574[(5'h10):(4'hf)] : ({reg582[(3'h4):(2'h3)],
                      {{reg623}, reg620, {reg620, reg603, reg603}},
                      reg603[(3'h6):(3'h5)]} || $unsigned($signed(reg570))));
              reg626 = reg582;
            end
          else
            begin
              reg622 = reg591;
              reg624 = (7'h57);
              reg625 <= $unsigned(reg623[(4'hd):(1'h1)]);
              reg626 = (reg626[(1'h0):(1'h0)] ?
                  ((~^(7'h40)) ?
                      reg591[(4'he):(4'h9)] : ($unsigned($unsigned(reg619)) ?
                          (reg577[(3'h6):(2'h3)] ?
                              $signed(reg603) : (reg579 ?
                                  reg612 : reg618)) : (((7'h4e) ?
                                  reg573 : reg579) ?
                              $signed((8'hb9)) : wire565))) : $signed((!$signed($signed((7'h40))))));
              reg627 = {$unsigned($unsigned((8'ha9)))};
              reg628 <= (^$signed(reg625));
              reg629 = ((+($signed((reg623 - reg621)) > reg581)) >> $signed($signed((reg623[(4'h8):(2'h3)] >= $unsigned(reg624)))));
            end
          for (forvar630 = (1'h0); (forvar630 < (3'h6)); forvar630 = (forvar630 + (1'h1)))
            begin
              reg631 <= (!reg567[(5'h14):(3'h5)]);
              reg632 <= (((!reg579) ?
                      {((reg623 ? reg582 : (7'h51)) ?
                              reg624[(2'h2):(1'h0)] : reg592[(4'hb):(3'h6)]),
                          (reg597 <= (reg588 + reg624))} : (forvar630 > reg595[(4'hc):(3'h6)])) ?
                  reg626 : $signed(reg591[(3'h4):(1'h1)]));
              reg633 <= $signed((!reg568));
              reg634 <= $unsigned(((wire565[(2'h2):(1'h1)] << $signed(reg582[(3'h4):(2'h3)])) ?
                  ({(reg621 && reg595), $signed(reg617), $signed(wire565)} ?
                      {$signed(wire565)} : reg566[(4'h8):(1'h1)]) : $signed(reg588)));
            end
          if ((($unsigned($signed(reg590)) || $signed($signed(wire562[(1'h1):(1'h1)]))) ?
              reg622[(4'hd):(4'h8)] : reg632))
            begin
              reg635 = $signed({$signed(((+reg576) + reg629)),
                  $unsigned(reg590),
                  reg621[(5'h1d):(5'h14)]});
            end
          else
            begin
              reg635 = $unsigned((~^$signed(reg634)));
              reg636 <= {(^(reg634[(3'h4):(2'h3)] > reg612))};
              reg637 <= ($unsigned((~&reg632)) ?
                  $unsigned((reg597 ?
                      (reg590 | wire564[(4'hd):(4'hd)]) : $signed(reg616))) : ($signed({reg624[(1'h0):(1'h0)],
                      ((8'hae) ? (8'hae) : reg601)}) + wire563[(1'h0):(1'h0)]));
            end
          if ($signed(reg627))
            begin
              reg638 <= $unsigned(reg579);
              reg639 <= {$unsigned(reg591)};
              reg640 = reg623;
              reg641 <= {((({reg573, reg632, (8'ha5)} ^~ {reg628}) ?
                      $unsigned((8'hbe)) : (~&reg617[(1'h0):(1'h0)])) | reg588[(1'h0):(1'h0)]),
                  ($unsigned(((reg582 <<< reg595) >> $signed((7'h4f)))) & ((~^{reg567,
                          (8'hb9),
                          wire565}) ?
                      $signed({reg620, reg612, reg619}) : (^(7'h56))))};
              reg642 <= {reg572,
                  (~|$signed(reg581[(1'h1):(1'h0)])),
                  $unsigned(reg576)};
            end
          else
            begin
              reg640 = {((~|$unsigned($signed(reg591))) != (+reg601)), reg625};
              reg641 <= (($unsigned($unsigned((^reg636))) ?
                      {{$unsigned(reg591), $unsigned(reg573), $signed(reg635)},
                          $signed(reg624)} : ((~|wire562) < (~|(!reg637)))) ?
                  {(((reg639 * (8'h9f)) ?
                              (reg616 ?
                                  reg629 : reg636) : (wire615 >> reg617)) ?
                          $unsigned({reg638,
                              reg591}) : ($signed(reg573) && reg588)),
                      $signed($unsigned((reg640 != reg590))),
                      (wire565[(1'h1):(1'h0)] >= reg567[(4'hb):(4'h8)])} : (+$signed((7'h46))));
              reg642 <= (~|reg626);
              reg643 <= ({$unsigned(((reg582 * wire563) >= (+reg597)))} ^~ (($signed($signed(reg597)) ?
                      reg626 : ((~|reg582) || $signed((7'h47)))) ?
                  reg582[(1'h0):(1'h0)] : (&$unsigned((wire605 ?
                      (7'h45) : wire615)))));
              reg644 <= (~|reg627);
              reg645 = (wire565 ?
                  {(reg634[(2'h3):(1'h0)] ?
                          reg581[(5'h1a):(4'h8)] : (&reg572))} : (~|((8'hac) ^ $unsigned($unsigned(reg601)))));
            end
        end
      else
        begin
          reg619 = ({((+((7'h42) ? reg592 : reg624)) ? (~&(8'hbf)) : reg645)} ?
              reg637 : $unsigned((^(!wire565))));
          reg621 <= $unsigned((forvar630[(4'h9):(2'h3)] ?
              reg570[(5'h19):(3'h5)] : {$unsigned({reg639})}));
          reg622 = ($signed(reg617[(4'ha):(4'ha)]) ?
              ($signed((reg579[(4'he):(1'h1)] ?
                  $signed((7'h4c)) : reg624[(4'h9):(3'h7)])) & (~|reg568[(5'h18):(4'hb)])) : (~|(~&$unsigned($unsigned(wire562)))));
          if ($signed(($unsigned((~&$unsigned(wire562))) * $unsigned($unsigned((reg601 ?
              reg642 : reg645))))))
            begin
              reg623 <= $unsigned(((~wire604[(4'h8):(1'h1)]) >>> reg624[(3'h6):(3'h4)]));
            end
          else
            begin
              reg623 <= ($signed(reg636[(5'h13):(3'h7)]) ?
                  wire605 : $signed(reg638[(4'h9):(1'h1)]));
            end
          if ({reg624,
              {(~^(wire563 ^ {wire605})),
                  (-$unsigned(((7'h58) ? reg590 : (8'ha2))))},
              reg590[(5'h11):(4'ha)]})
            begin
              reg624 = ($unsigned(($unsigned(reg566[(1'h1):(1'h1)]) ?
                      ((reg597 >>> reg571) == wire562) : $unsigned((^reg625)))) ?
                  reg620 : ({reg590, (7'h4f), (|(^~(8'h9e)))} ?
                      $signed(((reg574 ?
                          reg645 : reg632) >>> reg576)) : wire562[(3'h6):(2'h3)]));
              reg626 = (^$signed({reg621,
                  $signed($signed(wire562)),
                  ($unsigned(reg579) ?
                      (reg603 != reg629) : (reg634 ? reg597 : reg624))}));
              reg628 <= $unsigned($signed(($signed((!reg616)) ~^ ((reg619 < (8'hb0)) ^ wire562))));
              reg630 <= $unsigned(reg618);
              reg635 = $signed((({$unsigned(reg628)} ?
                      $unsigned({reg631,
                          forvar630,
                          reg570}) : $unsigned($signed(reg618))) ?
                  ({((8'hb7) && reg618)} & ({reg626, wire564, (8'hba)} ?
                      $signed(reg579) : {wire565,
                          reg622,
                          reg626})) : reg643[(4'hf):(1'h1)]));
              reg636 <= reg568[(3'h5):(1'h1)];
            end
          else
            begin
              reg624 = ($signed(reg628[(5'h16):(3'h6)]) ?
                  (wire604[(5'h12):(3'h4)] ^~ reg588) : $signed($unsigned((8'h9e))));
              reg626 = ($signed($unsigned((reg570[(4'hf):(3'h4)] ?
                  (reg639 ?
                      (8'ha4) : (8'hb8)) : (~^reg617)))) & $signed({((-reg603) ?
                      (^reg612) : $unsigned(reg620)),
                  reg626,
                  $signed({reg634})}));
              reg628 <= $unsigned($unsigned($signed(reg568[(4'h9):(2'h3)])));
            end
        end
      reg646 <= reg636[(5'h10):(2'h3)];
      for (forvar647 = (1'h0); (forvar647 < (3'h6)); forvar647 = (forvar647 + (1'h1)))
        begin
          for (forvar648 = (1'h0); (forvar648 < (1'h1)); forvar648 = (forvar648 + (1'h1)))
            begin
              reg649 <= reg597[(3'h6):(1'h1)];
              reg650 <= ($unsigned((~^($unsigned(reg588) ?
                  reg571[(1'h0):(1'h0)] : reg601))) > $unsigned((-(|$signed(reg597)))));
            end
          if (wire615)
            begin
              reg651 = $unsigned($signed($unsigned((reg630 ?
                  reg633[(5'h10):(3'h7)] : reg591[(2'h3):(2'h3)]))));
              reg652 <= ($unsigned((($unsigned((8'ha3)) > (reg628 * reg579)) & {(reg629 ^~ reg572)})) != (^~(wire563[(1'h1):(1'h0)] >> $unsigned((reg592 ?
                  reg616 : reg651)))));
              reg653 <= forvar647;
              reg654 = (-$signed((reg612[(3'h7):(3'h5)] - $signed((~^reg634)))));
              reg655 = (reg629 > (!(reg630 != $signed((~reg618)))));
              reg656 = (~^$signed((($signed(reg592) ?
                      $unsigned(reg644) : (8'ha2)) ?
                  ((wire615 == wire605) ^ $unsigned(reg635)) : $unsigned($unsigned((8'hb1))))));
            end
          else
            begin
              reg651 = (reg642[(5'h12):(3'h5)] ?
                  (8'ha6) : ((^wire562) ?
                      (($signed(reg628) >> (^(8'hbe))) ?
                          reg638 : reg628) : ((wire562[(1'h0):(1'h0)] + $unsigned(reg603)) ?
                          (&$unsigned(reg636)) : (~^(+reg567)))));
              reg654 = (&(+(&(~$signed(reg653)))));
            end
          reg657 <= $signed(reg629);
          reg658 <= (^reg566[(4'he):(2'h3)]);
          reg659 = $signed((&{($unsigned(reg626) ? reg649 : reg621),
              (((7'h54) ? reg597 : reg654) ?
                  $signed(reg567) : $signed(wire562))}));
          for (forvar660 = (1'h0); (forvar660 < (1'h0)); forvar660 = (forvar660 + (1'h1)))
            begin
              reg661 = $signed($signed($signed(((reg579 << (7'h4c)) > $unsigned((8'hae))))));
              reg662 = $signed($signed($unsigned(reg651)));
              reg663 <= $unsigned(reg643[(1'h1):(1'h1)]);
              reg664 = $signed($unsigned(reg628[(4'hc):(4'h8)]));
            end
        end
      if ({(8'hb3), (~&reg662[(4'h8):(3'h5)])})
        begin
          for (forvar665 = (1'h0); (forvar665 < (3'h4)); forvar665 = (forvar665 + (1'h1)))
            begin
              reg666 = ($unsigned(($unsigned(reg632[(1'h1):(1'h1)]) ?
                      reg591 : ((~^reg664) != $unsigned(reg651)))) ?
                  ($unsigned(reg576) ^~ wire565) : ($signed((~^(reg612 > reg642))) ?
                      (~|reg633[(2'h2):(2'h2)]) : (~reg663)));
            end
          for (forvar667 = (1'h0); (forvar667 < (2'h2)); forvar667 = (forvar667 + (1'h1)))
            begin
              reg668 <= reg574;
              reg669 <= ((reg577[(3'h7):(3'h7)] <<< forvar630) >= ($signed($unsigned($unsigned(reg603))) == ((~|(reg619 & reg625)) || {reg639[(3'h4):(3'h4)],
                  reg642[(5'h18):(5'h18)],
                  (reg661 ? reg639 : reg621)})));
              reg670 <= (!$unsigned((-$signed(reg624[(3'h5):(3'h4)]))));
              reg671 = $unsigned((((((8'h9f) ?
                      reg652 : reg622) >= reg624[(2'h3):(1'h0)]) != (((7'h58) ?
                      reg574 : reg632) * (forvar647 ? (8'hae) : forvar665))) ?
                  $signed(((forvar647 || reg634) ?
                      ((7'h55) ?
                          wire565 : reg628) : $unsigned(reg662))) : ({reg603,
                      reg627[(5'h17):(4'hb)],
                      (reg662 != reg582)} == $unsigned({wire604,
                      wire615,
                      reg624}))));
              reg672 = $unsigned({(((reg668 ? (8'h9f) : reg662) != (reg639 ?
                      (8'hac) : (8'hb9))) << $signed(reg626[(1'h1):(1'h0)])),
                  $signed($signed((reg627 ? reg573 : (8'hba)))),
                  ({forvar630, (reg651 || (8'hb2))} - reg592)});
              reg673 = reg570;
            end
          for (forvar674 = (1'h0); (forvar674 < (3'h4)); forvar674 = (forvar674 + (1'h1)))
            begin
              reg675 <= $unsigned(($signed($signed(reg649[(1'h1):(1'h0)])) ?
                  {{(~&reg621)}, ((~reg638) >>> reg624), reg643} : (!reg650)));
              reg676 = reg656[(4'h9):(3'h4)];
              reg677 <= $unsigned((-$signed((reg612[(2'h2):(1'h1)] ?
                  $unsigned(forvar630) : (reg662 ? reg628 : reg632)))));
              reg678 <= reg619[(3'h4):(2'h2)];
              reg679 <= (reg595[(3'h4):(1'h1)] <= reg675[(3'h5):(1'h1)]);
              reg680 <= reg567[(3'h4):(1'h0)];
            end
          reg681 = $unsigned((((reg633[(4'hd):(4'h9)] ?
              (wire604 == reg591) : (~reg638)) + ({wire563} & {reg680,
              (7'h49)})) && {($unsigned(reg626) ?
                  (reg628 ? reg595 : reg646) : reg634)}));
          reg682 = (reg629[(4'ha):(3'h5)] ? reg635 : reg664[(4'ha):(2'h3)]);
        end
      else
        begin
          if ((-{reg681[(3'h4):(1'h0)],
              ((reg651[(2'h3):(1'h0)] ?
                  {reg631, reg627, reg668} : reg597) <<< reg651[(3'h4):(3'h4)]),
              reg671[(5'h12):(4'hd)]}))
            begin
              reg665 = (^$signed($signed(reg678)));
              reg666 = reg616;
            end
          else
            begin
              reg667 <= ($unsigned((reg627 ?
                      $signed(reg656[(3'h6):(3'h4)]) : $signed($signed(forvar648)))) ?
                  ({$signed($signed(reg680)),
                      $signed(reg645),
                      $signed((reg680 != reg603))} && ((&{reg581,
                      reg641}) ~^ $signed(reg675[(3'h7):(2'h3)]))) : (8'hbe));
              reg668 <= reg582[(2'h2):(2'h2)];
              reg671 = (forvar665 ?
                  reg577 : $unsigned($unsigned(reg679[(1'h0):(1'h0)])));
              reg672 = (((7'h4b) > ({(~^reg630),
                  (~&reg635)} <<< reg632)) + (~^wire615[(4'hf):(1'h0)]));
              reg674 <= $signed({$signed(((&(8'hae)) ?
                      (-(7'h47)) : (reg591 ? reg669 : forvar660)))});
            end
        end
      for (forvar683 = (1'h0); (forvar683 < (3'h6)); forvar683 = (forvar683 + (1'h1)))
        begin
          for (forvar684 = (1'h0); (forvar684 < (2'h3)); forvar684 = (forvar684 + (1'h1)))
            begin
              reg685 <= ((reg653[(3'h4):(3'h4)] ~^ reg655[(4'h8):(3'h7)]) ?
                  $unsigned($unsigned(reg664[(3'h7):(3'h5)])) : $unsigned((7'h56)));
            end
          if (reg616[(1'h1):(1'h0)])
            begin
              reg686 = reg635[(4'ha):(1'h1)];
              reg687 = {{$unsigned({(reg643 ? reg581 : reg568)}),
                      $signed(reg590[(5'h10):(3'h4)]),
                      ($unsigned((~reg656)) ?
                          ((-reg626) ^ $signed((8'h9e))) : reg629[(3'h7):(3'h5)])}};
            end
          else
            begin
              reg686 = $signed((^($signed({(8'h9d), (8'hb6), reg652}) ?
                  $signed(wire564) : $signed(forvar684[(4'h8):(3'h6)]))));
              reg687 = $unsigned((^~($unsigned($signed(reg646)) ?
                  ($signed((8'hbf)) && forvar648[(3'h6):(2'h2)]) : (~&$signed(reg677)))));
              reg688 = {(8'ha7)};
              reg689 = (8'hb1);
              reg690 <= reg641;
              reg691 <= reg632;
              reg692 <= $unsigned(((reg592 ?
                      {reg632} : $signed(reg646[(4'hb):(4'h9)])) ?
                  {reg568[(1'h1):(1'h0)],
                      ((reg590 ? reg623 : reg631) ?
                          (~wire562) : (reg623 ?
                              reg679 : wire615))} : $signed($signed(((8'hb9) >> reg685)))));
            end
          if ((($unsigned($unsigned(forvar684[(2'h2):(1'h0)])) ?
                  (reg570 ^ (8'hba)) : reg643) ?
              (8'hb3) : (7'h48)))
            begin
              reg693 <= (^~$unsigned(reg621[(4'hd):(4'hc)]));
            end
          else
            begin
              reg694 = reg678[(4'h9):(3'h4)];
              reg695 <= {(+reg694)};
              reg696 <= (~&forvar630[(4'hb):(2'h3)]);
              reg697 <= ($signed({(+reg581),
                  reg592[(4'he):(4'he)],
                  reg619[(2'h3):(2'h3)]}) + (~|reg622[(4'he):(3'h7)]));
              reg698 = (reg641 * $unsigned({(reg566[(3'h5):(1'h1)] && reg678[(5'h19):(5'h11)])}));
              reg699 = (~reg650[(3'h7):(3'h4)]);
            end
          reg700 = $unsigned((forvar648 && $signed(reg622)));
          reg701 = $signed(reg645[(5'h13):(4'h9)]);
        end
    end
  module702 #() modinst1069 (wire1068, clk, reg669, reg678, reg582, reg637);
  assign wire1070 = ((reg567 || reg572[(3'h6):(2'h3)]) ?
                        ($signed(reg597) << reg638[(4'h9):(2'h2)]) : $unsigned((~$signed({reg618}))));
  assign wire1071 = (^~($signed((&(&wire604))) * (((wire564 ^~ reg592) ?
                        (+(7'h4f)) : (reg670 ?
                            reg597 : reg693)) << (reg668 * (reg588 ^~ reg696)))));
  assign wire1072 = reg595;
  assign wire1073 = ({$signed(((^reg576) ? (^~reg570) : $signed(reg577))),
                        reg588[(2'h2):(1'h1)]} || reg581[(4'hd):(1'h0)]);
  always
    @(posedge clk) begin
      if (((8'hbb) ?
          ($unsigned($unsigned({reg642,
              reg634,
              reg618})) == $unsigned(((^(7'h55)) ?
              reg691 : (8'haf)))) : reg595))
        begin
          if ($unsigned($signed((7'h4c))))
            begin
              reg1074 = reg576;
              reg1075 = reg631[(3'h4):(3'h4)];
              reg1076 = reg644;
              reg1077 <= $unsigned((((~^reg591) ?
                      (|reg657[(5'h11):(4'h9)]) : $unsigned(reg658)) ?
                  wire605 : reg567[(5'h12):(5'h11)]));
              reg1078 = (reg1076 ?
                  (!$unsigned($signed(((8'ha3) << wire563)))) : reg636[(3'h4):(2'h3)]);
              reg1079 = wire1068;
            end
          else
            begin
              reg1074 = reg650[(3'h7):(3'h7)];
              reg1077 <= reg636;
              reg1078 = $unsigned(reg592[(3'h5):(1'h0)]);
              reg1079 = ((!(+({(7'h45), reg570} == $signed(wire1068)))) ?
                  $signed(reg621) : $signed($unsigned(({reg653,
                      reg636,
                      reg677} << $signed(reg582)))));
            end
          reg1080 = {(reg696[(3'h4):(3'h4)] ?
                  $unsigned($signed(reg636[(1'h0):(1'h0)])) : (reg603 ?
                      $signed(reg644[(5'h1c):(4'ha)]) : ($unsigned((8'hbe)) > $signed(reg590)))),
              $signed(reg649[(4'h8):(2'h3)])};
        end
      else
        begin
          for (forvar1074 = (1'h0); (forvar1074 < (1'h1)); forvar1074 = (forvar1074 + (1'h1)))
            begin
              reg1075 = ($signed($signed(reg685[(3'h6):(3'h4)])) ?
                  (~|(8'hbc)) : reg576);
              reg1076 = {{$unsigned(({wire615} ? (8'hbd) : (~|(8'h9d)))),
                      (($signed(reg590) ^ reg680[(2'h3):(2'h3)]) || $unsigned($unsigned(reg652))),
                      reg643},
                  $signed($signed(((forvar1074 ? reg567 : wire1072) ?
                      reg642 : (reg1075 ? forvar1074 : reg623)))),
                  $signed(reg636)};
              reg1077 <= $signed({(~$signed(reg618[(4'hd):(2'h3)]))});
            end
        end
      reg1081 <= reg697[(4'hf):(4'h9)];
      for (forvar1082 = (1'h0); (forvar1082 < (3'h5)); forvar1082 = (forvar1082 + (1'h1)))
        begin
          reg1083 <= $unsigned(wire1070);
        end
      reg1084 = reg590[(5'h14):(4'hb)];
      if ({{reg642[(5'h14):(4'h8)],
              $unsigned(((reg574 >= reg668) ?
                  reg658[(3'h4):(3'h4)] : reg568[(5'h17):(5'h12)])),
              ($signed((reg642 ?
                  wire1072 : reg1084)) & wire1070[(5'h10):(4'hd)])},
          {reg644[(4'hc):(4'ha)],
              (~^reg566[(4'ha):(3'h5)]),
              reg639[(4'ha):(1'h1)]}})
        begin
          for (forvar1085 = (1'h0); (forvar1085 < (2'h3)); forvar1085 = (forvar1085 + (1'h1)))
            begin
              reg1086 <= reg574[(5'h13):(4'he)];
              reg1087 = (+(reg669 ?
                  $unsigned(reg695[(5'h13):(3'h6)]) : reg674[(1'h1):(1'h1)]));
              reg1088 = {wire1073,
                  ((((reg670 << reg588) << (8'ha8)) ?
                          ({wire605,
                              reg601,
                              reg678} && $signed(reg650)) : {reg693[(3'h4):(1'h0)],
                              $unsigned((7'h52)),
                              $signed(reg577)}) ?
                      (|(&$signed((7'h55)))) : ((^~reg675[(2'h3):(2'h3)]) >= wire563))};
            end
        end
      else
        begin
          reg1085 = $unsigned(reg658[(3'h6):(2'h2)]);
          reg1086 <= $unsigned(($signed(((reg680 ^ reg652) ?
                  reg603[(2'h3):(1'h1)] : ((7'h4a) ? reg616 : (7'h56)))) ?
              $unsigned(((reg1088 & reg1076) != $signed(reg590))) : $signed({(8'ha8)})));
          reg1087 = (^$unsigned($signed($signed($unsigned(reg690)))));
          reg1089 <= reg649[(2'h2):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      reg1090 <= $signed($unsigned(($signed($unsigned((7'h51))) ?
          (reg577[(1'h0):(1'h0)] ?
              (reg618 ? (7'h40) : wire1068) : ((8'ha6) ?
                  reg680 : wire563)) : $unsigned((reg1077 * reg570)))));
      if ((wire604 << (&($signed($unsigned(reg678)) ?
          (reg618 != reg675[(4'h8):(1'h1)]) : reg679[(3'h4):(1'h1)]))))
        begin
          if (reg633)
            begin
              reg1091 = $unsigned(($unsigned(reg649[(2'h3):(1'h0)]) * reg690));
            end
          else
            begin
              reg1092 <= $signed($unsigned($unsigned(reg695[(5'h15):(4'h9)])));
              reg1093 <= (reg663 <<< {($signed($signed(reg597)) ^ (reg677[(4'hf):(1'h1)] ?
                      {reg630, reg571} : ((8'hba) + reg574))),
                  {$signed((reg674 ^ (8'hbd))),
                      reg632[(2'h3):(1'h0)],
                      $unsigned({(8'ha0)})}});
              reg1094 <= (({reg630,
                      ((reg1089 ? reg663 : wire565) ?
                          reg668 : ((8'ha2) ?
                              reg668 : reg579))} ~^ ($unsigned((reg601 ?
                      reg577 : reg680)) >> {reg1090})) ?
                  ((~&$signed((^(8'hba)))) ^~ (~^((reg663 ?
                      reg693 : (8'ha3)) & (reg642 == reg628)))) : (7'h42));
              reg1095 <= ((^~$unsigned((^(^~reg628)))) >>> $unsigned({reg634,
                  {reg1086[(4'hb):(3'h7)]}}));
              reg1096 = $unsigned({$unsigned((~&$signed(reg1090))),
                  (^~reg633[(5'h19):(4'hd)]),
                  reg601[(4'h9):(3'h6)]});
              reg1097 <= (|reg590[(4'h8):(3'h6)]);
            end
        end
      else
        begin
          for (forvar1091 = (1'h0); (forvar1091 < (1'h1)); forvar1091 = (forvar1091 + (1'h1)))
            begin
              reg1092 <= $unsigned(reg638[(4'h8):(1'h1)]);
              reg1096 = reg588;
              reg1097 <= {(reg570 ?
                      {reg675,
                          (reg625 ?
                              $signed((7'h4c)) : reg630)} : $signed({(~&(7'h52)),
                          (reg625 ? (8'ha5) : reg649)})),
                  (reg581 != (reg566[(3'h4):(3'h4)] ?
                      $unsigned((+reg677)) : $unsigned($signed(wire562))))};
            end
          reg1098 <= (7'h58);
          for (forvar1099 = (1'h0); (forvar1099 < (1'h0)); forvar1099 = (forvar1099 + (1'h1)))
            begin
              reg1100 <= (^~$unsigned((!reg639)));
              reg1101 = reg595;
              reg1102 <= $signed((reg595[(4'hb):(3'h6)] ?
                  (~&reg1097[(3'h5):(1'h0)]) : $signed((~^reg588[(2'h2):(2'h2)]))));
              reg1103 = ($signed((wire565 == (&$unsigned(wire1068)))) <= $unsigned($signed(((reg582 ?
                  reg621 : reg1100) || wire562[(3'h5):(3'h5)]))));
            end
          reg1104 <= reg697[(4'h8):(1'h1)];
        end
      reg1105 <= reg679[(3'h4):(1'h0)];
      reg1106 <= ((($signed(reg574[(4'he):(1'h1)]) ?
              $signed((8'hab)) : $unsigned((~&(8'ha3)))) ?
          reg570[(5'h11):(3'h4)] : reg591) - ((7'h4d) && {$signed(reg693),
          $signed(reg632),
          wire1068[(4'ha):(3'h5)]}));
      for (forvar1107 = (1'h0); (forvar1107 < (1'h0)); forvar1107 = (forvar1107 + (1'h1)))
        begin
          reg1108 <= reg641[(4'h9):(3'h4)];
          reg1109 = $signed(($signed(((|reg674) >> (~wire615))) <<< ({$signed(reg571),
                  $signed((8'hbb))} ?
              (reg601[(5'h16):(5'h11)] ?
                  reg680[(3'h5):(2'h2)] : reg642[(4'hf):(4'hd)]) : (((7'h42) ?
                  reg573 : reg579) & (-wire604)))));
        end
    end
  assign wire1110 = ($signed($signed((~&reg590[(4'ha):(3'h7)]))) <= ((({reg643,
                                reg653,
                                reg1089} ?
                            (reg577 | reg603) : $unsigned(reg653)) >>> ((~^reg612) ?
                            (reg642 <<< wire563) : $unsigned(reg674))) ?
                        (8'hbb) : $signed($signed($signed(reg650)))));
  always
    @(posedge clk) begin
      if ((&((((wire615 && wire605) ~^ ((7'h41) ? reg1106 : reg579)) ?
          reg675 : $signed(reg697[(1'h0):(1'h0)])) || reg675[(2'h3):(2'h3)])))
        begin
          reg1111 = (((((!reg1102) <= (~wire1071)) ?
                  (7'h40) : $signed(reg582)) ?
              wire604 : (~reg571)) > reg646);
          reg1112 = $signed($unsigned(reg1104[(5'h15):(4'he)]));
        end
      else
        begin
          if ((^~($unsigned(($unsigned((7'h44)) ? $signed(wire1070) : reg634)) ?
              (($signed(reg641) >> reg685) ?
                  $unsigned(reg571) : $unsigned((reg571 + reg644))) : $unsigned(reg679[(4'h8):(2'h2)]))))
            begin
              reg1113 <= ((+(((reg652 & reg690) ?
                      (reg1090 < wire1070) : (-(7'h47))) & ((reg623 ?
                      reg650 : reg667) * (~reg650)))) ?
                  reg685 : (~reg568[(3'h7):(2'h3)]));
            end
          else
            begin
              reg1113 <= ((reg642 >> reg576) ?
                  ({{$signed(reg1089)}} ^~ ($signed((reg657 ?
                      (7'h51) : reg595)) ~^ reg643)) : $unsigned(reg646));
            end
        end
      for (forvar1114 = (1'h0); (forvar1114 < (1'h0)); forvar1114 = (forvar1114 + (1'h1)))
        begin
          for (forvar1115 = (1'h0); (forvar1115 < (2'h2)); forvar1115 = (forvar1115 + (1'h1)))
            begin
              reg1116 = ((8'ha6) <<< reg690);
              reg1117 = reg1086;
            end
          reg1118 <= $unsigned($unsigned(($signed($unsigned(reg597)) - ($signed(reg588) <<< $unsigned(reg1100)))));
          reg1119 = $signed($signed(((reg674 >> wire1110[(3'h6):(3'h5)]) + ((~reg1100) ?
              reg576 : wire565))));
        end
      for (forvar1120 = (1'h0); (forvar1120 < (3'h4)); forvar1120 = (forvar1120 + (1'h1)))
        begin
          reg1121 <= reg669[(2'h3):(2'h3)];
          for (forvar1122 = (1'h0); (forvar1122 < (3'h5)); forvar1122 = (forvar1122 + (1'h1)))
            begin
              reg1123 = {$signed((({(7'h4f), reg1092, (8'h9d)} ?
                      (reg643 > (8'had)) : {(8'ha3),
                          (7'h4e),
                          reg644}) || ((&reg670) ? {reg646} : (^~reg632))))};
              reg1124 = {$signed(reg625), reg625[(2'h2):(1'h1)]};
              reg1125 = ($signed((reg591[(3'h6):(3'h4)] ?
                      ({reg566} != $signed((8'hb7))) : ({reg1102,
                          reg1097,
                          (7'h44)} ~^ $unsigned(forvar1114)))) ?
                  reg643[(5'h14):(3'h4)] : (!{($unsigned((8'h9c)) < $unsigned((8'ha3))),
                      reg591[(4'h9):(3'h5)]}));
              reg1126 <= ((|(7'h48)) ?
                  ($signed(wire605[(5'h13):(3'h6)]) ^ (&(~|{reg595,
                      reg670,
                      reg690}))) : reg630);
              reg1127 = reg574;
            end
        end
      reg1128 = (~|(reg618[(3'h4):(3'h4)] ?
          reg668 : $signed(reg669[(5'h12):(4'h9)])));
      if ((~^wire1070))
        begin
          reg1129 = $unsigned((8'ha9));
          reg1130 <= ((reg1112 ?
                  {(reg568[(4'ha):(4'h9)] < {reg679, reg572}),
                      $signed((reg677 ? reg644 : reg643)),
                      $unsigned((reg1127 ?
                          reg1090 : reg577))} : $unsigned($unsigned((-(7'h46))))) ?
              $signed($signed($signed(reg1121))) : $signed(reg658[(2'h3):(2'h2)]));
          reg1131 <= $signed($unsigned(reg667));
          reg1132 <= (!reg691);
          for (forvar1133 = (1'h0); (forvar1133 < (1'h1)); forvar1133 = (forvar1133 + (1'h1)))
            begin
              reg1134 = reg1090;
              reg1135 = reg616[(5'h13):(5'h13)];
            end
          if ($unsigned(reg675))
            begin
              reg1136 = {(&(-((reg1123 ^~ forvar1122) | (~&reg612)))),
                  $unsigned(reg621)};
              reg1137 <= (forvar1114[(1'h0):(1'h0)] == reg573);
              reg1138 = (reg1134 ?
                  $signed(reg1119[(3'h4):(2'h2)]) : (reg674 | $unsigned(((|reg591) ~^ (reg1105 == forvar1115)))));
            end
          else
            begin
              reg1136 = $signed($signed($signed(reg1124)));
              reg1137 <= $signed(reg634[(2'h2):(2'h2)]);
              reg1139 <= {reg695,
                  ($unsigned((7'h52)) != (-$signed((reg1137 && reg650)))),
                  {reg603[(2'h3):(1'h0)], reg638[(3'h4):(3'h4)]}};
              reg1140 <= reg1121;
            end
        end
      else
        begin
          for (forvar1129 = (1'h0); (forvar1129 < (1'h1)); forvar1129 = (forvar1129 + (1'h1)))
            begin
              reg1130 <= ((reg639 ?
                      ((!$unsigned(reg1108)) * $unsigned(reg1129[(2'h3):(2'h2)])) : ($unsigned((reg649 ?
                              (7'h54) : reg1105)) ?
                          $unsigned($signed(reg1102)) : {$signed(reg1116),
                              reg574[(2'h3):(1'h1)]})) ?
                  {((~^(reg674 ? reg668 : reg658)) ?
                          reg677 : $unsigned(reg1113)),
                      (~((~&wire1071) ? (reg663 < (7'h4e)) : $signed((8'h9d)))),
                      {$unsigned((~reg1089))}} : $unsigned(reg1118));
              reg1131 <= (reg646 ?
                  $signed($unsigned(((reg675 < reg1105) >>> reg603[(2'h2):(1'h0)]))) : {reg638,
                      ((~&$unsigned(reg1077)) ?
                          {$unsigned(reg677)} : $signed((reg657 ?
                              reg644 : (8'hab)))),
                      $unsigned(reg630[(2'h3):(2'h3)])});
              reg1133 = $unsigned({reg574,
                  ({$signed((7'h42)),
                          (reg601 ? reg1092 : reg1118),
                          $unsigned(reg571)} ?
                      (~|$signed(reg618)) : reg1095[(3'h4):(1'h1)]),
                  (7'h45)});
              reg1134 = (+reg638[(3'h6):(3'h4)]);
              reg1137 <= reg1108;
            end
          reg1138 = ($signed($signed($signed((reg1077 * reg618)))) ?
              $signed((~|wire565)) : $signed(reg693[(3'h7):(3'h6)]));
          for (forvar1139 = (1'h0); (forvar1139 < (1'h1)); forvar1139 = (forvar1139 + (1'h1)))
            begin
              reg1140 <= reg577[(1'h0):(1'h0)];
              reg1141 <= $unsigned($unsigned((((|reg633) ?
                  wire563 : (~|reg669)) != reg1113[(2'h2):(2'h2)])));
              reg1142 = $unsigned(wire604[(3'h4):(3'h4)]);
              reg1143 = $unsigned(reg1118[(4'h8):(3'h6)]);
            end
          for (forvar1144 = (1'h0); (forvar1144 < (1'h1)); forvar1144 = (forvar1144 + (1'h1)))
            begin
              reg1145 = $signed(((((reg663 + (8'hb4)) ?
                  (reg1118 > reg1126) : (reg1086 ?
                      reg644 : reg1100)) >> reg690[(1'h1):(1'h1)]) - $unsigned((^~$signed(forvar1129)))));
              reg1146 = ((!reg572[(4'h9):(3'h7)]) ?
                  $unsigned($signed(reg1104)) : reg633);
              reg1147 <= (reg1095 ?
                  (7'h44) : $unsigned({($signed((8'hb9)) ?
                          $signed(reg1129) : {reg571, reg1128, reg570}),
                      (8'h9c)}));
              reg1148 = (($signed((|(reg1090 - reg1119))) ?
                  $signed(reg1118) : reg616[(5'h11):(4'h9)]) ~^ reg643[(2'h3):(2'h3)]);
              reg1149 = $signed(reg1128);
              reg1150 <= $signed((reg568 ?
                  $unsigned(reg1148[(5'h10):(3'h6)]) : reg1077));
            end
          if ((((~&wire1073[(4'hf):(1'h1)]) ?
                  $signed(reg1102) : (((|reg1138) * $unsigned(reg668)) ?
                      wire605 : reg1124[(4'he):(1'h1)])) ?
              ((7'h41) ?
                  $unsigned(forvar1122[(5'h12):(4'hb)]) : reg1102[(4'h8):(4'h8)]) : reg641))
            begin
              reg1151 = $unsigned((wire562 >= reg674));
            end
          else
            begin
              reg1152 <= (|forvar1129);
            end
        end
      for (forvar1153 = (1'h0); (forvar1153 < (1'h1)); forvar1153 = (forvar1153 + (1'h1)))
        begin
          reg1154 = (^reg566[(3'h6):(2'h3)]);
          if (reg679)
            begin
              reg1155 <= reg1108[(2'h2):(2'h2)];
              reg1156 <= {(|$signed($signed($unsigned(reg1095)))),
                  $unsigned($unsigned(reg1125[(2'h3):(2'h3)])),
                  reg576};
              reg1157 <= forvar1120;
              reg1158 = ({(reg631 ?
                          $signed(wire1072) : (reg650 ?
                              $signed((7'h54)) : reg680)),
                      $signed((^~$signed(reg1113)))} ?
                  ((((reg667 ? reg581 : reg1106) ?
                              (8'h9c) : {reg572, reg1090}) ?
                          ((reg643 ^~ forvar1114) ~^ {reg1125,
                              (8'hb1),
                              reg577}) : $unsigned((~|reg1086))) ?
                      ((reg649 ?
                          (wire565 & wire563) : $signed(reg1097)) <= $unsigned({reg652})) : ($unsigned(reg1155) ?
                          (reg612 ?
                              (~^reg1094) : {(8'hb8), (7'h54)}) : ({reg632} ?
                              (|reg650) : $signed(reg1131)))) : (reg1104[(4'hb):(2'h3)] && reg696[(3'h7):(2'h3)]));
              reg1159 = ((~^$signed(($signed(reg1147) << (reg616 ?
                      (8'hb7) : reg1089)))) ?
                  ((~(!$signed((8'hb6)))) != {((forvar1120 ?
                          reg643 : reg1077) | $unsigned(reg638)),
                      $signed(forvar1122[(5'h15):(2'h3)]),
                      (7'h4c)}) : reg1093);
              reg1160 <= (($signed(reg621[(5'h13):(5'h12)]) * {(reg628[(4'hf):(4'hd)] ?
                          forvar1115[(3'h4):(2'h2)] : $signed(reg633)),
                      {{(8'hb5), reg1106}, (~&reg1118)},
                      (&forvar1115[(1'h0):(1'h0)])}) ?
                  (&(-reg1093)) : ((8'hac) ?
                      wire562 : reg1102[(5'h12):(3'h6)]));
            end
          else
            begin
              reg1155 <= {($unsigned(reg1139) ?
                      reg1105[(3'h4):(2'h2)] : $unsigned($unsigned($signed((7'h58)))))};
              reg1156 <= reg601;
              reg1158 = $signed((-reg1116[(3'h6):(3'h5)]));
              reg1159 = (reg1141 ?
                  $unsigned({$unsigned((~reg588)),
                      (forvar1133[(1'h0):(1'h0)] >>> (reg577 ?
                          reg1098 : reg630)),
                      $signed($unsigned(wire563))}) : reg621);
              reg1160 <= reg643;
              reg1161 = (reg1158[(2'h2):(1'h1)] ?
                  (reg570 ?
                      $signed({$unsigned(wire565),
                          $signed(reg670)}) : {(+$unsigned(reg592)),
                          {(reg646 ? reg1136 : (8'ha9)),
                              $signed(reg1077),
                              $signed(reg592)}}) : ($unsigned(reg601) ?
                      (&($signed((7'h56)) ?
                          $signed(wire565) : (^~reg658))) : (^reg639)));
            end
          for (forvar1162 = (1'h0); (forvar1162 < (3'h4)); forvar1162 = (forvar1162 + (1'h1)))
            begin
              reg1163 <= $signed((reg634[(3'h4):(2'h2)] * (($unsigned(reg646) ?
                      $unsigned((8'hb5)) : (~&reg1119)) ?
                  {reg1158} : $unsigned(((7'h42) - reg653)))));
              reg1164 <= (reg628[(5'h10):(4'hb)] ?
                  $unsigned(($unsigned(wire1068[(5'h12):(3'h6)]) ?
                      $signed((-reg591)) : {(reg1138 ^ reg1077)})) : {reg570[(4'he):(4'hb)],
                      $unsigned({(reg634 + reg618), wire1072}),
                      $signed(((|wire562) * reg679[(4'ha):(3'h6)]))});
              reg1165 = (^reg592[(4'hf):(4'ha)]);
              reg1166 = (^(+$signed((reg1098 - ((7'h4e) ?
                  (8'hba) : (7'h46))))));
              reg1167 <= reg588[(1'h0):(1'h0)];
              reg1168 <= reg1124;
            end
          if ((reg1159[(1'h1):(1'h0)] & reg678))
            begin
              reg1169 = $signed(reg1117[(4'h8):(3'h7)]);
              reg1170 = $unsigned($unsigned({$signed(reg1081[(5'h12):(3'h4)])}));
              reg1171 <= (~&reg1090[(3'h5):(2'h3)]);
              reg1172 = reg1081;
              reg1173 <= $unsigned((+(reg576[(2'h2):(1'h0)] ?
                  {(reg674 ? reg1139 : reg1159),
                      (reg628 ?
                          reg1145 : (8'hb6))} : reg1128[(5'h11):(4'hf)])));
              reg1174 = ((&$signed($signed(reg1156[(4'h8):(3'h7)]))) && $signed(reg1102[(5'h10):(4'hb)]));
            end
          else
            begin
              reg1171 <= ({{{(reg1136 ? reg1152 : (8'hb3))},
                          $unsigned((~&reg1116)),
                          $signed(reg1098[(4'ha):(2'h2)])},
                      $unsigned(reg1138),
                      (($unsigned(reg566) ?
                              $signed(reg576) : {reg1151,
                                  wire1068,
                                  forvar1122}) ?
                          (7'h42) : $unsigned($signed(reg1139)))} ?
                  $signed($unsigned(reg652[(3'h7):(1'h1)])) : $signed(({{reg663,
                          reg1135,
                          forvar1153}} >> ((!reg1174) * (7'h54)))));
              reg1173 <= (~^$signed(reg1108[(5'h18):(4'h9)]));
              reg1175 <= reg1090;
            end
          reg1176 = reg646;
          reg1177 = (^~reg1118);
          for (forvar1178 = (1'h0); (forvar1178 < (3'h5)); forvar1178 = (forvar1178 + (1'h1)))
            begin
              reg1179 = $signed((~&reg649));
              reg1180 = reg1117;
              reg1181 <= reg1157;
              reg1182 <= {$signed(reg668[(4'h9):(2'h3)])};
              reg1183 = $unsigned(((((wire605 ? reg1102 : reg1136) ?
                  {reg601,
                      reg1155} : (reg1155 || reg631)) <<< reg597[(3'h4):(2'h3)]) + (~(8'hb0))));
              reg1184 = ((reg581 ?
                  $unsigned($unsigned($unsigned(reg1105))) : $signed($signed((!reg623)))) ^~ $signed((($signed(reg1134) > wire564) ?
                  ((reg1154 >> reg572) ?
                      reg1151[(1'h1):(1'h1)] : reg567) : (^~(8'had)))));
            end
        end
    end
  assign wire1185 = $signed(((-((reg636 ? reg633 : reg1126) >>> (reg571 ?
                        (8'hb7) : (8'haf)))) >>> (^~$signed(((7'h53) ?
                        reg695 : reg691)))));
  always
    @(posedge clk) begin
      if (reg685)
        begin
          if (reg632)
            begin
              reg1186 <= ((8'hbf) * reg590);
              reg1187 = reg1132;
              reg1188 <= (~|(({reg641[(3'h5):(3'h4)]} && $signed((wire565 != (7'h4b)))) >= (reg1092 ?
                  reg1094[(1'h0):(1'h0)] : $signed($unsigned(reg1077)))));
            end
          else
            begin
              reg1187 = reg590;
              reg1188 <= ((8'hb7) ?
                  {$unsigned((reg1187 <<< (&wire1070))),
                      $unsigned(reg1167[(3'h4):(1'h1)]),
                      ($signed(reg657[(4'hf):(2'h3)]) <= ($signed(reg690) ?
                          reg625 : reg1188[(2'h3):(2'h2)]))} : $unsigned((((~|reg1164) * reg678[(4'h9):(3'h7)]) ?
                      {$unsigned(wire564),
                          (reg639 ? reg1171 : reg590),
                          (reg571 == reg652)} : (~&reg1168[(4'hd):(3'h4)]))));
            end
          if (reg1171)
            begin
              reg1189 = (reg675[(4'h8):(3'h5)] <<< $unsigned(reg597));
              reg1190 = ((|({$signed(reg653),
                  $unsigned(reg1132),
                  (reg567 ?
                      wire1071 : reg592)} ^~ (reg1113 < {wire615}))) >= (+reg1139));
            end
          else
            begin
              reg1189 = (reg1126 ?
                  reg1150 : $signed(((-((7'h42) + reg643)) - ($unsigned(reg1150) ?
                      (|reg1094) : (~reg650)))));
              reg1191 <= $signed(((((!reg696) ~^ $signed(reg567)) ?
                      $signed($signed(reg588)) : $signed($unsigned(reg582))) ?
                  ((~^reg674) >> (~$unsigned(reg1164))) : (|(7'h57))));
              reg1192 = reg612[(4'he):(3'h4)];
              reg1193 = ($unsigned($signed($unsigned(reg693))) ^ ($unsigned($signed(wire1072[(4'h8):(3'h5)])) >= {$unsigned($signed(reg573)),
                  $signed((reg1106 ? reg1181 : (8'hae)))}));
              reg1194 <= $unsigned(($unsigned(($signed(reg1137) ?
                  {reg639, reg579} : (reg570 ?
                      reg612 : (7'h55)))) >= (+$signed((reg1140 ^ (8'hb9))))));
              reg1195 = (reg618[(4'h8):(4'h8)] & (($unsigned(reg573[(1'h1):(1'h1)]) >>> (^~reg1094[(5'h14):(1'h1)])) ?
                  (^{(reg597 < reg1126),
                      ((7'h54) ^ reg1168)}) : ((reg633[(3'h5):(2'h3)] ?
                      (~&reg1192) : reg621) * {reg1147[(3'h4):(2'h2)],
                      reg1092[(3'h4):(3'h4)],
                      (~&reg631)})));
            end
        end
      else
        begin
          reg1187 = $signed({(+$signed($signed(reg652))),
              (($unsigned(reg1086) * (^(7'h47))) ?
                  reg623 : $signed((reg637 && reg591)))});
          reg1188 <= (|reg1118[(4'hc):(1'h0)]);
          reg1191 <= (reg650 ? reg625 : wire1071);
          reg1194 <= (reg670 ?
              $signed($signed((reg1105 < reg1108))) : wire1070);
          if (reg571)
            begin
              reg1195 = $signed({reg690[(2'h2):(1'h0)],
                  $unsigned($signed({(8'ha7), (7'h53)})),
                  $unsigned({$signed((7'h41)), (wire564 >>> reg597)})});
              reg1196 = reg576[(2'h3):(2'h3)];
              reg1197 = wire1070[(5'h12):(4'h9)];
              reg1198 = reg572[(1'h1):(1'h0)];
            end
          else
            begin
              reg1195 = reg590;
              reg1199 <= (7'h54);
              reg1200 <= reg1108[(5'h10):(2'h2)];
              reg1201 <= reg601;
              reg1202 = $signed(reg1175);
              reg1203 = reg1105[(3'h4):(2'h2)];
              reg1204 = (~|$unsigned(((reg1140 * (reg1193 ? reg1104 : reg649)) ?
                  (wire1110 ?
                      (reg678 ?
                          reg597 : reg590) : (~^reg1094)) : ((reg597 < reg641) ?
                      (~|reg631) : (reg1194 & (7'h50))))));
            end
        end
      for (forvar1205 = (1'h0); (forvar1205 < (1'h1)); forvar1205 = (forvar1205 + (1'h1)))
        begin
          reg1206 <= (reg1167[(5'h12):(4'he)] ?
              (!reg591[(4'hd):(1'h0)]) : reg1118[(1'h0):(1'h0)]);
          for (forvar1207 = (1'h0); (forvar1207 < (3'h4)); forvar1207 = (forvar1207 + (1'h1)))
            begin
              reg1208 = (forvar1205[(1'h1):(1'h1)] ?
                  $unsigned(reg679[(4'ha):(3'h7)]) : ((reg601 < (reg642 ^~ $signed(reg1191))) ?
                      (($signed(reg690) ?
                              {(8'ha0), reg1201, reg1094} : (&forvar1205)) ?
                          {$signed(reg571),
                              reg644[(5'h17):(4'ha)]} : $signed($signed(reg582))) : {((reg646 >>> (8'hb4)) ?
                              (~&reg641) : (reg669 ^ reg1188)),
                          $unsigned($unsigned(reg588))}));
              reg1209 <= ((((-reg677[(2'h3):(1'h1)]) ?
                      $signed({(7'h57), reg643}) : (reg644 ?
                          reg1118 : $unsigned((7'h51)))) ?
                  reg1157[(3'h5):(1'h0)] : reg1077[(4'he):(3'h6)]) && ($unsigned(reg1186[(5'h10):(2'h3)]) ?
                  (~&{(reg639 ? reg1147 : reg571)}) : reg576));
              reg1210 <= $signed(($unsigned(reg642[(5'h12):(3'h5)]) ?
                  (reg1132[(5'h19):(4'h8)] - reg657[(4'hf):(3'h7)]) : $unsigned(reg1202)));
              reg1211 = ((!reg1193) ? (!reg579) : reg574[(3'h6):(3'h5)]);
              reg1212 = reg595;
              reg1213 <= $unsigned(reg628[(5'h10):(5'h10)]);
            end
          if ((($signed($unsigned($unsigned(reg695))) ?
                  ((reg668 ?
                      $signed((8'hb0)) : (|reg638)) ^~ reg1188) : $unsigned((^$signed((8'ha8))))) ?
              $unsigned(($unsigned($signed((8'hb8))) ?
                  ((reg1132 >>> (8'hb5)) ?
                      (reg642 - reg652) : $unsigned(reg1192)) : wire564)) : $signed((8'hbf))))
            begin
              reg1214 = (($signed({reg1196,
                      reg1098,
                      wire1068[(3'h7):(1'h0)]}) << $signed(reg1194[(4'he):(3'h7)])) ?
                  (~^reg667[(5'h12):(3'h5)]) : $unsigned($signed(reg1206[(5'h16):(5'h13)])));
              reg1215 = reg1190;
              reg1216 <= reg1163[(4'he):(3'h4)];
              reg1217 <= reg1152;
              reg1218 <= {$signed((((wire1185 ? reg675 : wire1073) ?
                          (~^(8'ha1)) : reg572[(3'h6):(2'h3)]) ?
                      reg693 : $signed((~&(7'h4f)))))};
            end
          else
            begin
              reg1214 = (-(reg668 - reg1104));
              reg1216 <= $signed(reg643);
              reg1217 <= $signed({$unsigned((^~(&reg1152))),
                  wire1185[(1'h0):(1'h0)]});
            end
          reg1219 <= $unsigned((-$unsigned({(wire1110 ? reg669 : reg1199),
              $signed(reg1214),
              reg630[(5'h12):(5'h10)]})));
        end
    end
  assign wire1220 = ($unsigned((reg1152 ^~ (8'ha9))) ?
                        $unsigned(((-(|reg631)) ?
                            $signed($signed(reg668)) : ((|reg631) ?
                                (~|reg1194) : wire615))) : ((($unsigned(reg582) ?
                                {reg1093} : (wire1110 <<< (7'h58))) || reg1081) ?
                            reg603 : ({$signed(reg668),
                                ((8'hae) & (7'h4e))} <= reg679[(1'h1):(1'h1)])));
  assign wire1221 = (reg1102[(1'h1):(1'h1)] ?
                        reg638[(3'h6):(3'h5)] : (reg670[(1'h0):(1'h0)] ?
                            {reg693,
                                {$signed((7'h45)),
                                    reg567}} : reg1106[(1'h1):(1'h0)]));
  always
    @(posedge clk) begin
      reg1222 = {{((~^$signed(wire615)) + $unsigned((|reg1201))),
              (|((reg1093 ? reg566 : (7'h52)) ?
                  $signed(wire1070) : (reg637 ? reg652 : reg590))),
              (+(+reg631))}};
      for (forvar1223 = (1'h0); (forvar1223 < (1'h0)); forvar1223 = (forvar1223 + (1'h1)))
        begin
          reg1224 <= $signed($unsigned((&($signed(reg658) << (8'hb8)))));
          for (forvar1225 = (1'h0); (forvar1225 < (2'h3)); forvar1225 = (forvar1225 + (1'h1)))
            begin
              reg1226 <= (reg696[(1'h0):(1'h0)] - ($signed((reg595[(4'ha):(4'ha)] ?
                  reg1194[(4'hf):(4'h8)] : reg1167[(4'ha):(4'h8)])) >>> ($signed((reg597 ?
                  (7'h43) : reg591)) ~^ ((wire1221 + reg1224) ~^ (~(8'hb1))))));
              reg1227 <= $unsigned((-(!wire1220)));
              reg1228 <= $signed(reg595);
              reg1229 <= (reg603[(2'h2):(1'h1)] >> $signed((^~((8'ha4) >>> $unsigned(wire604)))));
            end
          for (forvar1230 = (1'h0); (forvar1230 < (2'h2)); forvar1230 = (forvar1230 + (1'h1)))
            begin
              reg1231 = (reg670 ?
                  reg1152 : (((&$signed(reg632)) - ($signed(wire1185) ?
                          $unsigned(reg1139) : wire604[(4'hd):(3'h4)])) ?
                      $signed(((wire1185 >>> reg576) <<< $unsigned(reg652))) : reg1104[(4'hc):(2'h3)]));
              reg1232 <= $unsigned($signed(reg618[(3'h6):(1'h0)]));
              reg1233 <= (~(|({{reg1167, reg581, reg1218},
                      (!reg1201),
                      (~&wire1221)} ?
                  wire563 : $signed((reg695 ? reg1182 : (7'h40))))));
              reg1234 <= reg618[(1'h0):(1'h0)];
            end
          for (forvar1235 = (1'h0); (forvar1235 < (2'h3)); forvar1235 = (forvar1235 + (1'h1)))
            begin
              reg1236 = $signed((reg679 ?
                  $unsigned(($signed((8'hbd)) ?
                      reg1233 : (&wire605))) : (~reg1206)));
              reg1237 = (reg638[(2'h3):(2'h2)] ?
                  (!wire1070) : $signed({(reg1191[(1'h1):(1'h1)] && (+reg1077)),
                      $unsigned((~^reg1191))}));
              reg1238 <= $signed(reg1132[(5'h11):(1'h0)]);
              reg1239 = reg695;
              reg1240 <= (|(~^$unsigned($signed(wire565))));
              reg1241 = $signed(wire1220[(3'h5):(2'h2)]);
            end
          reg1242 = ($unsigned($unsigned(wire564[(4'hf):(4'h8)])) != (((reg1163 ?
              reg670[(1'h1):(1'h1)] : (^reg1104)) & ($signed(reg1228) ?
              (+reg1089) : (wire1070 ?
                  reg1132 : reg663))) == reg1209[(2'h3):(1'h1)]));
          if (wire1220[(5'h10):(4'h8)])
            begin
              reg1243 = (7'h55);
              reg1244 <= ({(($unsigned(reg1164) >>> reg636) ?
                      (reg630 ?
                          (reg1201 ?
                              reg674 : reg1182) : {reg1236}) : reg1243)} >> {wire1072});
              reg1245 <= (reg1108 >> reg652);
              reg1246 = reg579;
              reg1247 <= reg679[(2'h2):(1'h1)];
              reg1248 <= $signed(reg572);
              reg1249 <= reg1164;
            end
          else
            begin
              reg1243 = ($unsigned($unsigned(reg588[(1'h0):(1'h0)])) <<< reg667[(2'h3):(1'h0)]);
              reg1244 <= $unsigned((~|$signed((7'h50))));
            end
        end
      if ((reg572[(1'h1):(1'h0)] ?
          $unsigned((reg572[(3'h6):(2'h3)] << reg1155)) : {(((|reg1160) != (reg1224 ?
                  reg576 : reg1155)) > $unsigned($unsigned(reg1171))),
              $unsigned(((reg1246 ? reg668 : reg566) < (reg642 ?
                  reg1186 : reg572))),
              reg573}))
        begin
          for (forvar1250 = (1'h0); (forvar1250 < (2'h3)); forvar1250 = (forvar1250 + (1'h1)))
            begin
              reg1251 = $signed((8'hac));
              reg1252 <= {{(((reg1155 | reg649) ?
                          $unsigned(reg663) : {reg574,
                              reg1137}) != $signed(reg646[(4'hb):(3'h7)]))},
                  (reg1157[(2'h3):(2'h2)] >>> (^reg1147)),
                  $unsigned($signed(reg1147[(3'h5):(2'h2)]))};
              reg1253 <= (^((!(reg663[(3'h6):(2'h3)] >> $signed((7'h47)))) >> (((reg1175 <<< reg1241) ?
                  $unsigned(reg1121) : reg1239[(3'h5):(3'h4)]) >> reg1226[(3'h7):(2'h3)])));
              reg1254 = (~|$unsigned((!((^reg1100) == $signed(reg1232)))));
              reg1255 <= $unsigned($unsigned($unsigned((~^(~(8'ha9))))));
            end
          reg1256 <= (+$unsigned($unsigned($signed((reg1200 ?
              (7'h43) : reg1246)))));
          reg1257 = reg1090[(3'h6):(3'h6)];
          reg1258 = $signed((reg623 ?
              $unsigned((~|$unsigned(reg1231))) : reg1104[(3'h6):(1'h0)]));
          reg1259 = ({reg595[(4'h9):(3'h6)],
                  (($unsigned(reg590) ? wire605[(5'h1c):(4'he)] : reg1245) ?
                      $unsigned($signed((7'h45))) : reg693),
                  (8'hb5)} ?
              ((($unsigned(reg1233) ? reg1188 : reg1171[(2'h2):(1'h0)]) ?
                  (reg1229[(1'h1):(1'h1)] ?
                      reg1251 : reg658) : $unsigned($unsigned(reg690))) << ((-reg1094[(2'h2):(1'h1)]) <= (!(wire1071 ?
                  reg1237 : reg601)))) : $signed($signed(reg576[(3'h6):(3'h5)])));
          reg1260 <= wire1070[(5'h17):(5'h11)];
        end
      else
        begin
          reg1250 = {reg691[(4'h9):(4'h9)]};
          reg1251 = {$unsigned(reg1253)};
          if ($unsigned(($unsigned($signed($unsigned((7'h4b)))) >= (~&$signed($signed(reg1216))))))
            begin
              reg1254 = ((|(((reg667 ?
                          (7'h55) : reg1234) ^~ ((8'hbc) & wire562)) ?
                      reg1160 : reg634)) ?
                  (+(reg1168[(3'h5):(3'h4)] - (8'hbf))) : $signed(((8'ha8) ?
                      reg579[(4'ha):(3'h4)] : reg1224[(5'h15):(3'h5)])));
              reg1255 <= {((reg1252[(4'h9):(3'h6)] & wire564[(5'h11):(4'hf)]) >>> $unsigned({{reg692,
                          reg1131,
                          reg638},
                      (reg631 < wire1070)})),
                  (-(reg685[(4'hf):(1'h0)] > reg621)),
                  reg1186[(4'ha):(1'h1)]};
            end
          else
            begin
              reg1254 = $signed(reg1227);
              reg1257 = $signed(((~^reg630[(5'h16):(5'h12)]) ?
                  $unsigned(reg697[(4'h8):(3'h4)]) : {reg678[(5'h1a):(5'h19)],
                      ($unsigned(reg595) ?
                          {reg1113} : (wire1220 ? reg638 : (8'ha9))),
                      $unsigned({reg1253, reg1147})}));
              reg1260 <= {(&(wire1185[(1'h1):(1'h0)] ?
                      reg1243[(3'h5):(3'h5)] : (&$signed(reg577))))};
              reg1261 = (8'hba);
            end
          if ($signed(reg1199[(3'h4):(1'h0)]))
            begin
              reg1262 <= {(reg1083 ?
                      $signed($unsigned($unsigned(reg1206))) : ((+{wire604,
                              reg1150}) ?
                          ((reg1168 ?
                              (8'hb9) : reg623) - reg597) : $signed($signed(reg570))))};
              reg1263 <= (($signed($signed(forvar1230[(4'he):(3'h7)])) < (~|(reg621 ?
                  (reg1105 == (7'h4b)) : $unsigned(reg1250)))) ^~ ($signed($signed((reg1229 <<< (7'h4b)))) ^ (wire565 + wire1070)));
              reg1264 = ($signed(reg1130) ?
                  reg1132[(5'h12):(2'h2)] : {$unsigned($unsigned(reg1095))});
              reg1265 = $unsigned(forvar1230);
              reg1266 = ({$unsigned($signed((reg1219 ? reg1206 : reg1200))),
                      ((-{reg574, reg1219, reg1118}) ?
                          (~&(&reg685)) : $signed($signed(wire1185)))} ?
                  reg691[(4'ha):(3'h7)] : {$signed((+(|reg1234)))});
              reg1267 = (($signed($unsigned((&reg571))) ?
                  $unsigned($unsigned(reg1264[(3'h7):(3'h6)])) : (&{(reg642 <= reg690)})) & $signed($unsigned($signed(((7'h56) >>> reg1222)))));
              reg1268 <= reg1137;
            end
          else
            begin
              reg1262 <= {(reg1131 ?
                      $signed(reg1219[(4'hb):(2'h2)]) : {reg1251,
                          reg658[(1'h1):(1'h0)],
                          reg1155}),
                  reg674[(1'h1):(1'h1)],
                  reg1213[(3'h5):(2'h3)]};
              reg1263 <= (wire564 ?
                  $unsigned(($signed($unsigned(reg1167)) ?
                      ($signed(reg1218) - $signed(reg1105)) : $unsigned(reg1231[(3'h7):(3'h5)]))) : reg576[(3'h5):(1'h0)]);
              reg1264 = {(-$unsigned($unsigned({reg633}))),
                  ($signed(reg1121[(4'ha):(1'h0)]) ?
                      $unsigned($unsigned((reg680 == (8'hb6)))) : (wire1070[(2'h3):(2'h3)] ?
                          reg1163[(3'h5):(2'h2)] : (!$signed((8'haa)))))};
              reg1265 = $signed(reg601[(1'h0):(1'h0)]);
              reg1266 = (8'ha8);
            end
        end
      reg1269 <= $signed({reg632[(1'h1):(1'h1)],
          reg1106[(3'h4):(1'h1)],
          {((reg1224 && (8'ha3)) ? (~&reg670) : reg566[(4'hb):(3'h7)]),
              $signed($signed(reg1140))}});
    end
  assign wire1270 = (~|(((reg597[(3'h4):(3'h4)] >>> reg1219[(4'h9):(1'h0)]) ?
                        (~{wire563}) : reg1093[(2'h2):(1'h0)]) != $signed((|(reg637 ^~ reg1217)))));
  always
    @(posedge clk) begin
      if (reg1252)
        begin
          for (forvar1271 = (1'h0); (forvar1271 < (3'h5)); forvar1271 = (forvar1271 + (1'h1)))
            begin
              reg1272 <= (~&($signed((reg591 ?
                      {reg1086, (8'ha4), (8'h9e)} : $unsigned(reg1263))) ?
                  ({(reg601 ? reg568 : reg1269), (reg1219 >>> reg579)} ?
                      reg1089[(4'hc):(4'ha)] : (^~$signed(reg644))) : ((-(7'h4f)) ?
                      $signed($signed(reg1173)) : ($unsigned(reg1228) + $signed((7'h53))))));
              reg1273 = reg631[(3'h4):(2'h3)];
              reg1274 <= reg1113[(5'h10):(3'h5)];
              reg1275 <= reg1132[(5'h1b):(5'h11)];
            end
          if ((~|($signed($signed((reg603 | reg1210))) && (&reg603))))
            begin
              reg1276 = $signed($unsigned(((reg603[(2'h3):(1'h0)] && (~&reg1098)) ?
                  forvar1271 : ($signed(reg679) * (!reg601)))));
              reg1277 = (reg1155[(3'h4):(2'h2)] ?
                  $unsigned(($unsigned(reg1155[(4'h8):(2'h2)]) ?
                      (reg1168[(5'h10):(5'h10)] & reg697) : $signed((!(7'h42))))) : (8'ha8));
              reg1278 = $signed(reg1100);
            end
          else
            begin
              reg1276 = (reg597 ?
                  $signed(reg677) : (-(~(reg668[(5'h11):(3'h6)] < {reg625}))));
              reg1277 = {((8'ha3) >> {$unsigned(reg643[(4'he):(3'h7)])}),
                  ($signed(((reg1168 < (8'hbf)) ?
                      $unsigned(reg697) : (-(8'hb7)))) >= reg1089),
                  wire1270[(1'h0):(1'h0)]};
              reg1279 <= {(~^$signed(reg601[(4'h9):(4'h8)])),
                  (-$signed(reg1094))};
            end
        end
      else
        begin
          for (forvar1271 = (1'h0); (forvar1271 < (2'h3)); forvar1271 = (forvar1271 + (1'h1)))
            begin
              reg1273 = (-reg1253);
              reg1274 <= ($signed(((^reg641[(1'h0):(1'h0)]) ?
                  reg690[(3'h6):(3'h4)] : ((wire565 != (7'h4c)) > {reg653,
                      reg1094,
                      (8'ha6)}))) ^ ($signed($unsigned({reg1118,
                  (7'h53)})) * (&({reg1269} <= $signed((8'had))))));
              reg1275 <= ($signed({(~reg1089),
                  reg1194[(5'h1b):(5'h1b)],
                  (-$signed((7'h53)))}) ^~ $signed((((^reg1227) - $unsigned(wire1220)) >>> {(7'h47)})));
              reg1276 = reg1157[(5'h19):(4'hc)];
              reg1277 = $signed((($unsigned(reg623) - {(reg576 ?
                          reg1224 : reg616),
                      (reg1089 ^~ reg616),
                      (reg566 >> reg1248)}) ?
                  reg1273 : reg1106));
            end
          reg1279 <= {$signed(reg1077),
              reg1157[(5'h13):(5'h11)],
              $signed((!$unsigned($signed(reg1098))))};
          reg1280 <= reg1094[(4'hd):(2'h3)];
          if ($signed($signed(reg1216)))
            begin
              reg1281 = ((^$unsigned($unsigned((~&wire1073)))) > reg693[(3'h4):(2'h2)]);
              reg1282 <= reg1263;
              reg1283 <= reg1105;
            end
          else
            begin
              reg1282 <= $unsigned($unsigned({(^~reg1281),
                  {(^reg574)},
                  $signed(reg1240)}));
              reg1283 <= reg678;
              reg1284 <= $unsigned(($signed(reg1157[(4'hc):(4'ha)]) ?
                  $signed($signed((~^(8'h9d)))) : $unsigned(((reg1276 ?
                      (8'had) : reg567) != (reg1147 >>> reg1248)))));
            end
          for (forvar1285 = (1'h0); (forvar1285 < (3'h4)); forvar1285 = (forvar1285 + (1'h1)))
            begin
              reg1286 = (reg657[(3'h7):(1'h1)] ?
                  (~&($unsigned((reg1173 ?
                      reg1281 : reg1280)) ^ ((~^reg637) ~^ ((8'hb9) ~^ reg1150)))) : ((wire1221[(5'h1d):(4'hf)] <<< (^$unsigned(reg663))) == (7'h53)));
              reg1287 <= $unsigned((~|$unsigned(reg1163[(5'h11):(2'h2)])));
              reg1288 = reg1139[(1'h1):(1'h1)];
              reg1289 <= ({(|{(reg1108 ? (8'hae) : reg1286)})} ?
                  {$unsigned(reg697),
                      reg1248[(5'h11):(3'h6)]} : $signed($signed((reg566[(3'h6):(2'h2)] ^ (^(8'ha3))))));
              reg1290 = (((reg630 ?
                      ((-wire565) < (7'h53)) : $signed(reg1233)) ~^ ((-(reg1090 ?
                      (7'h47) : reg1287)) * $signed($unsigned(reg674)))) ?
                  $signed((&(+{reg1218, reg573, (8'hb2)}))) : reg1284);
              reg1291 = ((7'h51) ?
                  $signed(((|reg678) ?
                      reg1083 : (&$unsigned(wire615)))) : ($signed((~&$signed(reg693))) ?
                      $signed(reg1118) : reg642));
              reg1292 <= reg643;
            end
          for (forvar1293 = (1'h0); (forvar1293 < (1'h0)); forvar1293 = (forvar1293 + (1'h1)))
            begin
              reg1294 = ($unsigned(reg696[(3'h4):(2'h3)]) ?
                  $unsigned((~(reg668 ?
                      (^~reg1160) : $signed(reg1290)))) : (((reg1199[(2'h3):(1'h0)] || $signed(reg1286)) ?
                      $signed(reg1092) : reg1130) - $signed($signed($unsigned(reg1104)))));
              reg1295 = ($unsigned(($signed((|reg1152)) << reg1272[(2'h2):(2'h2)])) ?
                  ((!(^~reg693)) == {(reg1213[(1'h0):(1'h0)] ?
                          (+(7'h4d)) : (~^reg1173)),
                      reg677[(4'he):(3'h6)]}) : $unsigned((((reg1155 && (7'h50)) ?
                          $unsigned(reg1278) : reg576) ?
                      ({(7'h57), reg1284} == (reg1152 ?
                          reg1216 : reg1121)) : reg1137)));
              reg1296 = {(^~$unsigned($unsigned((reg1175 << reg1160)))),
                  $signed((reg621 ^ wire1270)),
                  ((~reg1175[(1'h1):(1'h1)]) - (reg603 ?
                      reg1269 : (wire1221 ?
                          $unsigned(reg693) : $unsigned(reg1106))))};
            end
          reg1297 = $unsigned(reg1295);
        end
      if (($signed($signed($unsigned((reg1233 >= reg1240)))) ?
          $signed($signed((reg1229 <<< $signed(reg1160)))) : $signed((!{reg577,
              reg1272[(3'h4):(3'h4)],
              reg1229}))))
        begin
          if ($unsigned((!((reg1181 != reg692[(5'h10):(5'h10)]) ?
              {(reg591 ?
                      reg597 : (8'h9d))} : $unsigned((reg1200 >= reg1121))))))
            begin
              reg1298 <= ((-reg1262) <= $unsigned($unsigned(reg1276[(5'h11):(4'hd)])));
              reg1299 = ((8'hb5) >= reg636[(5'h14):(4'hc)]);
              reg1300 <= $unsigned($unsigned(reg1083[(4'hf):(4'ha)]));
              reg1301 <= $unsigned($unsigned($unsigned((reg1232[(3'h7):(2'h2)] <= reg638))));
              reg1302 = $signed(reg1232[(4'h8):(2'h2)]);
              reg1303 = reg1157[(2'h2):(1'h0)];
              reg1304 = (reg1263 != $unsigned($signed($unsigned((reg650 ?
                  reg1256 : reg669)))));
            end
          else
            begin
              reg1298 <= (($unsigned({reg690, (reg1194 ? reg1090 : reg1206)}) ?
                      (({reg1277,
                          wire1185} == (reg1280 <<< reg1121)) > (&reg1291[(1'h1):(1'h1)])) : $signed($signed((^~reg644)))) ?
                  $unsigned(reg1245) : reg568[(2'h2):(1'h1)]);
              reg1300 <= ((^~(^$signed((~|wire565)))) < (^(~((wire565 <<< reg632) ?
                  (^~reg1213) : reg1200[(4'hb):(4'ha)]))));
              reg1302 = {((reg1276 ?
                          wire1070 : {reg697[(5'h10):(3'h7)], reg574}) ?
                      (({wire565} ~^ reg1276) <<< $signed(reg595)) : reg1302),
                  reg1233};
              reg1303 = reg1273[(4'hb):(4'ha)];
            end
          reg1305 = ($signed($signed(($signed(reg658) ?
                  (7'h44) : $signed((7'h56))))) ?
              (&(^$signed({reg1210}))) : reg1262[(3'h7):(1'h1)]);
          reg1306 <= reg1255;
          reg1307 = ((((~^wire1110[(3'h5):(3'h5)]) < (+$unsigned(reg1232))) ?
                  ($unsigned(reg616[(5'h1a):(2'h2)]) << {(reg1218 ?
                          wire564 : (8'h9f)),
                      (!reg1232)}) : reg1098[(4'h8):(4'h8)]) ?
              reg691 : (&(reg1156[(4'h8):(3'h6)] ?
                  $unsigned(reg571[(1'h1):(1'h1)]) : {(+(8'hb0))})));
          reg1308 = $unsigned(reg1171[(3'h4):(2'h3)]);
          if ($signed(reg653))
            begin
              reg1309 <= reg579;
              reg1310 <= $unsigned({$unsigned($signed(reg1248[(5'h12):(4'ha)])),
                  (~^({reg570, reg1137, reg652} ?
                      (reg668 ? reg1102 : reg566) : (-(8'hb3)))),
                  wire1270[(1'h0):(1'h0)]});
              reg1311 = ($signed($unsigned(((!(7'h56)) ?
                      (reg1094 ? reg1232 : reg1121) : $signed(reg1093)))) ?
                  reg1089[(3'h6):(1'h0)] : $unsigned(reg667[(4'hb):(3'h6)]));
              reg1312 = (reg1216[(5'h1d):(5'h18)] ?
                  ($unsigned($signed((reg1228 ?
                      reg692 : reg1299))) | {reg1106}) : reg579);
              reg1313 = $signed($unsigned(($unsigned((reg634 ?
                  reg677 : (8'hb8))) | ((!(8'ha0)) >>> $signed(reg1209)))));
              reg1314 <= $signed((+$signed((^~$unsigned(reg668)))));
              reg1315 <= reg1095[(3'h6):(2'h2)];
            end
          else
            begin
              reg1309 <= $unsigned($unsigned(($unsigned((-reg669)) >> (reg1228 & (~^reg1304)))));
              reg1310 <= reg1194;
              reg1314 <= reg1118;
              reg1316 = reg697;
              reg1317 = $signed(reg1213[(4'h8):(4'h8)]);
              reg1318 = ((reg1315[(5'h17):(5'h16)] > reg653[(3'h4):(2'h3)]) ?
                  (7'h52) : (~&$unsigned({$signed(reg675)})));
            end
        end
      else
        begin
          if ($unsigned($signed(reg1200)))
            begin
              reg1299 = ({(reg1289[(1'h0):(1'h0)] ?
                          reg1245 : $unsigned(reg637[(4'hb):(1'h0)]))} ?
                  forvar1293 : $signed(($unsigned($signed(reg668)) ^~ ((reg1089 ?
                          reg695 : (8'ha8)) ?
                      $unsigned(reg670) : reg1308))));
            end
          else
            begin
              reg1299 = (~|($signed(reg1252[(5'h10):(2'h3)]) || $unsigned($unsigned((reg1083 + wire1185)))));
            end
          reg1300 <= {reg595, reg1294, $unsigned(wire1185)};
          if (((({$unsigned(wire1220),
              reg1275[(1'h0):(1'h0)],
              (^reg1105)} > $signed((!reg618))) * $unsigned(((reg1226 & reg1150) ?
              reg568 : (8'hbc)))) ~^ ((-reg1160) <= reg1245)))
            begin
              reg1301 <= ($unsigned((($unsigned(wire1220) || reg680) ?
                      $signed($signed(reg572)) : $signed(reg641[(4'ha):(1'h0)]))) ?
                  (reg678 ~^ reg1182) : wire1220);
              reg1302 = reg697;
              reg1303 = (^((((reg1113 != reg649) ?
                      $unsigned(reg1160) : $unsigned(reg1150)) ^~ $signed((reg1102 << reg603))) ?
                  $signed({$unsigned((7'h48)),
                      reg1141,
                      reg1286[(5'h19):(4'ha)]}) : $signed((8'hb0))));
              reg1306 <= (reg567[(4'h9):(4'h9)] ?
                  {{{reg1290[(3'h7):(3'h5)], reg1255[(4'hc):(2'h3)]}},
                      $signed(reg597),
                      reg667[(1'h1):(1'h0)]} : (+(+reg1106[(3'h4):(3'h4)])));
              reg1309 <= (~|{{reg1182}, $unsigned((-reg675[(3'h5):(2'h2)]))});
            end
          else
            begin
              reg1302 = (+$signed((reg663[(1'h1):(1'h1)] ?
                  ((reg1126 ? reg1292 : reg1139) ?
                      (wire1070 ?
                          reg1186 : reg693) : $signed(reg1219)) : (wire1221 ?
                      {reg1318, reg577, reg1226} : $unsigned(reg1316)))));
              reg1306 <= ((($unsigned({reg679}) ?
                          reg568 : $signed($unsigned(reg1175))) ?
                      $unsigned($signed({reg1227})) : (|{{reg1253,
                              reg1201,
                              reg1260}})) ?
                  $signed({$unsigned((reg1217 ? reg653 : (8'hae))),
                      $signed(reg1227)}) : (~|(|$unsigned((reg603 <= reg603)))));
              reg1309 <= reg1274[(5'h19):(3'h7)];
              reg1310 <= reg1314;
            end
          for (forvar1311 = (1'h0); (forvar1311 < (1'h1)); forvar1311 = (forvar1311 + (1'h1)))
            begin
              reg1312 = (&((reg1113[(1'h1):(1'h1)] & ({wire1220, reg1140} ?
                  $signed(reg1274) : $signed(reg1218))) + (reg692 ?
                  (^~{(8'hb6), reg572, wire564}) : reg632)));
              reg1314 <= (reg658[(2'h2):(2'h2)] ?
                  (({(reg1141 < reg591),
                      $signed((8'h9e))} >> ($unsigned(reg1240) && (reg572 >= wire1270))) + ($unsigned((reg1132 >= wire562)) - $unsigned($signed(reg636)))) : $unsigned(reg680[(3'h7):(1'h1)]));
              reg1316 = {({reg1188,
                          (^reg1277),
                          $signed(reg1097[(3'h5):(2'h2)])} ?
                      reg1217 : (~|reg1229)),
                  (((&(~|reg653)) ?
                      $unsigned(reg638) : (|(reg638 << reg1217))) <<< $signed(wire1221[(3'h5):(3'h5)])),
                  (7'h4b)};
              reg1319 <= $signed((reg697 < (8'ha1)));
              reg1320 = (^(reg669 ?
                  $signed((7'h51)) : (~&$signed((~^reg1226)))));
              reg1321 = (~&((~|reg1298[(3'h7):(2'h3)]) ?
                  {((+reg1268) < (8'hb3)),
                      $signed(reg1273[(4'ha):(3'h5)]),
                      reg1295[(2'h3):(2'h2)]} : $unsigned(reg1181)));
            end
          reg1322 <= (&((reg1224[(5'h18):(3'h5)] ?
                  reg1320[(4'hc):(3'h6)] : ((~&reg1094) & (reg1289 - reg625))) ?
              ((reg1098[(1'h1):(1'h0)] << $unsigned(reg1291)) ?
                  (~|$signed((8'hbd))) : {(reg592 ?
                          forvar1285 : reg579)}) : ($signed({wire1071}) ?
                  (!$unsigned(reg1106)) : reg628[(5'h18):(3'h7)])));
        end
      if ($signed($signed($unsigned((|$unsigned(reg1281))))))
        begin
          reg1323 = ($unsigned($unsigned((((8'ha2) ?
                  reg1263 : reg641) == (+reg1157)))) ?
              ($unsigned($unsigned(reg1141)) ?
                  reg1094[(2'h3):(2'h3)] : (reg693 && $unsigned(((7'h44) ?
                      reg1284 : reg1167)))) : (((^(reg1256 ?
                      reg1093 : reg597)) ?
                  reg1314[(5'h15):(5'h14)] : reg1255[(4'he):(1'h0)]) >> reg1299[(5'h16):(5'h12)]));
        end
      else
        begin
          for (forvar1323 = (1'h0); (forvar1323 < (2'h2)); forvar1323 = (forvar1323 + (1'h1)))
            begin
              reg1324 <= reg566;
              reg1325 = reg597;
              reg1326 <= reg1318[(2'h2):(1'h0)];
              reg1327 = ((~&{$unsigned($signed(reg1132)),
                  $unsigned((reg1300 ?
                      wire563 : (8'h9d)))}) <= reg667[(2'h3):(2'h2)]);
              reg1328 <= (reg1232[(1'h0):(1'h0)] >>> $signed({reg1200[(1'h1):(1'h1)],
                  (reg1232 > reg692[(4'h9):(4'h9)]),
                  (8'hba)}));
              reg1329 = (~((~&$unsigned($signed(reg1290))) + (!reg663[(3'h5):(2'h2)])));
            end
          reg1330 = reg1275[(2'h2):(1'h1)];
          if ($unsigned($signed($unsigned(reg670[(2'h3):(1'h0)]))))
            begin
              reg1331 = ({reg570[(3'h6):(2'h2)],
                  reg1092[(5'h10):(4'h9)]} == (^reg582[(3'h6):(3'h4)]));
              reg1332 <= $unsigned($signed((((~&reg650) ?
                  $signed(reg1086) : reg1278[(1'h0):(1'h0)]) >= (reg612 == {(8'hb1)}))));
            end
          else
            begin
              reg1331 = $unsigned((8'ha6));
            end
          reg1333 <= reg1194;
          for (forvar1334 = (1'h0); (forvar1334 < (1'h1)); forvar1334 = (forvar1334 + (1'h1)))
            begin
              reg1335 <= reg1249[(5'h12):(4'he)];
              reg1336 = (~reg1206);
              reg1337 <= ((&$signed(((reg643 ? reg1092 : reg1095) ?
                  reg1298[(3'h5):(3'h5)] : reg1280))) >>> {$signed($unsigned((reg1227 >= reg591))),
                  reg566[(2'h3):(2'h2)]});
              reg1338 <= (7'h4a);
              reg1339 <= {($signed((^reg1305[(1'h1):(1'h1)])) ?
                      (-((!reg1199) <= (-reg1216))) : (~&((+reg582) ?
                          reg1132[(5'h14):(2'h2)] : $signed(reg1288))))};
            end
        end
      if (wire604[(5'h12):(4'hc)])
        begin
          if (wire1071[(2'h3):(2'h2)])
            begin
              reg1340 <= reg1233;
              reg1341 = reg1191;
              reg1342 <= $unsigned($unsigned($signed($signed($signed(reg1206)))));
              reg1343 <= (!wire604);
              reg1344 = (($unsigned($unsigned($signed(reg1244))) ?
                      (^((reg1130 <= reg667) | (reg1290 <= (8'hbb)))) : (((reg1291 != reg1325) & $unsigned(reg652)) ?
                          reg1326 : $signed($unsigned(reg595)))) ?
                  (reg1086 ?
                      ($unsigned($unsigned(reg612)) ?
                          reg1163[(4'ha):(2'h2)] : {(&reg1278)}) : $signed(reg653)) : (-(~reg1194)));
              reg1345 <= reg601[(5'h13):(5'h10)];
              reg1346 = reg601;
            end
          else
            begin
              reg1341 = reg669[(4'hf):(4'ha)];
              reg1344 = $unsigned($signed(reg1291[(3'h7):(1'h1)]));
              reg1346 = (reg568 ?
                  (^(^~$signed(reg1186))) : (reg1276 ?
                      $signed((((8'hbc) ? reg1186 : reg1171) ?
                          (reg1287 || (8'hb2)) : $unsigned(reg603))) : ((^reg1199[(1'h0):(1'h0)]) * reg1303[(2'h2):(1'h0)])));
              reg1347 <= (-$unsigned(reg1141));
            end
        end
      else
        begin
          reg1340 <= reg1191[(2'h3):(2'h3)];
        end
      for (forvar1348 = (1'h0); (forvar1348 < (1'h1)); forvar1348 = (forvar1348 + (1'h1)))
        begin
          reg1349 = ($signed(((-(reg1228 <<< reg1280)) | reg568)) && reg644[(5'h11):(4'ha)]);
          if ((reg1233[(2'h2):(1'h1)] >> reg1188[(3'h4):(2'h3)]))
            begin
              reg1350 = $signed((reg1118 ?
                  ((wire1270 || (reg1186 ?
                      reg1274 : reg591)) << wire1221[(5'h1b):(1'h1)]) : $unsigned(((~^(8'h9f)) | reg1218[(1'h1):(1'h0)]))));
              reg1351 <= {(({((7'h54) + reg1137),
                      $unsigned(reg1336)} && reg612) << reg1295[(2'h2):(1'h0)])};
              reg1352 <= $unsigned(reg570);
              reg1353 <= $unsigned((7'h44));
            end
          else
            begin
              reg1350 = ($signed(((+reg1350) ?
                      $signed({reg690, reg1238}) : reg1253)) ?
                  $unsigned(wire1070[(3'h6):(1'h1)]) : ($unsigned(reg1104[(3'h5):(3'h5)]) | wire562[(3'h6):(2'h3)]));
              reg1354 = (reg1338[(2'h3):(2'h2)] > (({reg1328[(2'h2):(1'h1)],
                      $unsigned(reg1156)} ?
                  {$unsigned(reg1171),
                      $signed(reg643)} : reg566[(2'h3):(1'h0)]) > reg1227[(4'h8):(3'h4)]));
              reg1355 <= reg1132[(4'hb):(3'h6)];
              reg1356 <= reg1152[(2'h3):(1'h0)];
            end
        end
    end
  assign wire1357 = reg1188;
  assign wire1358 = $unsigned(((|$signed(reg1081)) >>> $unsigned({reg1139[(2'h3):(2'h3)],
                        (reg652 || reg592),
                        $unsigned((8'hb0))})));
  assign wire1359 = $unsigned({wire605[(3'h4):(1'h1)],
                        $signed(reg1173[(3'h7):(3'h5)])});
  always
    @(posedge clk) begin
      reg1360 = $unsigned((((reg588[(1'h1):(1'h1)] + $unsigned((8'hb6))) - (reg1090[(4'h9):(2'h2)] == (reg582 <<< reg1089))) ?
          (($unsigned(wire1359) <<< reg1210) >>> (&(7'h4b))) : $unsigned(reg1234[(1'h1):(1'h1)])));
    end
  assign wire1361 = reg1098[(4'h9):(2'h2)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module702
#(parameter param1067 = (^~(&((^(+(7'h43))) << (((8'hb9) || (7'h4b)) == (+(8'ha5)))))))
(y, clk, wire706, wire705, wire704, wire703);
  output wire [(32'h1794):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire706;
  input wire signed [(4'hd):(1'h0)] wire705;
  input wire [(4'hb):(1'h0)] wire704;
  input wire signed [(4'he):(1'h0)] wire703;
  wire signed [(4'hc):(1'h0)] wire1007;
  wire signed [(4'hc):(1'h0)] wire1006;
  wire [(3'h4):(1'h0)] wire1005;
  wire [(4'hb):(1'h0)] wire825;
  wire signed [(3'h6):(1'h0)] wire709;
  wire [(2'h3):(1'h0)] wire708;
  wire [(5'h10):(1'h0)] wire707;
  reg signed [(5'h11):(1'h0)] reg1060 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1056 = (1'h0);
  reg [(4'h9):(1'h0)] reg1055 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1053 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1048 = (1'h0);
  reg [(2'h2):(1'h0)] reg1044 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1043 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1042 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1039 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1038 = (1'h0);
  reg [(5'h14):(1'h0)] reg1037 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1035 = (1'h0);
  reg [(4'he):(1'h0)] reg1034 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1033 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1031 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1026 = (1'h0);
  reg [(4'hf):(1'h0)] reg1025 = (1'h0);
  reg [(3'h7):(1'h0)] reg1024 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1023 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1022 = (1'h0);
  reg [(3'h7):(1'h0)] reg1020 = (1'h0);
  reg [(5'h17):(1'h0)] reg1018 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1015 = (1'h0);
  reg [(3'h4):(1'h0)] reg1013 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1009 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1004 = (1'h0);
  reg [(4'hf):(1'h0)] reg1003 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1000 = (1'h0);
  reg [(5'h10):(1'h0)] reg998 = (1'h0);
  reg [(5'h10):(1'h0)] reg994 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg985 = (1'h0);
  reg [(5'h1e):(1'h0)] reg984 = (1'h0);
  reg [(3'h5):(1'h0)] reg983 = (1'h0);
  reg [(5'h17):(1'h0)] reg982 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg979 = (1'h0);
  reg [(5'h18):(1'h0)] reg978 = (1'h0);
  reg [(5'h1e):(1'h0)] reg976 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg974 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg972 = (1'h0);
  reg [(5'h1f):(1'h0)] reg969 = (1'h0);
  reg [(5'h16):(1'h0)] reg965 = (1'h0);
  reg [(5'h14):(1'h0)] reg962 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg961 = (1'h0);
  reg [(2'h2):(1'h0)] reg956 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg954 = (1'h0);
  reg [(3'h7):(1'h0)] reg950 = (1'h0);
  reg [(3'h7):(1'h0)] reg948 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg943 = (1'h0);
  reg [(2'h2):(1'h0)] reg941 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg938 = (1'h0);
  reg [(5'h1c):(1'h0)] reg928 = (1'h0);
  reg [(5'h14):(1'h0)] reg934 = (1'h0);
  reg [(3'h4):(1'h0)] reg933 = (1'h0);
  reg [(3'h7):(1'h0)] reg932 = (1'h0);
  reg [(2'h3):(1'h0)] reg930 = (1'h0);
  reg [(4'hf):(1'h0)] reg929 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg926 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg925 = (1'h0);
  reg [(2'h3):(1'h0)] reg923 = (1'h0);
  reg [(4'h8):(1'h0)] reg919 = (1'h0);
  reg [(4'he):(1'h0)] reg913 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg911 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg909 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg908 = (1'h0);
  reg [(4'h8):(1'h0)] reg907 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg905 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg901 = (1'h0);
  reg [(5'h12):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg898 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg894 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg892 = (1'h0);
  reg [(4'h8):(1'h0)] reg891 = (1'h0);
  reg [(5'h1e):(1'h0)] reg887 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg886 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg885 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg881 = (1'h0);
  reg [(4'hb):(1'h0)] reg880 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg878 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg877 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg875 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg874 = (1'h0);
  reg [(3'h5):(1'h0)] reg872 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg870 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg869 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg868 = (1'h0);
  reg [(2'h2):(1'h0)] reg862 = (1'h0);
  reg [(5'h1f):(1'h0)] reg863 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg859 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg849 = (1'h0);
  reg [(5'h1c):(1'h0)] reg855 = (1'h0);
  reg [(2'h3):(1'h0)] reg854 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg853 = (1'h0);
  reg signed [(4'he):(1'h0)] reg846 = (1'h0);
  reg signed [(4'he):(1'h0)] reg842 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg841 = (1'h0);
  reg [(5'h14):(1'h0)] reg840 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg838 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg836 = (1'h0);
  reg [(5'h1a):(1'h0)] reg833 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg832 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg831 = (1'h0);
  reg [(5'h10):(1'h0)] reg827 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg824 = (1'h0);
  reg [(5'h15):(1'h0)] reg821 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg820 = (1'h0);
  reg [(4'ha):(1'h0)] reg819 = (1'h0);
  reg [(5'h14):(1'h0)] reg815 = (1'h0);
  reg [(4'hf):(1'h0)] reg814 = (1'h0);
  reg [(5'h1b):(1'h0)] reg810 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg809 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg808 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg807 = (1'h0);
  reg [(3'h6):(1'h0)] reg790 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg802 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg801 = (1'h0);
  reg [(2'h3):(1'h0)] reg800 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg799 = (1'h0);
  reg [(5'h17):(1'h0)] reg797 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg795 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg791 = (1'h0);
  reg [(5'h1a):(1'h0)] reg784 = (1'h0);
  reg [(5'h1f):(1'h0)] reg779 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg778 = (1'h0);
  reg [(5'h19):(1'h0)] reg777 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg776 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg775 = (1'h0);
  reg [(5'h1a):(1'h0)] reg773 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg770 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg769 = (1'h0);
  reg [(5'h11):(1'h0)] reg768 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg766 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg761 = (1'h0);
  reg [(2'h2):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg756 = (1'h0);
  reg [(5'h1c):(1'h0)] reg755 = (1'h0);
  reg [(5'h11):(1'h0)] reg754 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg752 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg750 = (1'h0);
  reg [(4'hd):(1'h0)] reg749 = (1'h0);
  reg [(4'ha):(1'h0)] reg747 = (1'h0);
  reg [(2'h2):(1'h0)] reg746 = (1'h0);
  reg [(4'he):(1'h0)] reg742 = (1'h0);
  reg [(5'h1a):(1'h0)] reg741 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg740 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg738 = (1'h0);
  reg [(5'h1d):(1'h0)] reg737 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg733 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg732 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg726 = (1'h0);
  reg [(2'h3):(1'h0)] reg724 = (1'h0);
  reg [(5'h1d):(1'h0)] reg720 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg715 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg714 = (1'h0);
  reg [(4'hd):(1'h0)] reg713 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1066 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1065 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1064 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1063 = (1'h0);
  reg [(4'hc):(1'h0)] reg1062 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1061 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1059 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1058 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1057 = (1'h0);
  reg [(2'h2):(1'h0)] reg1054 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1052 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1051 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1049 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1047 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1046 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1045 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1041 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar1040 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1036 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1032 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1030 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1029 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1028 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1027 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1021 = (1'h0);
  reg [(5'h14):(1'h0)] reg1019 = (1'h0);
  reg [(4'he):(1'h0)] reg1017 = (1'h0);
  reg [(2'h2):(1'h0)] reg1016 = (1'h0);
  reg [(4'he):(1'h0)] reg1014 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1012 = (1'h0);
  reg [(3'h6):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1010 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1008 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1002 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1001 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg999 = (1'h0);
  reg [(4'h9):(1'h0)] reg997 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg996 = (1'h0);
  reg [(5'h12):(1'h0)] reg995 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg993 = (1'h0);
  reg [(2'h3):(1'h0)] forvar992 = (1'h0);
  reg [(4'hf):(1'h0)] reg991 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg990 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg989 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar988 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg987 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg986 = (1'h0);
  reg [(4'hc):(1'h0)] reg981 = (1'h0);
  reg [(3'h6):(1'h0)] reg980 = (1'h0);
  reg [(5'h16):(1'h0)] reg977 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar975 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg973 = (1'h0);
  reg [(3'h4):(1'h0)] reg971 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg970 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg968 = (1'h0);
  reg [(5'h18):(1'h0)] forvar967 = (1'h0);
  reg [(2'h2):(1'h0)] reg966 = (1'h0);
  reg [(5'h13):(1'h0)] reg964 = (1'h0);
  reg [(4'hf):(1'h0)] reg963 = (1'h0);
  reg [(4'hb):(1'h0)] reg960 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg959 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg958 = (1'h0);
  reg [(4'hb):(1'h0)] forvar957 = (1'h0);
  reg [(5'h15):(1'h0)] reg955 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg953 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar952 = (1'h0);
  reg [(5'h16):(1'h0)] reg951 = (1'h0);
  reg [(3'h7):(1'h0)] reg949 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg947 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg946 = (1'h0);
  reg [(4'ha):(1'h0)] reg945 = (1'h0);
  reg [(5'h16):(1'h0)] forvar944 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg942 = (1'h0);
  reg [(4'he):(1'h0)] reg940 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg939 = (1'h0);
  reg [(5'h11):(1'h0)] reg937 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar936 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg935 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg931 = (1'h0);
  reg [(3'h4):(1'h0)] forvar928 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg927 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg924 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg922 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar921 = (1'h0);
  reg [(2'h2):(1'h0)] reg920 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg918 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg917 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg916 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg915 = (1'h0);
  reg [(2'h2):(1'h0)] reg914 = (1'h0);
  reg [(3'h4):(1'h0)] reg912 = (1'h0);
  reg [(4'he):(1'h0)] reg910 = (1'h0);
  reg [(5'h14):(1'h0)] forvar895 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar910 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg906 = (1'h0);
  reg [(5'h12):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg902 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg899 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg897 = (1'h0);
  reg [(5'h12):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg893 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg890 = (1'h0);
  reg [(5'h1f):(1'h0)] reg889 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg888 = (1'h0);
  reg [(5'h12):(1'h0)] reg884 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg883 = (1'h0);
  reg [(5'h12):(1'h0)] reg882 = (1'h0);
  reg [(5'h16):(1'h0)] forvar879 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg876 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg873 = (1'h0);
  reg [(5'h1b):(1'h0)] reg871 = (1'h0);
  reg [(5'h19):(1'h0)] forvar867 = (1'h0);
  reg [(5'h15):(1'h0)] reg866 = (1'h0);
  reg [(4'he):(1'h0)] forvar858 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg857 = (1'h0);
  reg [(5'h16):(1'h0)] reg865 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg864 = (1'h0);
  reg [(5'h19):(1'h0)] forvar862 = (1'h0);
  reg [(5'h1b):(1'h0)] reg861 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg860 = (1'h0);
  reg [(3'h5):(1'h0)] reg858 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar857 = (1'h0);
  reg [(5'h14):(1'h0)] reg856 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg852 = (1'h0);
  reg [(5'h15):(1'h0)] reg851 = (1'h0);
  reg [(5'h15):(1'h0)] reg850 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar849 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg848 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg847 = (1'h0);
  reg [(5'h17):(1'h0)] reg845 = (1'h0);
  reg [(5'h18):(1'h0)] reg844 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg843 = (1'h0);
  reg [(5'h14):(1'h0)] reg839 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg837 = (1'h0);
  reg [(4'h8):(1'h0)] reg835 = (1'h0);
  reg [(5'h19):(1'h0)] forvar834 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg830 = (1'h0);
  reg [(4'ha):(1'h0)] forvar829 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg828 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar826 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg823 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg822 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg818 = (1'h0);
  reg [(5'h1c):(1'h0)] reg817 = (1'h0);
  reg [(5'h1a):(1'h0)] reg816 = (1'h0);
  reg [(5'h14):(1'h0)] reg813 = (1'h0);
  reg [(4'he):(1'h0)] reg812 = (1'h0);
  reg [(4'hf):(1'h0)] reg811 = (1'h0);
  reg [(4'h9):(1'h0)] reg806 = (1'h0);
  reg [(5'h11):(1'h0)] reg805 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg804 = (1'h0);
  reg [(4'ha):(1'h0)] reg803 = (1'h0);
  reg [(5'h10):(1'h0)] reg798 = (1'h0);
  reg [(5'h10):(1'h0)] reg796 = (1'h0);
  reg [(5'h1a):(1'h0)] reg794 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg793 = (1'h0);
  reg [(4'hd):(1'h0)] reg792 = (1'h0);
  reg [(3'h5):(1'h0)] forvar790 = (1'h0);
  reg [(5'h1a):(1'h0)] reg789 = (1'h0);
  reg [(3'h5):(1'h0)] reg788 = (1'h0);
  reg [(5'h10):(1'h0)] reg787 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar786 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg785 = (1'h0);
  reg [(4'h9):(1'h0)] reg783 = (1'h0);
  reg [(5'h12):(1'h0)] reg782 = (1'h0);
  reg [(4'hf):(1'h0)] forvar781 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg765 = (1'h0);
  reg [(5'h10):(1'h0)] forvar758 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar741 = (1'h0);
  reg [(5'h1d):(1'h0)] reg780 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg774 = (1'h0);
  reg [(5'h1e):(1'h0)] reg772 = (1'h0);
  reg [(4'h8):(1'h0)] reg771 = (1'h0);
  reg [(5'h11):(1'h0)] reg767 = (1'h0);
  reg [(5'h13):(1'h0)] forvar765 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg764 = (1'h0);
  reg [(5'h10):(1'h0)] reg763 = (1'h0);
  reg [(5'h18):(1'h0)] reg762 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg760 = (1'h0);
  reg [(4'h8):(1'h0)] reg758 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg757 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg753 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg751 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg748 = (1'h0);
  reg [(3'h7):(1'h0)] reg745 = (1'h0);
  reg [(5'h19):(1'h0)] reg744 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg743 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg739 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg736 = (1'h0);
  reg [(5'h13):(1'h0)] reg735 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg734 = (1'h0);
  reg [(5'h17):(1'h0)] reg731 = (1'h0);
  reg [(5'h10):(1'h0)] reg730 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg729 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg728 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg727 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg725 = (1'h0);
  reg [(4'hb):(1'h0)] forvar723 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar722 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg721 = (1'h0);
  reg [(5'h1a):(1'h0)] reg719 = (1'h0);
  reg [(4'h8):(1'h0)] reg718 = (1'h0);
  reg [(4'he):(1'h0)] reg717 = (1'h0);
  reg [(5'h17):(1'h0)] reg712 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar711 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg710 = (1'h0);
  assign y = {wire1007,
                 wire1006,
                 wire1005,
                 wire825,
                 wire709,
                 wire708,
                 wire707,
                 reg1060,
                 reg1056,
                 reg1055,
                 reg1053,
                 reg1050,
                 reg1048,
                 reg1044,
                 reg1043,
                 reg1042,
                 reg1039,
                 reg1038,
                 reg1037,
                 reg1035,
                 reg1034,
                 reg1033,
                 reg1031,
                 reg1026,
                 reg1025,
                 reg1024,
                 reg1023,
                 reg1022,
                 reg1020,
                 reg1018,
                 reg1015,
                 reg1013,
                 reg1009,
                 reg1004,
                 reg1003,
                 reg1000,
                 reg998,
                 reg994,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg979,
                 reg978,
                 reg976,
                 reg974,
                 reg972,
                 reg969,
                 reg965,
                 reg962,
                 reg961,
                 reg956,
                 reg954,
                 reg950,
                 reg948,
                 reg943,
                 reg941,
                 reg938,
                 reg928,
                 reg934,
                 reg933,
                 reg932,
                 reg930,
                 reg929,
                 reg926,
                 reg925,
                 reg923,
                 reg919,
                 reg913,
                 reg911,
                 reg909,
                 reg908,
                 reg907,
                 reg905,
                 reg903,
                 reg901,
                 reg900,
                 reg898,
                 reg894,
                 reg892,
                 reg891,
                 reg887,
                 reg886,
                 reg885,
                 reg881,
                 reg880,
                 reg878,
                 reg877,
                 reg875,
                 reg874,
                 reg872,
                 reg870,
                 reg869,
                 reg868,
                 reg862,
                 reg863,
                 reg859,
                 reg849,
                 reg855,
                 reg854,
                 reg853,
                 reg846,
                 reg842,
                 reg841,
                 reg840,
                 reg838,
                 reg836,
                 reg833,
                 reg832,
                 reg831,
                 reg827,
                 reg824,
                 reg821,
                 reg820,
                 reg819,
                 reg815,
                 reg814,
                 reg810,
                 reg809,
                 reg808,
                 reg807,
                 reg790,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 reg797,
                 reg795,
                 reg791,
                 reg784,
                 reg779,
                 reg778,
                 reg777,
                 reg776,
                 reg775,
                 reg773,
                 reg770,
                 reg769,
                 reg768,
                 reg766,
                 reg761,
                 reg759,
                 reg756,
                 reg755,
                 reg754,
                 reg752,
                 reg750,
                 reg749,
                 reg747,
                 reg746,
                 reg742,
                 reg741,
                 reg740,
                 reg738,
                 reg737,
                 reg733,
                 reg732,
                 reg726,
                 reg724,
                 reg720,
                 reg716,
                 reg715,
                 reg714,
                 reg713,
                 reg1066,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1059,
                 forvar1058,
                 forvar1057,
                 reg1054,
                 reg1052,
                 reg1051,
                 forvar1049,
                 forvar1047,
                 reg1046,
                 reg1045,
                 reg1041,
                 forvar1040,
                 forvar1036,
                 reg1032,
                 reg1030,
                 reg1029,
                 forvar1028,
                 reg1027,
                 reg1021,
                 reg1019,
                 reg1017,
                 reg1016,
                 reg1014,
                 forvar1012,
                 reg1011,
                 reg1010,
                 reg1008,
                 reg1002,
                 reg1001,
                 reg999,
                 reg997,
                 reg996,
                 reg995,
                 reg993,
                 forvar992,
                 reg991,
                 reg990,
                 reg989,
                 forvar988,
                 reg987,
                 reg986,
                 reg981,
                 reg980,
                 reg977,
                 forvar975,
                 reg973,
                 reg971,
                 reg970,
                 reg968,
                 forvar967,
                 reg966,
                 reg964,
                 reg963,
                 reg960,
                 reg959,
                 reg958,
                 forvar957,
                 reg955,
                 reg953,
                 forvar952,
                 reg951,
                 reg949,
                 reg947,
                 reg946,
                 reg945,
                 forvar944,
                 reg942,
                 reg940,
                 reg939,
                 reg937,
                 forvar936,
                 reg935,
                 reg931,
                 forvar928,
                 reg927,
                 reg924,
                 reg922,
                 forvar921,
                 reg920,
                 reg918,
                 reg917,
                 reg916,
                 reg915,
                 reg914,
                 reg912,
                 reg910,
                 forvar895,
                 forvar910,
                 reg906,
                 reg904,
                 reg902,
                 reg899,
                 reg897,
                 reg896,
                 reg895,
                 reg893,
                 reg890,
                 reg889,
                 reg888,
                 reg884,
                 reg883,
                 reg882,
                 forvar879,
                 reg876,
                 reg873,
                 reg871,
                 forvar867,
                 reg866,
                 forvar858,
                 reg857,
                 reg865,
                 reg864,
                 forvar862,
                 reg861,
                 reg860,
                 reg858,
                 forvar857,
                 reg856,
                 reg852,
                 reg851,
                 reg850,
                 forvar849,
                 reg848,
                 reg847,
                 reg845,
                 reg844,
                 reg843,
                 reg839,
                 reg837,
                 reg835,
                 forvar834,
                 reg830,
                 forvar829,
                 reg828,
                 forvar826,
                 reg823,
                 reg822,
                 reg818,
                 reg817,
                 reg816,
                 reg813,
                 reg812,
                 reg811,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg798,
                 reg796,
                 reg794,
                 reg793,
                 reg792,
                 forvar790,
                 reg789,
                 reg788,
                 reg787,
                 forvar786,
                 reg785,
                 reg783,
                 reg782,
                 forvar781,
                 reg765,
                 forvar758,
                 forvar741,
                 reg780,
                 reg774,
                 reg772,
                 reg771,
                 reg767,
                 forvar765,
                 reg764,
                 reg763,
                 reg762,
                 reg760,
                 reg758,
                 reg757,
                 reg753,
                 reg751,
                 reg748,
                 reg745,
                 reg744,
                 reg743,
                 reg739,
                 reg736,
                 reg735,
                 reg734,
                 reg731,
                 reg730,
                 reg729,
                 reg728,
                 reg727,
                 reg725,
                 forvar723,
                 forvar722,
                 reg721,
                 reg719,
                 reg718,
                 reg717,
                 reg712,
                 forvar711,
                 reg710,
                 (1'h0)};
  assign wire707 = wire706;
  assign wire708 = (+wire707);
  assign wire709 = wire706[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg710 = $unsigned(wire705[(1'h1):(1'h0)]);
      for (forvar711 = (1'h0); (forvar711 < (3'h4)); forvar711 = (forvar711 + (1'h1)))
        begin
          if (wire707)
            begin
              reg712 = ((((!$signed(forvar711)) || ((wire709 ?
                      (8'hb7) : wire703) + {reg710,
                      (8'ha6)})) >> $unsigned(((+wire706) ~^ (~|wire703)))) ?
                  (^(8'had)) : (wire709 ^ reg710[(1'h0):(1'h0)]));
            end
          else
            begin
              reg712 = (wire703 < ($unsigned(wire703[(3'h7):(3'h5)]) ?
                  wire709[(1'h1):(1'h1)] : (wire708 ?
                      $unsigned(((8'hab) > wire703)) : $unsigned(wire705))));
              reg713 <= $signed((+$signed(((wire709 ~^ wire708) ?
                  reg712[(4'h9):(4'h9)] : $signed((8'hb7))))));
              reg714 <= ((7'h44) <= wire703);
            end
          if (reg712)
            begin
              reg715 <= {(wire708[(1'h0):(1'h0)] ? {(|wire703)} : (7'h4d)),
                  {{reg712, $signed((wire705 | reg710)), wire708}, reg712},
                  $unsigned((~^(7'h4c)))};
              reg716 <= reg714[(2'h2):(2'h2)];
              reg717 = $unsigned((($signed((~(8'h9c))) >= (reg712[(4'hc):(4'ha)] ?
                      (wire704 ? reg714 : reg714) : (+wire705))) ?
                  {wire704[(4'hb):(3'h4)],
                      ((wire706 + (8'h9e)) ?
                          $signed(reg714) : $signed(forvar711)),
                      forvar711} : $unsigned(wire708)));
              reg718 = ($unsigned({$signed(reg717),
                      $signed($signed((8'hb2))),
                      ($unsigned(wire703) ?
                          (wire707 ?
                              forvar711 : wire706) : $unsigned(reg713))}) ?
                  ((((wire705 ?
                      wire705 : wire709) < (~|wire706)) ^~ $signed(wire708)) ~^ (&($unsigned(wire704) ?
                      reg712 : (~|wire709)))) : $signed(wire703));
              reg719 = (|{((wire708[(2'h3):(1'h0)] ^~ (reg713 ?
                          reg715 : reg710)) ?
                      reg717[(3'h5):(1'h1)] : {$unsigned(reg716),
                          (wire708 || wire707),
                          $signed(wire703)})});
              reg720 <= ((^~reg717[(4'hd):(3'h5)]) ?
                  (|$unsigned(reg716[(1'h0):(1'h0)])) : $signed({(&$signed(reg714)),
                      reg710[(4'h9):(3'h5)]}));
            end
          else
            begin
              reg715 <= wire703;
              reg716 <= reg713[(4'h9):(2'h3)];
              reg717 = ($signed(reg715[(3'h6):(3'h6)]) >= $signed((&(+{reg712,
                  (8'ha7)}))));
              reg718 = ($signed(reg717) != (($unsigned($unsigned(reg719)) ?
                      (7'h40) : ($unsigned(reg717) ?
                          (forvar711 * reg712) : reg712)) ?
                  $unsigned($signed($unsigned((8'h9f)))) : wire708[(2'h3):(2'h2)]));
            end
          reg721 = wire704[(3'h7):(1'h1)];
        end
      for (forvar722 = (1'h0); (forvar722 < (2'h2)); forvar722 = (forvar722 + (1'h1)))
        begin
          for (forvar723 = (1'h0); (forvar723 < (3'h6)); forvar723 = (forvar723 + (1'h1)))
            begin
              reg724 <= ((~&((wire709 ?
                  wire708 : wire704[(3'h6):(1'h0)]) && $signed((~&reg710)))) || $signed(wire707[(1'h0):(1'h0)]));
              reg725 = $signed((reg716[(1'h1):(1'h0)] ?
                  (((forvar723 ?
                      reg713 : wire709) ^ forvar711) && (reg713 * (reg713 ?
                      reg710 : reg717))) : (reg714 ?
                      ($signed(forvar723) ?
                          {reg716,
                              forvar723} : $unsigned(reg718)) : wire708[(2'h2):(2'h2)])));
              reg726 <= (~{((-wire704[(1'h0):(1'h0)]) ?
                      (wire705 ?
                          (-wire706) : wire707[(5'h10):(1'h1)]) : ({reg725,
                          reg725} >= $signed(wire705))),
                  ((+reg719) >> reg715[(4'ha):(3'h7)]),
                  (((~&(8'hb1)) ?
                      $signed(wire703) : $unsigned(reg717)) << wire708[(2'h2):(2'h2)])});
              reg727 = forvar711[(4'hd):(2'h2)];
              reg728 = (($signed((+$signed(forvar722))) ?
                      reg717 : $unsigned(wire708)) ?
                  $unsigned($signed($unsigned((^~wire706)))) : ((-$unsigned((~^(8'ha4)))) >= $unsigned(forvar723[(2'h2):(1'h1)])));
              reg729 = reg721;
              reg730 = ($unsigned(($signed((8'ha2)) ?
                  {(reg721 <<< reg718),
                      (~|reg724),
                      reg721} : reg727[(3'h7):(3'h7)])) >> $unsigned(((forvar722 ?
                  (|wire706) : (-wire705)) >>> $unsigned({(7'h58),
                  forvar711}))));
            end
          if (reg719)
            begin
              reg731 = $unsigned(((((7'h48) ?
                          $unsigned(reg724) : $signed(wire705)) ?
                      $unsigned($signed((8'hbb))) : $signed(reg729)) ?
                  (~^((reg729 ? wire704 : (8'ha7)) ?
                      {reg712, reg718} : {wire708,
                          reg720})) : (~^$signed($signed(reg720)))));
              reg732 <= $unsigned((~^wire705));
              reg733 <= ({forvar722, reg719[(3'h6):(3'h5)]} ?
                  $unsigned(({(reg718 ?
                          reg716 : wire703)} || reg728[(4'h9):(2'h3)])) : $signed(reg725[(3'h6):(1'h1)]));
              reg734 = reg726[(3'h4):(2'h2)];
              reg735 = reg712;
              reg736 = reg714[(2'h2):(2'h2)];
              reg737 <= reg733[(5'h15):(5'h11)];
            end
          else
            begin
              reg731 = (!(+(($signed((7'h46)) - (|reg717)) < ((reg715 ~^ forvar711) * (reg718 ?
                  reg736 : reg732)))));
              reg732 <= $unsigned($unsigned((~&($unsigned(reg710) - $signed(wire704)))));
              reg734 = forvar711[(3'h7):(3'h5)];
              reg735 = $unsigned($signed({{(wire703 ^ (7'h58)),
                      forvar711[(4'hb):(4'h9)]}}));
            end
          reg738 <= (((reg717 ? ({reg710} ~^ (^~(8'hb2))) : reg713) ?
                  (($unsigned(reg718) ?
                      ((7'h41) ?
                          reg718 : (8'h9c)) : $unsigned(reg725)) < $signed((reg735 ?
                      reg724 : reg728))) : $unsigned($unsigned(reg715))) ?
              ((((reg728 ? wire709 : reg729) >> $unsigned((8'hba))) ?
                  {(^wire706),
                      reg724[(2'h3):(1'h0)],
                      reg737[(5'h18):(1'h1)]} : ($unsigned((7'h49)) ?
                      (8'ha9) : (^~forvar711))) - reg724[(1'h0):(1'h0)]) : $signed((reg732[(4'h8):(3'h4)] ?
                  $unsigned($unsigned((7'h48))) : (8'h9f))));
        end
      reg739 = $unsigned($unsigned($signed(reg715)));
      if ($signed($unsigned({(~reg715)})))
        begin
          if (reg716[(2'h2):(1'h0)])
            begin
              reg740 <= $unsigned($signed((8'hb2)));
              reg741 <= (reg738[(4'hc):(4'ha)] ?
                  (wire709[(1'h0):(1'h0)] ?
                      ($signed(reg724) ?
                          $unsigned($unsigned(reg726)) : reg726) : reg734[(4'hf):(4'h9)]) : (~|reg713));
              reg742 <= $unsigned((^~(8'hb2)));
              reg743 = (reg721 + $signed($unsigned($signed($signed(reg742)))));
              reg744 = $signed(($unsigned({reg710, (8'hb6), reg739}) ?
                  $signed($unsigned((^~(7'h43)))) : $unsigned(reg710[(4'h9):(1'h1)])));
              reg745 = ((~^{$unsigned((reg728 >= wire703))}) ^ $unsigned(reg730));
            end
          else
            begin
              reg743 = $signed(wire708[(1'h1):(1'h0)]);
              reg746 <= wire707[(3'h6):(3'h6)];
              reg747 <= reg744;
            end
          if ($signed(reg735))
            begin
              reg748 = reg739;
              reg749 <= reg725[(3'h6):(3'h5)];
              reg750 <= {(~reg726),
                  $unsigned((~((reg745 ?
                      reg728 : reg726) ^ $unsigned(reg730))))};
              reg751 = ((|reg739[(2'h2):(1'h0)]) ?
                  (reg727[(5'h14):(3'h4)] ?
                      ((8'ha4) ?
                          wire704[(1'h0):(1'h0)] : $unsigned({forvar723})) : (8'ha7)) : $signed({($signed(reg728) ?
                          reg732[(5'h10):(3'h4)] : reg747)}));
              reg752 <= (reg750[(4'hc):(3'h5)] ?
                  $unsigned((&$signed(wire703[(3'h7):(2'h3)]))) : ({{reg721[(2'h2):(2'h2)],
                              wire708,
                              $signed(reg751)},
                          ((&reg745) & (+reg739))} ?
                      reg718 : reg743[(5'h15):(4'ha)]));
            end
          else
            begin
              reg749 <= ($signed((reg745 < (reg720[(3'h7):(3'h5)] >= (+reg744)))) + reg725);
              reg751 = $unsigned((reg715[(1'h0):(1'h0)] ?
                  ((reg724[(1'h1):(1'h0)] << (8'ha7)) != (~reg729)) : (~(!(reg736 < reg750)))));
              reg753 = ($unsigned(reg749) <<< ($unsigned(wire707) ?
                  reg737[(4'hf):(4'hf)] : $signed(reg747)));
              reg754 <= (7'h50);
              reg755 <= ($signed(reg737) ? reg743 : reg741[(4'hc):(1'h0)]);
              reg756 <= $signed((^~reg727[(2'h2):(1'h1)]));
              reg757 = (({wire705,
                      (reg727[(5'h10):(4'hc)] ?
                          reg728[(4'ha):(1'h1)] : (wire708 ? reg740 : reg728)),
                      reg743} ?
                  (forvar722 - ((+wire705) ?
                      ((8'ha3) ? reg712 : reg727) : (forvar711 ?
                          reg727 : (8'h9d)))) : (~((reg710 ? wire709 : reg731) ?
                      $signed(reg720) : $signed((7'h4d))))) < (($unsigned({reg736,
                      wire706}) ?
                  (^$signed(reg732)) : (-(reg718 ?
                      (7'h51) : reg718))) > reg734));
            end
          reg758 = $unsigned(reg738[(3'h4):(1'h1)]);
          if ($signed((wire708[(2'h2):(1'h1)] <<< ((reg733[(5'h11):(4'hf)] ^~ $unsigned((8'hb2))) << reg727[(3'h5):(1'h1)]))))
            begin
              reg759 <= $signed($unsigned((((reg719 ? reg719 : reg715) ?
                      $unsigned(reg720) : {reg717, reg710}) ?
                  $signed((reg719 >> reg713)) : reg753[(1'h1):(1'h0)])));
              reg760 = {$unsigned(($signed($signed(reg727)) | $unsigned((reg725 ?
                      reg713 : reg753)))),
                  (~&$unsigned(((reg754 ? reg756 : reg745) ?
                      {(8'hae), forvar722, wire703} : (~|reg725)))),
                  (reg717 ?
                      (forvar711 <= $signed((reg736 ?
                          (7'h4d) : reg715))) : reg752[(1'h0):(1'h0)])};
            end
          else
            begin
              reg759 <= {$signed($unsigned($unsigned((reg728 <= reg759)))),
                  (reg751 ? forvar723 : reg740[(4'h8):(4'h8)]),
                  (&(^~reg719))};
              reg760 = (!$signed(($unsigned((reg731 ?
                  forvar723 : reg753)) > (&(reg757 ? (8'h9e) : reg718)))));
              reg761 <= $unsigned((~&{(reg751 ?
                      (forvar723 ? (8'haa) : forvar711) : reg758),
                  ((reg740 ? reg720 : reg760) ? (~|reg720) : reg724)}));
              reg762 = $unsigned((^($signed((&reg738)) != $signed($unsigned(reg758)))));
              reg763 = (reg720 << (reg758[(1'h0):(1'h0)] ?
                  ((~|(reg737 > reg748)) || (reg747[(4'h9):(3'h5)] ?
                      $signed(reg730) : (wire703 ?
                          reg720 : reg749))) : (^(~^reg736[(2'h2):(1'h0)]))));
              reg764 = (~|(reg755[(5'h13):(1'h0)] <<< $unsigned((8'ha4))));
            end
          for (forvar765 = (1'h0); (forvar765 < (1'h0)); forvar765 = (forvar765 + (1'h1)))
            begin
              reg766 <= (reg749[(1'h1):(1'h0)] ?
                  $unsigned((^$signed((!reg753)))) : ($signed(($signed(reg725) ?
                          (reg763 & reg736) : $signed(reg756))) ?
                      $signed(((wire708 > reg747) >>> $unsigned((8'hbc)))) : (((forvar723 ?
                                  (7'h57) : (8'ha6)) ?
                              (~&reg717) : $unsigned((8'ha7))) ?
                          (!reg760) : ((^~reg715) >>> ((8'ha0) << wire708)))));
              reg767 = {$unsigned(({(7'h4f),
                      (reg757 ?
                          reg735 : reg724)} - $signed(wire707[(4'h9):(1'h1)]))),
                  {$signed({$signed(reg724)})}};
              reg768 <= reg756;
              reg769 <= $unsigned((~&reg736));
              reg770 <= (7'h44);
              reg771 = reg766;
            end
          reg772 = (&$unsigned((reg751 ?
              reg728[(2'h2):(1'h1)] : $unsigned((forvar765 ?
                  reg754 : reg741)))));
          if ((7'h47))
            begin
              reg773 <= reg725;
              reg774 = wire709;
            end
          else
            begin
              reg773 <= ($signed(($signed(reg718[(4'h8):(3'h4)]) ?
                  forvar765 : forvar722[(4'h9):(3'h6)])) == (reg753[(1'h1):(1'h0)] ?
                  reg743 : (reg721 ^~ reg729[(4'he):(2'h3)])));
              reg775 <= {(8'hba),
                  $unsigned((8'ha2)),
                  {$unsigned(((~&reg733) >>> (~^(7'h46)))),
                      ((|(reg766 > reg721)) ?
                          $signed(reg774) : $signed(((8'h9e) - reg742))),
                      reg710[(4'hc):(4'hc)]}};
              reg776 <= reg724;
              reg777 <= ($signed($signed($signed((+reg745)))) ?
                  (-$signed(($unsigned(reg732) ^~ reg717))) : forvar711[(2'h2):(2'h2)]);
              reg778 <= reg770;
              reg779 <= (($unsigned(($signed(reg761) == {wire708})) ?
                  ($signed($unsigned(reg778)) * (8'hb7)) : wire703) >= reg712);
              reg780 = reg720;
            end
        end
      else
        begin
          reg740 <= ($unsigned(reg724) ~^ $signed(reg755[(5'h18):(3'h5)]));
          for (forvar741 = (1'h0); (forvar741 < (3'h4)); forvar741 = (forvar741 + (1'h1)))
            begin
              reg743 = $unsigned($signed($signed((reg746 - (-reg767)))));
            end
          reg746 <= $signed({$signed($signed((wire705 > reg721))),
              $signed(forvar741),
              reg741});
          if (reg724[(1'h1):(1'h0)])
            begin
              reg747 <= $unsigned($unsigned(reg716));
              reg748 = (^$signed((reg737[(5'h13):(4'hf)] ?
                  reg718[(2'h3):(2'h2)] : (reg778 ?
                      (reg749 ? wire706 : reg747) : (-reg746)))));
              reg749 <= (~$unsigned({$signed($signed(reg773)),
                  reg764[(3'h4):(2'h2)],
                  $unsigned($unsigned(reg755))}));
              reg751 = ($unsigned((8'had)) - (reg751[(4'hb):(2'h3)] <= {((7'h55) ?
                      reg710 : (reg769 ? reg769 : forvar765)),
                  ($signed(reg759) ?
                      ((7'h55) ? (7'h46) : forvar723) : $unsigned(reg753)),
                  (^$unsigned(reg728))}));
            end
          else
            begin
              reg747 <= (~&reg742[(3'h7):(3'h7)]);
              reg749 <= reg752;
              reg751 = (($unsigned(reg777) >> reg772) ?
                  reg761[(4'ha):(4'ha)] : ($unsigned({(reg713 ?
                          (8'hb0) : reg770),
                      (reg737 ^~ (8'hb4)),
                      reg740}) <<< {$unsigned((-reg719)), $unsigned(wire704)}));
              reg752 <= $unsigned(($unsigned({(reg717 ? reg739 : reg750),
                  $unsigned(reg720)}) != reg764[(1'h0):(1'h0)]));
              reg754 <= wire704[(3'h5):(2'h2)];
              reg757 = ($unsigned({((reg741 - reg772) ?
                          (reg768 ? reg762 : forvar765) : {forvar723,
                              reg724,
                              reg745})}) ?
                  $signed((((reg735 ? forvar723 : reg740) == (forvar741 ?
                          forvar723 : reg744)) ?
                      ($unsigned(forvar723) ?
                          reg720 : reg733[(5'h1c):(1'h0)]) : reg740)) : ($signed($unsigned((!forvar765))) ?
                      $unsigned((8'hbe)) : reg720));
            end
          for (forvar758 = (1'h0); (forvar758 < (3'h4)); forvar758 = (forvar758 + (1'h1)))
            begin
              reg759 <= (reg775[(5'h13):(5'h13)] ?
                  ({$unsigned($unsigned((8'ha9))), (~(^(7'h53)))} ?
                      (8'ha5) : $signed(((-reg718) ?
                          (-reg767) : (reg748 ?
                              reg738 : reg753)))) : ((|((reg754 <<< reg759) ?
                          (8'ha6) : ((8'hb3) != reg736))) ?
                      (((7'h4b) ?
                          (reg717 ?
                              reg755 : reg772) : ((8'ha8) & reg767)) >>> ((^reg716) ?
                          (reg747 << (7'h51)) : $unsigned(reg747))) : ((7'h52) ?
                          ((+reg755) || $signed(reg737)) : $unsigned($signed(forvar722)))));
              reg760 = $unsigned((reg725 ?
                  $unsigned($unsigned({reg752,
                      reg776,
                      reg776})) : ($signed((reg760 >= reg756)) ?
                      $signed({(7'h46)}) : $unsigned(reg760[(4'h8):(3'h5)]))));
            end
          if (reg744)
            begin
              reg762 = reg736;
              reg763 = (-reg750[(2'h3):(1'h0)]);
              reg764 = $unsigned(($unsigned($signed((~^reg769))) ?
                  (reg760 >>> $unsigned($signed(reg715))) : $unsigned(reg720[(5'h12):(2'h2)])));
              reg765 = (reg735 ?
                  reg768 : (reg772 ?
                      (($signed(reg748) <= (reg777 > reg756)) ?
                          ((reg737 ^ reg730) ?
                              {(8'hb5),
                                  reg780,
                                  reg725} : $signed((8'hbb))) : ((reg778 ^~ reg778) ?
                              $signed(reg757) : $signed(reg720))) : $unsigned({(~^reg761),
                          (reg754 ^ reg772)})));
              reg767 = $unsigned({($signed(reg737) == reg729),
                  reg761[(2'h2):(1'h1)]});
              reg771 = ($signed(forvar722) ?
                  ((|$unsigned($unsigned(forvar722))) * $signed(({reg731,
                          reg772,
                          (7'h43)} ?
                      ((8'hac) >> reg775) : $signed(forvar758)))) : reg764[(1'h1):(1'h1)]);
            end
          else
            begin
              reg762 = (^~$unsigned($signed({$signed((7'h48)),
                  {reg747, reg714},
                  wire708[(1'h1):(1'h1)]})));
              reg766 <= {(reg741[(5'h18):(4'hc)] ?
                      reg750[(4'hb):(4'h9)] : forvar723),
                  $unsigned(((|((8'had) <= reg712)) ?
                      reg760[(3'h4):(3'h4)] : (+{reg712, reg779, (8'hbb)}))),
                  ((($signed(reg743) ?
                          reg748 : (reg721 != reg726)) <<< (7'h46)) ?
                      (~|(~&(reg769 ^ reg731))) : ($unsigned($unsigned((8'hb4))) || $unsigned((&reg745))))};
              reg767 = $signed(((reg717[(1'h0):(1'h0)] ?
                      (~^reg738) : wire703[(4'hd):(4'h9)]) ?
                  $unsigned((+$unsigned(reg710))) : reg730[(4'hb):(3'h6)]));
              reg771 = $unsigned((reg758[(2'h2):(1'h1)] ^~ reg755));
              reg772 = {$unsigned(reg757), (8'hbe), (8'ha2)};
              reg773 <= reg760[(5'h1c):(5'h11)];
              reg775 <= {(8'ha3), $unsigned($signed(wire705[(4'hc):(4'h8)]))};
            end
        end
      for (forvar781 = (1'h0); (forvar781 < (3'h4)); forvar781 = (forvar781 + (1'h1)))
        begin
          reg782 = ($signed($signed((8'h9c))) != (+(|(7'h41))));
          reg783 = (7'h54);
          reg784 <= (+(reg759[(1'h0):(1'h0)] > reg753));
          reg785 = reg745;
          for (forvar786 = (1'h0); (forvar786 < (3'h4)); forvar786 = (forvar786 + (1'h1)))
            begin
              reg787 = (~&(7'h4b));
            end
          reg788 = reg721;
        end
    end
  always
    @(posedge clk) begin
      reg789 = (((7'h46) ?
              (~|(wire703 - $signed(wire703))) : (($signed(reg726) ?
                      (8'ha8) : $unsigned(wire709)) ?
                  reg740 : ($unsigned(reg741) << reg770))) ?
          reg714 : ($signed((reg741 >>> wire706[(3'h5):(1'h0)])) ?
              (~^reg713) : $unsigned(((reg778 <= reg766) ?
                  $signed(reg746) : reg732[(5'h18):(5'h18)]))));
      if (($unsigned(reg749) ?
          (-($unsigned(wire704[(3'h7):(3'h4)]) ?
              wire705[(1'h0):(1'h0)] : ($signed((7'h46)) * $unsigned(reg720)))) : reg776))
        begin
          for (forvar790 = (1'h0); (forvar790 < (2'h2)); forvar790 = (forvar790 + (1'h1)))
            begin
              reg791 <= {wire707,
                  $unsigned(({reg742} ?
                      (reg714 ?
                          $signed(reg740) : $unsigned(reg746)) : $signed($signed(reg724))))};
              reg792 = $signed({($signed((reg715 | reg750)) ?
                      ({reg766, reg746} ?
                          reg747[(2'h3):(1'h0)] : (|(8'hbf))) : {((7'h55) == reg732)}),
                  reg726,
                  reg778});
              reg793 = reg714[(1'h0):(1'h0)];
            end
          reg794 = reg741[(5'h14):(5'h10)];
          if ((reg715 ^~ {(reg759 ? reg773 : (^reg746[(2'h2):(2'h2)])),
              wire709}))
            begin
              reg795 <= (reg777 ?
                  (reg726[(3'h6):(1'h0)] ^~ (~^$signed((+reg775)))) : (8'hab));
              reg796 = $signed($unsigned((|{{reg738, reg775}})));
              reg797 <= reg779[(3'h6):(1'h0)];
              reg798 = (8'h9e);
              reg799 <= (-reg766);
            end
          else
            begin
              reg795 <= reg740[(1'h0):(1'h0)];
              reg797 <= $signed(reg778[(3'h6):(2'h3)]);
              reg799 <= $signed(($unsigned($unsigned($unsigned((8'haf)))) ?
                  $signed($signed({reg754,
                      reg733})) : (($signed(reg793) && $signed(reg724)) ?
                      ((reg754 ?
                          wire709 : reg793) ^~ (~wire707)) : reg768[(1'h1):(1'h1)])));
              reg800 <= reg755[(3'h7):(3'h5)];
              reg801 <= (7'h40);
              reg802 <= ($signed(wire705) * ($unsigned((reg715 ?
                      $unsigned(wire707) : $signed(wire706))) ?
                  wire706[(5'h10):(4'he)] : $unsigned((((8'ha7) ?
                          reg776 : reg795) ?
                      $signed(reg769) : $unsigned(reg766)))));
            end
        end
      else
        begin
          if (reg802)
            begin
              reg790 <= (-$signed((reg746[(2'h2):(1'h1)] | $signed($signed(reg766)))));
              reg792 = $unsigned(wire708[(1'h0):(1'h0)]);
              reg793 = (~^{{((+reg800) ?
                          (reg726 ~^ reg752) : reg761[(1'h1):(1'h1)]),
                      {reg746},
                      (|{reg795})}});
              reg795 <= reg766[(5'h11):(4'hb)];
              reg796 = (~&((~|((8'h9e) ? (8'hb8) : $unsigned(reg790))) ?
                  $unsigned(forvar790) : (reg716 ?
                      ((!(8'hb9)) ?
                          reg769 : reg750) : $signed($unsigned((8'hb6))))));
              reg798 = reg797[(4'h8):(2'h3)];
              reg803 = reg740;
            end
          else
            begin
              reg790 <= $signed($unsigned($signed((8'ha0))));
              reg792 = reg756;
              reg795 <= reg773[(4'ha):(4'h9)];
              reg796 = reg750;
              reg798 = $unsigned((!$unsigned((~^(^reg775)))));
              reg803 = (~reg713);
              reg804 = ((|(^$unsigned(reg754[(4'he):(4'hd)]))) - (reg784 ?
                  ($unsigned($signed((7'h4f))) ?
                      $unsigned((8'ha8)) : $unsigned(reg755[(1'h0):(1'h0)])) : ((reg794[(5'h16):(1'h0)] ?
                      ((7'h53) ?
                          reg750 : reg713) : reg799) >>> $unsigned($signed(reg747)))));
            end
          reg805 = $signed((({$unsigned(reg747)} >> reg797[(5'h13):(4'he)]) ?
              ((!$unsigned(reg768)) - reg713) : ((^$signed(reg733)) - reg715[(4'hb):(3'h4)])));
          if ((~|$unsigned(reg766[(5'h10):(4'hf)])))
            begin
              reg806 = reg803;
              reg807 <= reg756;
              reg808 <= wire708;
              reg809 <= (~^reg755[(2'h2):(1'h1)]);
            end
          else
            begin
              reg807 <= $signed({$unsigned(((^reg724) ?
                      {reg716, reg777} : (reg807 < (8'ha7)))),
                  $unsigned((8'hab))});
            end
          if ($signed(wire704))
            begin
              reg810 <= $signed((((((8'hb2) != wire706) ?
                  reg726[(4'hc):(1'h1)] : (reg742 * wire704)) <= ((8'hb8) ?
                  (reg778 ? reg798 : reg756) : (reg793 >> reg807))) ^ reg756));
              reg811 = (({forvar790[(3'h4):(2'h2)]} << reg773) != (~^{(((7'h46) ?
                      reg807 : reg732) != $signed(reg777))}));
              reg812 = (reg798[(4'h8):(1'h0)] && ((8'h9f) > (~|$unsigned(reg801))));
              reg813 = ($unsigned(((&reg754[(4'h9):(3'h7)]) ?
                      $signed((~|reg790)) : reg770)) ?
                  reg811[(4'hc):(4'h9)] : $signed(($signed((forvar790 ^ reg714)) >>> (+(reg741 ~^ (8'ha7))))));
            end
          else
            begin
              reg811 = {($unsigned($unsigned((-reg773))) ?
                      (-(reg769 >= (~&reg756))) : ((&(reg714 ~^ reg756)) == ($unsigned(reg749) ~^ reg716))),
                  ({reg746[(2'h2):(1'h1)],
                          ($unsigned(reg778) & $unsigned(reg714))} ?
                      (~$unsigned((|reg810))) : $signed(reg747)),
                  {(^{(reg775 && wire704), $unsigned(reg766)}),
                      reg713,
                      reg801}};
              reg814 <= reg795;
              reg815 <= $signed($signed((7'h42)));
              reg816 = {((($signed(reg810) ? $signed((7'h52)) : forvar790) ?
                      ((reg800 ? reg740 : reg807) >= {reg789,
                          reg713,
                          reg740}) : (^(~^(8'hb6)))) - $unsigned(reg792[(4'ha):(3'h7)]))};
              reg817 = ($unsigned((^~(^~reg779[(5'h14):(4'hc)]))) ?
                  reg816 : (reg816 ?
                      {(~&(reg794 ? (7'h4f) : reg815)),
                          ((!reg805) ? reg796 : (8'had)),
                          ($signed(reg792) ?
                              (reg716 != (7'h4f)) : reg789)} : reg747[(4'h8):(4'h8)]));
              reg818 = (8'hb8);
            end
          if ($unsigned(($signed($unsigned(reg807)) ?
              reg741[(2'h2):(2'h2)] : reg715[(4'hb):(1'h1)])))
            begin
              reg819 <= $signed(reg750[(4'hb):(2'h3)]);
              reg820 <= (((|(reg761[(3'h7):(2'h2)] ?
                          $unsigned(reg816) : reg811[(4'h8):(3'h6)])) ?
                      {reg733} : {($unsigned(reg804) ?
                              reg778[(4'h8):(3'h7)] : (&reg737)),
                          ((reg814 ? reg770 : reg766) & (~^reg742))}) ?
                  reg801 : wire708);
              reg821 <= (~|((8'hae) || (~(&{(7'h58)}))));
              reg822 = (($unsigned(wire709) && {$unsigned((reg737 ^~ reg773)),
                  ($signed(reg759) <<< (&wire703)),
                  ($signed(reg726) ?
                      $signed(reg778) : $unsigned(reg715))}) ^ reg716[(1'h1):(1'h1)]);
              reg823 = ($unsigned($unsigned(({reg801} | reg752))) * (!wire709[(2'h3):(1'h0)]));
            end
          else
            begin
              reg819 <= ((reg749 ?
                      $unsigned($signed(reg769)) : {$unsigned(reg779),
                          (reg713 ? (reg822 >>> (7'h57)) : $signed(wire706)),
                          (!reg796)}) ?
                  reg738[(4'hf):(1'h1)] : $signed($signed(({reg714} ?
                      reg790[(3'h5):(1'h0)] : (reg755 ~^ reg792)))));
            end
        end
      reg824 <= {reg794[(5'h11):(4'he)],
          ((($signed(wire709) ? (-reg738) : reg775) << wire705) ?
              reg821 : ({reg732[(5'h1e):(5'h17)],
                  (-reg806),
                  (&wire706)} == $unsigned((~reg790))))};
    end
  assign wire825 = (-((reg801[(1'h1):(1'h1)] ?
                       $unsigned(((7'h40) << reg732)) : (reg815[(3'h6):(3'h5)] ?
                           reg770[(4'hb):(4'hb)] : (wire709 != reg799))) >= {reg777}));
  always
    @(posedge clk) begin
      for (forvar826 = (1'h0); (forvar826 < (1'h1)); forvar826 = (forvar826 + (1'h1)))
        begin
          reg827 <= $unsigned($signed(reg809[(5'h13):(1'h1)]));
          reg828 = (8'haf);
          for (forvar829 = (1'h0); (forvar829 < (3'h5)); forvar829 = (forvar829 + (1'h1)))
            begin
              reg830 = reg768;
              reg831 <= reg750;
            end
          reg832 <= ((reg820 ?
              forvar829 : $signed($unsigned((7'h47)))) < {reg726, (7'h41)});
          reg833 <= reg778[(3'h5):(1'h1)];
          for (forvar834 = (1'h0); (forvar834 < (3'h5)); forvar834 = (forvar834 + (1'h1)))
            begin
              reg835 = reg720[(4'hd):(4'hd)];
              reg836 <= (~&$unsigned(reg759[(1'h1):(1'h0)]));
              reg837 = ((-reg830[(3'h4):(1'h1)]) ?
                  reg819[(4'h8):(2'h3)] : reg810);
              reg838 <= reg836;
              reg839 = (^wire825);
              reg840 <= $unsigned((~($unsigned($signed(reg720)) ?
                  ((^~(8'hba)) ?
                      $unsigned(reg828) : (reg714 <<< reg833)) : ((reg824 || reg779) ?
                      $signed(reg766) : $unsigned(wire825)))));
              reg841 <= (({reg784[(2'h3):(1'h1)]} < {$signed(reg838),
                  reg819}) <= $signed(reg755));
            end
        end
      if (reg795[(4'h8):(3'h4)])
        begin
          if ($signed(reg766[(5'h17):(4'hc)]))
            begin
              reg842 <= reg777[(4'he):(3'h4)];
              reg843 = (&reg769);
              reg844 = reg775[(3'h7):(1'h1)];
              reg845 = (^reg814[(3'h6):(1'h0)]);
              reg846 <= reg715[(4'hd):(3'h7)];
              reg847 = (reg814[(1'h1):(1'h1)] ?
                  reg742 : (-$signed(reg839[(4'ha):(3'h5)])));
              reg848 = $signed((~(reg756 ?
                  (reg724 ?
                      ((7'h4e) > (7'h55)) : reg807) : $signed((|reg828)))));
            end
          else
            begin
              reg842 <= (+$signed($unsigned(reg779[(4'h9):(2'h3)])));
              reg843 = (((~reg841[(4'h8):(4'h8)]) ?
                  forvar826 : ($unsigned($unsigned(reg832)) ^ {$signed(reg726),
                      (&wire825),
                      (reg713 <= reg761)})) | (|$unsigned(($signed(reg761) + $unsigned(reg732)))));
              reg846 <= {reg769[(3'h4):(1'h1)]};
            end
          for (forvar849 = (1'h0); (forvar849 < (2'h3)); forvar849 = (forvar849 + (1'h1)))
            begin
              reg850 = (reg820 ?
                  $signed($unsigned($signed((wire825 ?
                      reg830 : wire704)))) : (8'hbd));
              reg851 = (-reg807[(5'h12):(5'h12)]);
              reg852 = $unsigned(({$unsigned((reg761 <<< forvar834)),
                  $unsigned((+reg726))} - wire704[(3'h7):(3'h7)]));
              reg853 <= $unsigned({$unsigned((^reg852[(2'h2):(1'h1)])),
                  $unsigned(((reg820 <<< wire709) * (!reg848))),
                  (~|$unsigned(reg842[(2'h2):(2'h2)]))});
            end
          reg854 <= $signed(reg838[(2'h3):(1'h1)]);
          reg855 <= $unsigned(reg846);
        end
      else
        begin
          if ($signed({reg838[(1'h0):(1'h0)]}))
            begin
              reg842 <= reg848[(2'h3):(2'h3)];
              reg843 = (!$unsigned((-(8'hbb))));
            end
          else
            begin
              reg843 = ($unsigned((((&wire706) ?
                  $signed(reg800) : {reg847,
                      reg852}) ^~ (&reg791))) ^ (~|($unsigned((7'h48)) ?
                  reg759 : $signed((reg844 <= (8'hb3))))));
              reg844 = (-{(reg837 ?
                      (reg855 >= reg814[(4'ha):(2'h2)]) : (reg855[(1'h1):(1'h1)] ?
                          (!reg847) : (reg852 ? reg831 : (7'h40)))),
                  (7'h43)});
            end
          if (((^(+$signed(reg716))) ?
              $signed({$unsigned((+reg713)),
                  (7'h4b)}) : $signed($unsigned(reg844[(4'hc):(3'h7)]))))
            begin
              reg846 <= forvar826;
              reg847 = (($signed(($signed(reg759) | wire708)) ?
                  (-{(-wire704)}) : $signed($unsigned({reg845,
                      (8'had),
                      reg808}))) >= reg775);
              reg848 = $signed(reg777[(1'h1):(1'h0)]);
              reg849 <= reg850;
              reg850 = ((~^($unsigned($signed((7'h54))) + ((reg779 ?
                          reg761 : reg855) ?
                      $signed(reg740) : (8'haf)))) ?
                  reg773[(2'h2):(1'h1)] : ((&($signed(reg776) ?
                          $signed(wire709) : $unsigned(reg838))) ?
                      $unsigned((wire704[(1'h1):(1'h0)] ?
                          (reg797 ^ reg832) : reg852[(3'h5):(2'h3)])) : ($signed({reg746}) >>> reg759[(2'h2):(1'h1)])));
              reg851 = (+((~|((reg841 == (8'hba)) ?
                      (~reg773) : (reg769 - reg831))) ?
                  (reg747 ?
                      $unsigned((^(8'h9f))) : (^~(reg821 ?
                          reg853 : reg840))) : {{reg713[(1'h1):(1'h0)],
                          reg724[(1'h1):(1'h1)],
                          $unsigned(reg791)}}));
            end
          else
            begin
              reg846 <= {$signed(((forvar829 ?
                      reg773 : reg784) - ($unsigned(reg840) < reg828[(2'h2):(2'h2)]))),
                  (reg754 ?
                      {reg844[(1'h0):(1'h0)],
                          (8'hbe)} : ((-$unsigned(reg830)) <= ($unsigned(reg809) - $signed(reg724)))),
                  $unsigned($unsigned((~$signed(wire705))))};
              reg847 = (((&reg790[(1'h0):(1'h0)]) ^ reg843[(1'h1):(1'h1)]) && ((+((reg742 && reg755) != reg720)) ?
                  (|{(-reg841),
                      (reg778 && (8'hb6)),
                      wire709[(3'h5):(2'h2)]}) : ($signed($unsigned(reg810)) > $unsigned((|reg845)))));
              reg848 = (reg852 ?
                  reg850[(5'h15):(5'h10)] : reg790[(2'h2):(2'h2)]);
              reg850 = forvar826;
              reg851 = $signed((7'h53));
              reg852 = (reg827[(4'he):(1'h0)] ?
                  $unsigned({$unsigned((~forvar849)),
                      $signed(((8'h9c) ? reg754 : (7'h44))),
                      ($signed((8'hbf)) ?
                          $signed(reg716) : reg752[(2'h2):(2'h2)])}) : (reg820[(2'h3):(2'h2)] ?
                      (&(&$signed((7'h49)))) : ({(reg841 ? reg777 : reg761),
                              (forvar829 ? reg732 : wire709),
                              $unsigned(reg776)} ?
                          ($signed((7'h54)) ?
                              (reg831 ?
                                  wire709 : reg714) : reg840) : $unsigned(reg831))));
            end
          reg856 = $signed(reg843[(2'h2):(1'h1)]);
        end
      if ((-$signed($signed($unsigned($signed((8'hb6)))))))
        begin
          for (forvar857 = (1'h0); (forvar857 < (3'h4)); forvar857 = (forvar857 + (1'h1)))
            begin
              reg858 = $signed(($signed((!$unsigned(reg799))) * $unsigned((~(reg854 ^~ reg840)))));
              reg859 <= (($unsigned(reg715[(4'hc):(3'h7)]) ?
                      reg844[(5'h13):(5'h12)] : $unsigned((reg838[(2'h3):(2'h3)] & reg801[(3'h4):(1'h1)]))) ?
                  $unsigned($signed((~^(forvar849 ?
                      wire704 : reg856)))) : $unsigned(reg838[(1'h0):(1'h0)]));
            end
          reg860 = {(reg715[(3'h5):(2'h2)] ?
                  {((reg819 ? reg795 : reg724) + $signed(reg799)),
                      $signed((reg761 & reg845)),
                      reg801} : (^$unsigned((reg831 ? wire708 : (7'h4a))))),
              $unsigned((~(7'h51))),
              reg720[(4'h9):(1'h0)]};
          reg861 = ($signed(reg837[(4'hb):(3'h4)]) ?
              $signed((~&($unsigned(reg715) ?
                  reg742[(1'h1):(1'h1)] : reg746[(2'h2):(1'h0)]))) : $unsigned($signed((reg724 > reg801))));
          for (forvar862 = (1'h0); (forvar862 < (1'h1)); forvar862 = (forvar862 + (1'h1)))
            begin
              reg863 <= $unsigned($signed({$unsigned((^reg840)),
                  (+$signed(reg836))}));
              reg864 = $signed(reg847[(4'h9):(3'h7)]);
            end
          reg865 = reg800[(2'h2):(2'h2)];
        end
      else
        begin
          reg857 = ($unsigned(($unsigned($signed(reg851)) ^ reg845)) ?
              reg848[(4'ha):(4'ha)] : ($signed(((reg846 & reg784) + (reg713 * reg828))) || (^reg848[(4'h8):(1'h1)])));
          for (forvar858 = (1'h0); (forvar858 < (1'h1)); forvar858 = (forvar858 + (1'h1)))
            begin
              reg859 <= reg846[(3'h4):(3'h4)];
              reg862 <= $signed($signed(reg791));
              reg864 = ((($unsigned(reg740[(4'hf):(4'h9)]) >= reg795[(4'hf):(4'h8)]) ?
                  $signed($signed((+(8'hb0)))) : $signed(reg775)) >> ((((reg839 >= reg821) && reg750) == ((+forvar858) ?
                  ((7'h52) >>> (8'ha1)) : $unsigned(reg726))) * (8'hbd)));
              reg865 = $unsigned($unsigned((7'h53)));
              reg866 = $signed(({(-$signed(reg768))} ?
                  (reg855 + (reg795 ?
                      reg842[(3'h7):(2'h3)] : $signed(reg740))) : reg768[(4'he):(1'h0)]));
            end
          for (forvar867 = (1'h0); (forvar867 < (1'h0)); forvar867 = (forvar867 + (1'h1)))
            begin
              reg868 <= (~|($unsigned($unsigned((+reg852))) && reg831[(3'h6):(3'h5)]));
              reg869 <= $unsigned(reg833[(5'h18):(4'hc)]);
              reg870 <= (reg851[(3'h6):(1'h1)] ?
                  ((7'h44) == ((~$unsigned(forvar862)) ?
                      (reg821 ? (~|reg720) : $unsigned(reg784)) : (reg852 ?
                          (reg801 & forvar829) : $signed(reg836)))) : $signed({$unsigned($signed(reg777)),
                      reg720,
                      reg856}));
              reg871 = (reg820[(4'h8):(1'h1)] ?
                  ((reg746 ? reg831 : reg855) ?
                      {$unsigned(reg713[(4'h9):(4'h8)]),
                          ({(8'hb9), reg808} ?
                              {reg724} : $unsigned(forvar867))} : reg720[(4'hb):(4'h9)]) : ($unsigned(((reg766 != wire705) ^~ {reg863,
                          reg777,
                          reg846})) ?
                      reg759[(1'h1):(1'h0)] : (((!reg756) ?
                              forvar858[(2'h2):(1'h1)] : reg713) ?
                          $signed(reg738[(5'h19):(5'h10)]) : (8'hb1))));
            end
          if ({$unsigned((((reg775 ? reg842 : (7'h46)) ?
                  {reg720} : (reg824 ? reg768 : reg855)) - {$signed(forvar867),
                  $unsigned(reg802),
                  reg808[(5'h1a):(5'h13)]}))})
            begin
              reg872 <= $unsigned(($signed((~^(reg837 ?
                  reg800 : reg791))) >= reg863));
            end
          else
            begin
              reg873 = (+(^(^~$signed(reg746[(1'h0):(1'h0)]))));
              reg874 <= reg838[(1'h1):(1'h0)];
              reg875 <= $unsigned(reg814);
              reg876 = $signed($signed($signed(({reg732} ?
                  $unsigned(forvar834) : $signed(wire705)))));
              reg877 <= reg845[(1'h0):(1'h0)];
            end
          reg878 <= $unsigned(reg770[(4'hd):(4'hc)]);
          for (forvar879 = (1'h0); (forvar879 < (3'h4)); forvar879 = (forvar879 + (1'h1)))
            begin
              reg880 <= reg797[(5'h12):(4'h9)];
              reg881 <= reg715[(3'h4):(2'h2)];
            end
        end
      if ((((reg769 << {(forvar858 | reg858)}) ~^ reg756) ?
          $signed(($signed({(7'h58)}) || ((|reg838) ?
              (reg836 * reg864) : reg759[(2'h2):(1'h1)]))) : $signed((~|$signed((^~wire707))))))
        begin
          reg882 = (((~^reg746) ?
                  (({(8'h9c), reg849} ?
                          $signed(reg843) : (reg795 ? reg877 : (7'h56))) ?
                      (!$unsigned((7'h56))) : $signed(reg856[(5'h10):(4'he)])) : (|$unsigned((8'hb1)))) ?
              (~|wire709) : reg841[(1'h0):(1'h0)]);
          reg883 = $unsigned(($unsigned(($signed(reg773) | reg749[(2'h2):(2'h2)])) & (~^reg724[(1'h0):(1'h0)])));
          if ($signed($unsigned(($signed((reg869 ? reg828 : reg759)) ?
              reg870 : $unsigned((~&reg848))))))
            begin
              reg884 = reg845;
              reg885 <= $signed($signed($unsigned(reg860[(3'h6):(1'h0)])));
              reg886 <= (!$signed((~^((reg724 ?
                  wire703 : reg773) >> {reg737}))));
              reg887 <= reg862;
              reg888 = $signed((~^(~^reg855)));
              reg889 = reg845[(5'h12):(4'hb)];
              reg890 = (-reg807[(3'h6):(3'h6)]);
            end
          else
            begin
              reg885 <= ({reg799[(3'h7):(1'h1)],
                      (~^(~^{reg833})),
                      reg801[(2'h2):(2'h2)]} ?
                  reg720 : {reg799, $signed(reg784[(5'h16):(4'hc)])});
              reg888 = reg773[(5'h18):(3'h7)];
              reg889 = ($signed(($signed(((7'h4c) ? reg861 : reg791)) ?
                  reg801 : reg777[(3'h4):(1'h1)])) < forvar849[(3'h7):(3'h4)]);
              reg891 <= $unsigned(reg877[(2'h2):(1'h1)]);
            end
          reg892 <= reg854;
          if (($signed($unsigned($signed((8'haf)))) >= $signed($unsigned({(&reg821)}))))
            begin
              reg893 = ((^~reg820) ?
                  ((7'h40) < (&reg715)) : (~|{reg886, $signed((^~reg873))}));
              reg894 <= (($unsigned($signed(reg884[(1'h0):(1'h0)])) ?
                      reg888[(1'h0):(1'h0)] : $unsigned(($unsigned(reg801) != $unsigned(reg766)))) ?
                  ((wire709[(2'h3):(2'h3)] < $unsigned((-reg887))) ^ {$unsigned(reg855),
                      reg714[(2'h2):(2'h2)],
                      reg755[(5'h10):(3'h4)]}) : $unsigned((($signed(reg768) && {reg726,
                          reg770}) ?
                      {reg864[(4'h8):(3'h7)],
                          $signed(reg738),
                          reg846[(4'he):(3'h6)]} : reg716[(2'h3):(2'h2)])));
              reg895 = reg750;
              reg896 = (~&(&reg746));
              reg897 = (reg777 ~^ (reg847[(2'h2):(2'h2)] ? reg713 : reg870));
            end
          else
            begin
              reg894 <= (&(8'h9e));
              reg898 <= reg838[(2'h2):(2'h2)];
              reg899 = forvar834[(3'h7):(1'h0)];
              reg900 <= reg884;
              reg901 <= ((~&$unsigned($unsigned($unsigned((8'hb3))))) ?
                  reg733 : {$unsigned($signed(reg797[(3'h4):(3'h4)])),
                      {(~(8'hb2)),
                          ((reg877 & forvar862) ?
                              ((7'h42) ? reg883 : reg836) : {wire704,
                                  (8'h9f),
                                  forvar862}),
                          reg838[(2'h3):(1'h0)]}});
            end
          if (reg854[(2'h2):(1'h1)])
            begin
              reg902 = reg833[(2'h2):(2'h2)];
              reg903 <= (~|reg819);
              reg904 = reg843[(3'h7):(3'h4)];
              reg905 <= reg860;
              reg906 = wire704;
              reg907 <= ((wire708[(1'h1):(1'h1)] ?
                      (reg897[(2'h2):(2'h2)] ?
                          (|$unsigned(reg900)) : ($signed((8'ha2)) || $unsigned(reg810))) : {($signed(reg824) == wire708[(2'h3):(2'h2)])}) ?
                  (($signed((wire825 >>> reg810)) ^ $signed($signed(reg888))) ?
                      (($unsigned((8'ha5)) ^~ $unsigned(reg724)) & ($unsigned(reg733) ?
                          $unsigned(reg852) : {reg888,
                              forvar879})) : $unsigned(($signed(reg863) ?
                          (reg755 ?
                              wire705 : reg872) : (reg862 ~^ (7'h45))))) : (|{($signed(reg790) ?
                          (reg889 ? reg846 : reg898) : (reg847 < reg873)),
                      $unsigned($unsigned(reg905))}));
            end
          else
            begin
              reg903 <= (~|(reg885 ? reg840 : {reg749}));
              reg905 <= reg850;
              reg907 <= forvar829;
              reg908 <= $signed(reg776[(2'h2):(1'h1)]);
              reg909 <= ({{((reg905 >>> reg808) ^~ (reg894 ?
                          forvar857 : reg778)),
                      {(reg773 ~^ reg859),
                          $signed(reg750)}}} << (((reg892[(1'h0):(1'h0)] < (~^reg843)) ~^ reg897) ?
                  ((~(reg768 || reg859)) <<< ((|forvar879) ?
                      $signed(reg874) : (reg892 ?
                          reg902 : (8'haa)))) : (($signed(reg821) || $unsigned(reg752)) ?
                      wire709[(2'h2):(2'h2)] : ($unsigned(reg784) ?
                          forvar834[(4'ha):(3'h4)] : $unsigned(reg844)))));
            end
          for (forvar910 = (1'h0); (forvar910 < (3'h6)); forvar910 = (forvar910 + (1'h1)))
            begin
              reg911 <= {($unsigned(reg779) ?
                      $signed(reg836[(4'ha):(4'h9)]) : (reg900[(3'h7):(2'h3)] < ((&reg878) ?
                          {forvar849, reg801, reg875} : $signed(reg740)))),
                  (&reg885[(3'h5):(1'h1)])};
            end
        end
      else
        begin
          if (reg795[(4'hb):(3'h4)])
            begin
              reg885 <= (($unsigned(reg808[(3'h4):(2'h2)]) ^~ {(+(forvar849 ?
                      (8'ha7) : reg855))}) - (-reg716));
              reg888 = (($unsigned(($signed(forvar849) <= reg778[(3'h5):(1'h0)])) >= reg828[(4'he):(2'h3)]) ?
                  $unsigned(($signed(reg890[(4'hf):(3'h6)]) ?
                      reg824 : $unsigned(((8'ha1) && reg853)))) : ($signed((~reg740)) ^ reg894[(1'h1):(1'h1)]));
              reg889 = ((&$signed($signed($unsigned(reg847)))) ?
                  $unsigned(({(~wire709),
                      $unsigned(reg901)} | ($unsigned(reg852) ?
                      reg807 : $unsigned(forvar867)))) : (-reg854));
              reg890 = $unsigned({reg833[(5'h18):(3'h7)]});
              reg891 <= ({reg903,
                  $signed(((^~reg820) <= (~^reg905))),
                  (+{reg892[(2'h3):(1'h0)],
                      (!(7'h40))})} & wire825[(2'h3):(2'h2)]);
              reg893 = forvar910[(1'h1):(1'h1)];
            end
          else
            begin
              reg885 <= ((reg800[(1'h1):(1'h0)] > (~|(^~$signed(reg716)))) || $signed($unsigned(reg857[(4'hf):(2'h2)])));
              reg888 = $signed(reg878);
              reg889 = ($signed((~|reg835[(3'h7):(3'h6)])) ?
                  (((+reg877) ? reg908[(5'h14):(5'h14)] : $unsigned(reg715)) ?
                      $unsigned(reg909[(3'h5):(2'h2)]) : ($signed($signed(reg716)) ?
                          $signed((reg890 ?
                              reg777 : reg756)) : (+(-reg724)))) : reg891[(3'h5):(2'h2)]);
              reg890 = (((!(reg909[(3'h7):(1'h1)] < reg715[(3'h4):(1'h0)])) ?
                      $signed((~^(reg773 ?
                          reg881 : reg887))) : (^~($unsigned(reg749) >= $unsigned(reg904)))) ?
                  $signed(reg846) : ({((^reg908) ?
                              ((8'h9c) ? forvar857 : wire709) : {reg800,
                                  reg835,
                                  reg872}),
                          $signed($unsigned(reg830))} ?
                      reg874[(3'h7):(3'h4)] : (reg824[(3'h7):(3'h4)] ?
                          $unsigned(reg766[(2'h2):(1'h0)]) : (!(7'h53)))));
            end
          reg894 <= {$signed((&(|$signed((7'h4b))))),
              $unsigned(reg855),
              reg895};
          for (forvar895 = (1'h0); (forvar895 < (2'h3)); forvar895 = (forvar895 + (1'h1)))
            begin
              reg898 <= $unsigned(reg884[(5'h12):(1'h0)]);
              reg900 <= reg907;
              reg901 <= (8'ha5);
              reg903 <= (reg830 <<< (8'ha6));
              reg905 <= $signed(reg797);
              reg907 <= (reg880[(1'h1):(1'h1)] ?
                  reg899[(3'h7):(2'h3)] : reg904[(2'h2):(2'h2)]);
              reg910 = (~|($unsigned((7'h44)) ?
                  reg838 : (((reg756 == wire706) >>> $unsigned(reg855)) - $unsigned(reg738))));
            end
          reg912 = {$signed({($signed(reg894) - $unsigned(reg892)),
                  $unsigned((|(8'ha3)))}),
              $signed(reg909)};
          reg913 <= ({forvar826[(2'h3):(1'h1)],
              $signed(reg819[(4'h8):(3'h6)]),
              reg842} | $unsigned(({((8'h9f) ? (7'h40) : reg820)} ?
              reg901[(5'h12):(4'he)] : $unsigned((+reg849)))));
          if (({$signed(reg815[(3'h7):(3'h4)]),
                  $signed(reg841[(1'h0):(1'h0)]),
                  reg827[(2'h2):(2'h2)]} ?
              reg809 : $unsigned(reg857[(2'h3):(2'h2)])))
            begin
              reg914 = reg860;
              reg915 = ($signed($unsigned($signed($signed(reg715)))) * $signed((!reg907[(3'h4):(1'h0)])));
              reg916 = ($signed((~^reg737)) * (reg815[(3'h4):(1'h0)] - {reg892,
                  ((-forvar829) + (forvar879 ? reg756 : reg833)),
                  (wire703 ? reg809 : (reg843 ? reg819 : reg756))}));
              reg917 = wire706[(5'h12):(5'h10)];
              reg918 = (^~(!reg835));
              reg919 <= ($unsigned((reg750[(1'h0):(1'h0)] ?
                  $unsigned($signed((7'h4b))) : $unsigned((reg775 ?
                      reg770 : reg891)))) ~^ (~|$signed(((reg821 >>> reg726) ?
                  {(7'h45)} : (reg766 ? reg884 : (8'hb7))))));
            end
          else
            begin
              reg919 <= ($signed($unsigned($unsigned((-reg894)))) << (reg801 ^~ (!reg880[(1'h0):(1'h0)])));
            end
          reg920 = {$signed(forvar895[(4'hf):(3'h7)])};
        end
      for (forvar921 = (1'h0); (forvar921 < (2'h2)); forvar921 = (forvar921 + (1'h1)))
        begin
          if (reg824[(4'hb):(3'h4)])
            begin
              reg922 = ((~{reg913,
                  (((8'hbd) ?
                      reg887 : forvar895) >= reg860[(4'he):(2'h2)])}) == $unsigned(($signed((reg773 ?
                  reg910 : reg770)) << reg883[(4'ha):(4'h8)])));
            end
          else
            begin
              reg922 = $unsigned($signed($unsigned(((forvar910 ?
                  reg759 : reg878) != (wire825 ? reg824 : reg898)))));
              reg923 <= (reg922[(1'h1):(1'h0)] << reg903);
              reg924 = (($signed((~^reg901)) ?
                      (reg892[(4'hc):(4'ha)] ?
                          (-(~wire703)) : reg885) : reg912[(1'h0):(1'h0)]) ?
                  (8'hb6) : {$unsigned(($signed(forvar826) != forvar862[(3'h5):(3'h4)]))});
              reg925 <= reg779;
              reg926 <= reg838[(1'h1):(1'h0)];
              reg927 = ($unsigned((forvar829[(1'h0):(1'h0)] - ($unsigned(reg913) >> reg860[(2'h3):(1'h0)]))) ?
                  (8'ha2) : $unsigned((+(~^reg741))));
            end
        end
      if ((^reg849))
        begin
          for (forvar928 = (1'h0); (forvar928 < (3'h6)); forvar928 = (forvar928 + (1'h1)))
            begin
              reg929 <= {reg853};
              reg930 <= reg733[(1'h1):(1'h1)];
              reg931 = {reg870[(5'h10):(4'he)]};
              reg932 <= (!({((8'ha4) << wire705[(3'h6):(1'h0)])} != {$signed(reg899),
                  (&$unsigned((8'ha3))),
                  $signed((-(8'hbc)))}));
              reg933 <= $unsigned($signed((-{reg800[(2'h3):(1'h1)]})));
            end
          reg934 <= (((~&reg810[(4'hf):(3'h6)]) ?
                  ($unsigned(reg925) << reg810) : reg918) ?
              ({($unsigned(reg887) << reg882[(4'he):(4'h8)]),
                      {((8'h9c) ? reg874 : reg807),
                          (forvar826 ? reg909 : reg881)}} ?
                  $unsigned($signed($signed(reg841))) : $unsigned(({(8'hb8),
                          reg827,
                          wire707} ?
                      reg889 : ((7'h40) - forvar858)))) : ((({reg931,
                          reg821,
                          reg831} ?
                      $unsigned(reg769) : (reg831 ?
                          reg819 : reg740)) ^ reg916[(1'h0):(1'h0)]) ?
                  $signed(((reg832 ^ reg924) ?
                      reg904[(5'h10):(4'hf)] : reg861)) : reg797));
        end
      else
        begin
          reg928 <= $unsigned((({reg875} ?
              (|$unsigned(forvar862)) : reg895) << $unsigned(($signed(reg824) || $signed(reg768)))));
          reg929 <= (&$unsigned($signed((reg904 || (reg741 ?
              forvar858 : reg801)))));
          reg930 <= $signed($signed(({(+reg899), $unsigned(reg899)} ?
              wire705 : $signed((reg928 ~^ reg872)))));
          reg932 <= reg776;
          reg935 = ($unsigned(reg871[(4'h8):(3'h6)]) && reg844[(4'hd):(1'h0)]);
          for (forvar936 = (1'h0); (forvar936 < (3'h6)); forvar936 = (forvar936 + (1'h1)))
            begin
              reg937 = $signed($signed((($signed(reg880) > (!reg871)) ^ (!reg747[(2'h3):(2'h2)]))));
              reg938 <= (+$unsigned(({(|reg923)} ~^ ({reg914} ?
                  ((8'ha5) ^~ reg926) : reg832))));
              reg939 = reg922;
              reg940 = $signed({(|{(reg815 ? reg863 : reg939),
                      (reg778 | reg911),
                      $unsigned(reg884)})});
              reg941 <= ((reg755 ?
                      $signed(((~|reg855) ?
                          (reg933 ? (8'hbb) : reg737) : (reg885 ?
                              (8'hbf) : reg836))) : $unsigned(reg755)) ?
                  wire704[(3'h5):(1'h0)] : {({reg880[(4'h8):(3'h5)],
                          reg841[(1'h0):(1'h0)],
                          reg831} + ((reg809 >= reg784) & reg750))});
              reg942 = (($unsigned($signed(reg724)) ?
                  reg853 : ((7'h40) ?
                      reg902[(5'h1a):(5'h16)] : $unsigned($signed(reg761)))) < $unsigned({(reg799[(4'h8):(3'h6)] ?
                      reg738[(5'h10):(3'h4)] : reg885),
                  $signed((reg754 ? reg918 : reg881)),
                  reg837[(2'h3):(2'h3)]}));
              reg943 <= (~^({reg893[(3'h4):(2'h2)], (|((7'h43) >= reg872))} ?
                  ((~|(~^(7'h4d))) ?
                      $signed((reg854 ?
                          forvar879 : forvar895)) : reg713[(4'h8):(2'h3)]) : {reg933[(3'h4):(1'h0)]}));
            end
        end
      for (forvar944 = (1'h0); (forvar944 < (3'h4)); forvar944 = (forvar944 + (1'h1)))
        begin
          if (reg912)
            begin
              reg945 = reg894[(1'h0):(1'h0)];
              reg946 = $signed((reg913[(3'h7):(3'h5)] + (8'hb1)));
              reg947 = $unsigned(reg900);
              reg948 <= $unsigned($signed(((&{forvar921,
                  reg930,
                  reg853}) == $signed($unsigned(reg742)))));
            end
          else
            begin
              reg945 = $signed({$signed((^wire707)), forvar826});
              reg946 = ((((~(8'ha7)) ?
                          forvar834 : (reg835[(4'h8):(3'h6)] > forvar928[(3'h4):(1'h1)])) ?
                      $unsigned(((-(7'h4f)) ?
                          (reg853 + reg768) : reg776)) : reg750) ?
                  (reg899[(3'h7):(1'h1)] ?
                      reg755[(4'hd):(1'h0)] : reg874[(3'h6):(1'h0)]) : reg898[(4'hf):(4'h8)]);
            end
          reg949 = reg831[(2'h2):(2'h2)];
          reg950 <= (~|wire703);
          reg951 = (~^((&$unsigned((reg752 ?
              (7'h48) : reg903))) <<< {(forvar857 ^~ $signed((8'hb9))),
              (reg891[(3'h5):(1'h1)] ? {forvar895} : (reg897 >>> (8'hbe)))}));
        end
    end
  always
    @(posedge clk) begin
      for (forvar952 = (1'h0); (forvar952 < (3'h6)); forvar952 = (forvar952 + (1'h1)))
        begin
          reg953 = (^~{(((~|reg775) ~^ (reg838 <= reg802)) ?
                  ($unsigned((8'hbf)) ?
                      (reg777 ? reg791 : reg737) : {reg930,
                          reg898,
                          reg819}) : reg747[(2'h3):(1'h0)]),
              {wire708,
                  $signed((reg800 - wire703)),
                  $signed((reg827 ? reg862 : reg713))},
              ((~^(^~reg737)) ?
                  $unsigned(((7'h4b) ^~ reg878)) : $signed((reg903 ?
                      reg737 : reg784)))});
          if ((^~reg759))
            begin
              reg954 <= ((^(($unsigned((7'h42)) ?
                      reg797[(5'h14):(4'h8)] : $signed(reg842)) ?
                  (reg755 <<< reg934) : (8'hb6))) == (^(reg820 >= reg754)));
            end
          else
            begin
              reg955 = $unsigned(reg859);
              reg956 <= (~|((reg911 == ($signed((8'haf)) ?
                      $unsigned(reg863) : $signed(reg862))) ?
                  ($unsigned((~^reg777)) ?
                      (reg854 || (wire704 ?
                          reg900 : reg846)) : $unsigned($unsigned(reg943))) : ($signed($unsigned((7'h4d))) ^ $unsigned((8'hae)))));
            end
          for (forvar957 = (1'h0); (forvar957 < (1'h0)); forvar957 = (forvar957 + (1'h1)))
            begin
              reg958 = (+(+reg732[(5'h1b):(4'hb)]));
              reg959 = reg795[(4'he):(3'h6)];
              reg960 = $signed((~|reg929[(4'hf):(1'h1)]));
              reg961 <= reg815;
              reg962 <= ((~&reg810[(5'h13):(5'h11)]) ?
                  (reg749 ? reg752 : (^(~&(^~reg742)))) : wire705);
              reg963 = {reg909[(1'h0):(1'h0)], reg953[(1'h0):(1'h0)]};
              reg964 = (($unsigned(((reg773 | reg886) && reg746[(1'h1):(1'h1)])) ?
                      (((7'h56) ? $signed(reg862) : $signed(reg713)) ?
                          $unsigned(reg752[(2'h2):(2'h2)]) : $unsigned((reg900 ?
                              reg880 : reg802))) : (reg752[(2'h2):(1'h1)] ?
                          (8'hb5) : reg740)) ?
                  $signed(reg715) : ((((reg752 << reg869) ?
                      {reg766,
                          reg862} : $signed((8'hbb))) > reg773) ~^ (-forvar952)));
            end
          reg965 <= reg740[(1'h0):(1'h0)];
        end
      reg966 = {((((reg911 ? reg815 : reg770) ? (~^reg891) : reg891) ?
              $unsigned({reg859, reg881, (7'h44)}) : {{wire706, reg716},
                  reg863[(5'h1d):(4'h9)]}) >= ((reg726[(4'hd):(4'h8)] ?
                  reg752 : (reg965 ? reg909 : reg849)) ?
              reg961 : ({reg801, (7'h57), reg901} ?
                  (+forvar952) : (~^reg800))))};
      if ((7'h4a))
        begin
          for (forvar967 = (1'h0); (forvar967 < (3'h5)); forvar967 = (forvar967 + (1'h1)))
            begin
              reg968 = ({{reg814, (reg801 ? reg726 : reg807[(4'hf):(4'hd)])}} ?
                  $signed((((reg815 ? reg943 : reg894) * reg740) && (^~(reg777 ?
                      reg841 : forvar957)))) : reg814[(3'h5):(3'h5)]);
              reg969 <= (($signed((+(wire703 <<< (8'hbe)))) >> $unsigned($unsigned($signed((7'h4d))))) & (reg875[(4'hb):(3'h5)] ?
                  $unsigned(((reg732 * reg821) || (reg784 != reg750))) : (reg808 ?
                      reg755[(4'he):(4'hd)] : (((8'ha8) == reg761) < (reg766 ?
                          (7'h54) : reg799)))));
              reg970 = {reg925[(2'h3):(1'h0)]};
              reg971 = reg898;
              reg972 <= ((^reg759) ? reg749[(1'h1):(1'h0)] : reg754);
              reg973 = $signed($unsigned({((8'haf) >= wire707),
                  ($unsigned(reg950) ? $unsigned(reg885) : $signed(reg797)),
                  $unsigned(reg908)}));
              reg974 <= (((^$signed(reg750[(3'h6):(3'h6)])) + $signed((!{(8'ha9),
                  reg930}))) ^~ (($unsigned($signed(reg775)) ?
                      $unsigned(reg964[(5'h10):(1'h1)]) : reg746[(1'h0):(1'h0)]) ?
                  {reg933[(1'h0):(1'h0)],
                      reg790[(2'h3):(2'h3)],
                      (~^$signed(reg724))} : reg925[(1'h1):(1'h0)]));
            end
          for (forvar975 = (1'h0); (forvar975 < (3'h5)); forvar975 = (forvar975 + (1'h1)))
            begin
              reg976 <= reg720[(5'h1b):(4'hb)];
              reg977 = reg732[(5'h17):(3'h7)];
              reg978 <= $unsigned({$signed(((reg778 ?
                      reg746 : reg943) >> $unsigned(reg953))),
                  ($signed((reg964 ~^ reg836)) != $signed($signed(reg737)))});
              reg979 <= {(((^~$unsigned((7'h40))) ?
                      ({reg859, reg726, wire707} ?
                          (-reg930) : (reg741 ?
                              reg819 : reg928)) : $signed($signed(reg777))) == $unsigned((~^$signed(wire707))))};
              reg980 = reg859;
            end
          if (reg824)
            begin
              reg981 = $signed({wire704[(1'h1):(1'h0)],
                  ((reg738[(5'h19):(4'h8)] ?
                      (reg769 >= wire705) : $signed(reg887)) >= ({reg964,
                          wire709} ?
                      (reg854 ? reg870 : reg954) : reg814))});
              reg982 <= reg715;
              reg983 <= (((reg776 ?
                          ((reg982 ?
                              reg740 : reg877) << (reg824 ^~ (7'h4c))) : $signed(reg907)) ?
                      $signed($signed($signed(reg800))) : ($unsigned((&reg875)) != ((+(8'h9d)) << reg842))) ?
                  reg752[(2'h2):(2'h2)] : ((&((|(7'h4b)) + wire709)) ?
                      $unsigned($signed((+reg956))) : (reg797 - $unsigned((reg982 & forvar957)))));
              reg984 <= reg969;
              reg985 <= wire708[(2'h3):(2'h3)];
              reg986 = ($signed(reg934[(4'hd):(3'h5)]) & ((reg892 ~^ $signed(reg872[(1'h1):(1'h1)])) ?
                  reg943[(1'h0):(1'h0)] : $signed(reg756[(5'h14):(4'h8)])));
              reg987 = (~^((reg955[(2'h3):(2'h3)] ?
                      reg842[(3'h5):(2'h3)] : ($unsigned(reg961) + $unsigned(forvar957))) ?
                  (reg885 ?
                      $unsigned((reg901 | reg973)) : reg715[(4'h8):(3'h5)]) : $unsigned((reg953[(1'h1):(1'h0)] ?
                      reg752[(2'h2):(1'h1)] : (|reg972)))));
            end
          else
            begin
              reg982 <= (wire706[(2'h2):(1'h0)] >= (7'h52));
              reg986 = $unsigned($unsigned((({reg720} ^ reg754[(3'h7):(1'h0)]) != reg720)));
            end
          for (forvar988 = (1'h0); (forvar988 < (1'h0)); forvar988 = (forvar988 + (1'h1)))
            begin
              reg989 = $unsigned({((~(reg901 & (8'ha2))) <<< reg941),
                  reg892[(4'hb):(3'h4)],
                  reg963[(1'h0):(1'h0)]});
              reg990 = ({reg973[(4'h8):(3'h6)],
                  ((-(reg863 ? reg877 : reg872)) ?
                      reg859 : {reg800,
                          (reg770 >= reg913)})} ^~ (^$unsigned(((8'hbf) ?
                  {reg976, reg756} : $signed(reg713)))));
              reg991 = wire704;
            end
          for (forvar992 = (1'h0); (forvar992 < (1'h1)); forvar992 = (forvar992 + (1'h1)))
            begin
              reg993 = (!($unsigned({$signed(reg932),
                      $unsigned(reg820),
                      reg832[(3'h5):(1'h1)]}) ?
                  ({reg810, (reg815 + reg877), (+reg870)} ?
                      ((reg755 ?
                          reg909 : reg715) || (8'ha8)) : (~reg769)) : ((~&(-reg738)) && $signed((^~reg863)))));
              reg994 <= {$unsigned($unsigned($signed($unsigned(reg894))))};
              reg995 = $signed((~|(($signed(reg981) ?
                  (reg990 && reg732) : reg950[(3'h6):(3'h5)]) != $signed((reg715 && reg979)))));
              reg996 = $signed((reg833[(1'h1):(1'h1)] ?
                  $signed($unsigned(reg926)) : $signed((((7'h48) ?
                      reg971 : reg881) == $unsigned(reg854)))));
              reg997 = (~$unsigned((((wire709 ? reg971 : (8'hb8)) != (reg872 ?
                      reg815 : (7'h4b))) ?
                  (!{reg779}) : (!((8'ha3) ? reg881 : reg933)))));
              reg998 <= $signed(reg832);
            end
          if ((reg891 ^~ {(|(!reg807[(4'he):(4'hd)])),
              ($signed(reg800[(2'h2):(1'h0)]) ?
                  forvar975[(4'hb):(1'h0)] : reg982[(4'hb):(2'h2)]),
              ((reg981 ? reg877[(3'h4):(2'h2)] : (+reg779)) ?
                  reg926[(5'h15):(4'h9)] : $unsigned(reg795[(1'h0):(1'h0)]))}))
            begin
              reg999 = reg778;
              reg1000 <= (reg832 & ({reg933, reg997[(2'h2):(2'h2)]} ?
                  $unsigned((reg986 ?
                      (^(8'hba)) : (forvar975 ?
                          reg886 : reg849))) : {$unsigned((reg775 <<< (7'h55))),
                      $signed({reg713, reg824})}));
            end
          else
            begin
              reg1000 <= (($unsigned(({(8'hb1),
                  reg980,
                  reg732} ^~ (~^(8'hbc)))) <= {({reg840, reg715} ?
                      (reg885 ? reg928 : forvar975) : (!reg994)),
                  $unsigned(((7'h48) >> (8'hae))),
                  $unsigned((reg819 | wire708))}) ^~ (!reg870[(5'h11):(1'h1)]));
              reg1001 = (reg855 * (&$signed((~|((7'h41) && reg963)))));
              reg1002 = (reg869 ?
                  (^~{$unsigned(reg885[(2'h3):(1'h1)]),
                      $signed((wire705 ~^ wire709))}) : (~$signed((-{reg973,
                      reg968}))));
              reg1003 <= $unsigned({$signed($unsigned($signed(reg737)))});
              reg1004 <= $signed($signed(reg887[(5'h11):(1'h1)]));
            end
        end
      else
        begin
          for (forvar967 = (1'h0); (forvar967 < (3'h6)); forvar967 = (forvar967 + (1'h1)))
            begin
              reg968 = {$unsigned($signed($signed((reg838 ?
                      reg913 : reg960))))};
              reg969 <= $signed($signed($signed(reg965)));
              reg970 = $unsigned($unsigned($signed($signed((reg909 <= reg960)))));
              reg972 <= reg875;
            end
          reg973 = $unsigned($signed(reg808));
        end
    end
  assign wire1005 = (|(!reg854[(2'h2):(1'h0)]));
  assign wire1006 = (wire705 ~^ reg754);
  assign wire1007 = $signed(wire705);
  always
    @(posedge clk) begin
      reg1008 = ($signed($unsigned($unsigned((^~reg726)))) >>> $signed(reg820));
      reg1009 <= $unsigned(reg827[(4'hc):(2'h2)]);
      reg1010 = (reg770 ?
          $unsigned((($unsigned(reg853) >> (reg752 ?
              reg726 : reg891)) << reg961)) : (($signed($unsigned((8'h9c))) ?
              $signed({reg740, reg737}) : (!((8'ha5) ?
                  reg872 : wire706))) ~^ $signed((^(reg773 != (8'ha5))))));
      reg1011 = $signed((($signed((+reg925)) >>> reg855[(4'h9):(3'h4)]) ?
          ((reg1000[(4'ha):(1'h0)] ? (~(7'h58)) : (~|reg750)) ?
              (|((8'hb8) == wire1007)) : $signed((-reg943))) : ($signed($unsigned((7'h47))) >= $unsigned((reg994 ?
              reg909 : reg928)))));
    end
  always
    @(posedge clk) begin
      for (forvar1012 = (1'h0); (forvar1012 < (1'h0)); forvar1012 = (forvar1012 + (1'h1)))
        begin
          if ((^~$unsigned($signed({(reg849 ? reg807 : reg797),
              ((7'h48) > wire707)}))))
            begin
              reg1013 <= ($signed($signed(reg819[(3'h7):(3'h6)])) ?
                  ((reg810 ?
                      ($signed((8'ha7)) >>> $signed(reg998)) : reg900[(4'hf):(1'h1)]) == $signed((^~(8'ha9)))) : (|reg827));
              reg1014 = $signed({reg1000[(3'h5):(2'h2)],
                  reg821[(5'h15):(1'h1)]});
              reg1015 <= (-$signed(reg815));
              reg1016 = (^~(8'hba));
              reg1017 = $signed({$signed($unsigned({reg726}))});
            end
          else
            begin
              reg1013 <= reg979;
              reg1015 <= ((((+(reg998 ? reg875 : reg901)) ?
                  (~$unsigned(reg950)) : (+$signed(reg929))) ^~ ((reg800 ?
                  $unsigned(reg878) : $signed(reg842)) == reg827)) || {reg948,
                  (~|reg741)});
              reg1016 = reg979[(4'h8):(1'h1)];
              reg1018 <= ($unsigned((~(7'h56))) ?
                  reg770 : (~&$signed($signed((-(8'hb6))))));
              reg1019 = $unsigned($unsigned((!reg948)));
              reg1020 <= (((wire705[(4'h9):(4'h8)] <= ($signed(reg911) ?
                      (reg801 ^~ reg819) : (reg713 ?
                          reg913 : wire1007))) < reg978) ?
                  (reg747[(3'h6):(3'h6)] ?
                      reg832[(1'h1):(1'h0)] : reg892[(5'h15):(4'he)]) : {(reg1013 ~^ (reg938[(4'he):(3'h6)] | ((8'ha9) != reg747)))});
            end
          if (reg819)
            begin
              reg1021 = $unsigned(reg930);
              reg1022 <= (!reg928[(4'hf):(3'h4)]);
              reg1023 <= (8'ha6);
              reg1024 <= (({$signed($signed(wire707)),
                      reg750,
                      reg974[(3'h7):(3'h5)]} > (~&reg827[(3'h6):(3'h4)])) ?
                  $unsigned(reg810[(5'h11):(1'h0)]) : ((7'h48) ?
                      (reg815 ?
                          $unsigned($signed(reg941)) : reg824[(3'h4):(3'h4)]) : {$signed(reg800),
                          ($unsigned((7'h4f)) >>> $unsigned(reg797))}));
            end
          else
            begin
              reg1021 = {reg919[(1'h1):(1'h0)],
                  reg892,
                  ($signed($signed($unsigned((7'h4d)))) ?
                      {$signed({(8'hbd), reg738}),
                          (~^reg875[(4'hc):(3'h7)])} : wire704[(1'h1):(1'h0)])};
              reg1022 <= reg962;
            end
          reg1025 <= $unsigned(wire1006);
          reg1026 <= $signed((reg976 ^~ $signed((8'ha8))));
          reg1027 = reg814;
        end
      for (forvar1028 = (1'h0); (forvar1028 < (3'h6)); forvar1028 = (forvar1028 + (1'h1)))
        begin
          if ({$unsigned((^($signed(reg840) ?
                  {reg983, reg815, reg994} : (^~reg923)))),
              $unsigned((((~reg713) ? (^~reg900) : (8'hb5)) ?
                  reg779[(5'h1b):(3'h7)] : $signed(reg1003[(3'h4):(2'h3)])))})
            begin
              reg1029 = (~|$signed(((reg713[(3'h4):(1'h1)] && (~|reg863)) != $signed({reg775,
                  reg880}))));
              reg1030 = $signed(reg849[(3'h6):(1'h1)]);
            end
          else
            begin
              reg1031 <= $signed((reg1009[(5'h15):(1'h1)] ?
                  (+reg790) : (reg720 ? reg777[(1'h0):(1'h0)] : (|reg969))));
              reg1032 = $signed(wire1007);
              reg1033 <= {((((reg901 || reg854) ?
                      $unsigned(reg815) : (reg878 == reg875)) >>> (~&$unsigned(reg738))) ^~ $signed(reg894[(1'h0):(1'h0)])),
                  (($signed($unsigned(reg930)) ^~ ((-reg985) & {reg1003,
                      reg911,
                      reg716})) > (reg720 * ($signed(reg869) ?
                      reg737 : reg820[(1'h0):(1'h0)])))};
              reg1034 <= $signed($unsigned(reg1026));
              reg1035 <= $unsigned(($unsigned(((7'h4d) ?
                  (reg1034 < (8'hb8)) : reg1014[(4'h8):(2'h2)])) << ((reg854[(2'h2):(1'h0)] ~^ (+reg907)) ?
                  reg1029[(3'h7):(3'h4)] : ($unsigned(reg1032) ?
                      {reg891} : (reg1019 ? reg854 : reg853)))));
            end
          for (forvar1036 = (1'h0); (forvar1036 < (3'h5)); forvar1036 = (forvar1036 + (1'h1)))
            begin
              reg1037 <= ((reg807[(2'h3):(2'h3)] + (^~$signed($signed(reg824)))) << ((+{(reg885 << reg994),
                      reg982,
                      reg907[(3'h6):(3'h5)]}) ?
                  (($unsigned((8'haa)) ^ {(7'h53), reg911, reg954}) ?
                      {(wire1006 + reg840)} : ($signed((8'ha3)) ?
                          (reg974 ?
                              reg907 : reg761) : (-reg784))) : reg819[(2'h2):(2'h2)]));
              reg1038 <= $signed((^~((~|{reg775, reg1015, reg833}) ?
                  reg901 : $signed($signed(reg724)))));
            end
          reg1039 <= (reg824 ? reg1029[(5'h12):(5'h10)] : (!reg842));
          for (forvar1040 = (1'h0); (forvar1040 < (3'h6)); forvar1040 = (forvar1040 + (1'h1)))
            begin
              reg1041 = (!(({$signed(reg892)} * ((~reg943) ?
                  {reg956,
                      reg755,
                      reg808} : (reg842 & reg928))) != (($signed(reg956) ^~ $unsigned(reg1026)) ?
                  (7'h43) : wire708)));
              reg1042 <= $signed((|reg1031));
              reg1043 <= (forvar1036[(4'h9):(4'h9)] ^~ reg903[(5'h14):(1'h1)]);
              reg1044 <= (8'hb8);
              reg1045 = (!reg1003[(3'h6):(3'h5)]);
              reg1046 = $signed(wire1007);
            end
        end
      for (forvar1047 = (1'h0); (forvar1047 < (3'h5)); forvar1047 = (forvar1047 + (1'h1)))
        begin
          reg1048 <= reg768[(4'hd):(4'hd)];
          for (forvar1049 = (1'h0); (forvar1049 < (2'h3)); forvar1049 = (forvar1049 + (1'h1)))
            begin
              reg1050 <= $signed((-($signed({reg862}) ?
                  reg872[(3'h5):(1'h0)] : ($signed(reg820) ?
                      (8'ha1) : {reg954}))));
              reg1051 = $unsigned(((reg784 ~^ $signed({(7'h55)})) ?
                  $signed(((reg976 ?
                      (8'ha0) : reg773) ^ (|reg737))) : (((reg776 ?
                      (8'hb2) : reg941) ^~ (reg887 + reg815)) <<< $signed($unsigned(reg797)))));
              reg1052 = ((|reg756[(4'ha):(2'h2)]) ?
                  ((8'h9d) <<< reg1046) : reg983);
              reg1053 <= $unsigned(((reg983 ?
                      reg985 : reg1050[(5'h1d):(5'h1a)]) ?
                  ($signed((reg1021 ?
                      forvar1028 : reg1026)) > {$unsigned(reg775),
                      reg824,
                      $unsigned(reg831)}) : ((reg841 ?
                          (reg732 || (8'h9f)) : (reg905 ? (7'h48) : reg1033)) ?
                      $signed((-reg950)) : $unsigned({(8'hb8), wire706}))));
              reg1054 = reg894;
              reg1055 <= $unsigned(reg1033);
              reg1056 <= reg868;
            end
        end
      for (forvar1057 = (1'h0); (forvar1057 < (1'h0)); forvar1057 = (forvar1057 + (1'h1)))
        begin
          for (forvar1058 = (1'h0); (forvar1058 < (2'h3)); forvar1058 = (forvar1058 + (1'h1)))
            begin
              reg1059 = $signed($signed($unsigned(reg1044[(1'h1):(1'h0)])));
              reg1060 <= $unsigned($signed($signed(((-reg868) ?
                  (reg1052 && reg749) : reg972))));
              reg1061 = reg749[(4'hb):(4'h9)];
              reg1062 = reg797[(4'he):(2'h2)];
              reg1063 = ($signed(reg1056) | ((({reg911, (8'hb9)} ?
                      (wire708 ?
                          reg831 : reg1045) : $signed(reg862)) & (&$signed(reg754))) ?
                  (reg1050 ?
                      ($unsigned(reg1060) ?
                          $unsigned(reg1055) : ((8'hbc) & reg799)) : (~|reg934)) : (~^(wire709 ?
                      (!reg979) : (~&reg969)))));
              reg1064 = $signed((|$unsigned((reg1042 > (8'hae)))));
              reg1065 = $signed($signed(($unsigned((reg750 >>> reg1045)) ?
                  {((7'h44) ? reg755 : reg1009),
                      reg934[(4'ha):(3'h4)]} : $unsigned(reg790))));
            end
          reg1066 = $unsigned(reg859[(2'h3):(2'h3)]);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1695  (y, clk, wire1699, wire1698, wire1697, wire1696);
  output wire [(32'h1525):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire1699;
  input wire signed [(5'h19):(1'h0)] wire1698;
  input wire [(5'h18):(1'h0)] wire1697;
  input wire signed [(3'h5):(1'h0)] wire1696;
  wire signed [(5'h16):(1'h0)] wire2892;
  wire signed [(5'h12):(1'h0)] wire2891;
  wire signed [(5'h12):(1'h0)] wire2890;
  wire signed [(5'h14):(1'h0)] wire2889;
  wire signed [(5'h1d):(1'h0)] wire2887;
  wire signed [(5'h18):(1'h0)] wire2876;
  wire [(4'he):(1'h0)] wire2864;
  wire signed [(4'h9):(1'h0)] wire2863;
  wire signed [(3'h4):(1'h0)] wire2823;
  wire signed [(5'h12):(1'h0)] wire2822;
  wire [(3'h7):(1'h0)] wire2821;
  wire [(3'h7):(1'h0)] wire2820;
  wire signed [(5'h1e):(1'h0)] wire2730;
  wire [(5'h1b):(1'h0)] wire2729;
  wire [(5'h11):(1'h0)] wire2728;
  wire signed [(5'h19):(1'h0)] wire2688;
  wire [(5'h1c):(1'h0)] wire2635;
  wire [(2'h3):(1'h0)] wire1725;
  wire [(5'h1e):(1'h0)] wire1724;
  wire [(5'h18):(1'h0)] wire1723;
  wire [(5'h15):(1'h0)] wire1722;
  reg [(5'h16):(1'h0)] reg2945 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2941 = (1'h0);
  reg [(5'h11):(1'h0)] reg2936 = (1'h0);
  reg [(4'hc):(1'h0)] reg2935 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2933 = (1'h0);
  reg [(4'h8):(1'h0)] reg2932 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2925 = (1'h0);
  reg [(4'ha):(1'h0)] reg2923 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2922 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2920 = (1'h0);
  reg [(5'h11):(1'h0)] reg2918 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2914 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2908 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2907 = (1'h0);
  reg [(3'h6):(1'h0)] reg2904 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2902 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2900 = (1'h0);
  reg [(4'hb):(1'h0)] reg1755 = (1'h0);
  reg [(4'hb):(1'h0)] reg1754 = (1'h0);
  reg [(5'h14):(1'h0)] reg1752 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1749 = (1'h0);
  reg [(5'h17):(1'h0)] reg1748 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1747 = (1'h0);
  reg [(4'hd):(1'h0)] reg1746 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1744 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1736 = (1'h0);
  reg [(5'h19):(1'h0)] reg1735 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1734 = (1'h0);
  reg [(3'h7):(1'h0)] reg1731 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1729 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1728 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1720 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1718 = (1'h0);
  reg [(3'h4):(1'h0)] reg1712 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1711 = (1'h0);
  reg [(5'h19):(1'h0)] reg1707 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1702 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1700 = (1'h0);
  reg [(5'h12):(1'h0)] reg2637 = (1'h0);
  reg [(3'h5):(1'h0)] reg2638 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2640 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2641 = (1'h0);
  reg [(3'h5):(1'h0)] reg2692 = (1'h0);
  reg [(5'h13):(1'h0)] reg2693 = (1'h0);
  reg [(3'h4):(1'h0)] reg2694 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2696 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2702 = (1'h0);
  reg [(4'hf):(1'h0)] reg2703 = (1'h0);
  reg [(4'he):(1'h0)] reg2705 = (1'h0);
  reg [(5'h10):(1'h0)] reg2707 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2708 = (1'h0);
  reg [(2'h3):(1'h0)] reg2711 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2713 = (1'h0);
  reg [(5'h14):(1'h0)] reg2719 = (1'h0);
  reg [(5'h15):(1'h0)] reg2725 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2726 = (1'h0);
  reg [(5'h11):(1'h0)] reg2731 = (1'h0);
  reg [(5'h15):(1'h0)] reg2734 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2735 = (1'h0);
  reg [(4'hb):(1'h0)] reg2736 = (1'h0);
  reg [(5'h11):(1'h0)] reg2737 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2740 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2741 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2742 = (1'h0);
  reg [(5'h14):(1'h0)] reg2743 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2746 = (1'h0);
  reg [(5'h14):(1'h0)] reg2747 = (1'h0);
  reg [(4'hf):(1'h0)] reg2749 = (1'h0);
  reg [(5'h17):(1'h0)] reg2751 = (1'h0);
  reg [(5'h11):(1'h0)] reg2752 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2753 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2758 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2759 = (1'h0);
  reg [(3'h5):(1'h0)] reg2762 = (1'h0);
  reg [(4'ha):(1'h0)] reg2765 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2766 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2768 = (1'h0);
  reg [(5'h15):(1'h0)] reg2772 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2773 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2776 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2784 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2789 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2791 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2795 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2799 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2803 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2804 = (1'h0);
  reg [(3'h6):(1'h0)] reg2806 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2807 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2809 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2810 = (1'h0);
  reg [(4'h8):(1'h0)] reg2811 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2813 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2814 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2815 = (1'h0);
  reg [(5'h12):(1'h0)] reg2817 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2824 = (1'h0);
  reg [(4'hb):(1'h0)] reg2827 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2828 = (1'h0);
  reg [(4'ha):(1'h0)] reg2831 = (1'h0);
  reg [(5'h12):(1'h0)] reg2835 = (1'h0);
  reg [(2'h3):(1'h0)] reg2836 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2841 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2843 = (1'h0);
  reg [(5'h15):(1'h0)] reg2845 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2850 = (1'h0);
  reg [(5'h15):(1'h0)] reg2851 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2853 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2854 = (1'h0);
  reg [(4'hc):(1'h0)] reg2856 = (1'h0);
  reg [(5'h14):(1'h0)] reg2859 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2860 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2861 = (1'h0);
  reg [(3'h6):(1'h0)] reg2866 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2871 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2872 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2873 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2875 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2944 = (1'h0);
  reg [(3'h5):(1'h0)] reg2943 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2942 = (1'h0);
  reg [(3'h4):(1'h0)] reg2940 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2939 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2938 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2937 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2930 = (1'h0);
  reg [(5'h15):(1'h0)] reg2934 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2931 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2930 = (1'h0);
  reg [(2'h3):(1'h0)] reg2929 = (1'h0);
  reg [(4'he):(1'h0)] reg2928 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2927 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2926 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2924 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2921 = (1'h0);
  reg [(2'h3):(1'h0)] reg2919 = (1'h0);
  reg [(2'h2):(1'h0)] reg2917 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2916 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2915 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2913 = (1'h0);
  reg [(5'h13):(1'h0)] reg2912 = (1'h0);
  reg [(2'h2):(1'h0)] reg2911 = (1'h0);
  reg [(2'h3):(1'h0)] reg2910 = (1'h0);
  reg [(2'h2):(1'h0)] reg2909 = (1'h0);
  reg [(5'h19):(1'h0)] reg2906 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2905 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2903 = (1'h0);
  reg [(5'h12):(1'h0)] reg2901 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2899 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2898 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2897 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2896 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2895 = (1'h0);
  reg [(4'ha):(1'h0)] reg2894 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2893 = (1'h0);
  reg [(5'h13):(1'h0)] reg2874 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2870 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2869 = (1'h0);
  reg [(2'h2):(1'h0)] reg2868 = (1'h0);
  reg [(5'h19):(1'h0)] reg2867 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2865 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2862 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2858 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2857 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2855 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2852 = (1'h0);
  reg [(4'hc):(1'h0)] reg2849 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2848 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2847 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2847 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2846 = (1'h0);
  reg [(5'h18):(1'h0)] reg2844 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar2838 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2842 = (1'h0);
  reg [(4'hc):(1'h0)] reg2840 = (1'h0);
  reg [(2'h3):(1'h0)] reg2839 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2838 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2837 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2834 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2833 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2832 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2830 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2829 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2826 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2825 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2819 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2818 = (1'h0);
  reg [(4'ha):(1'h0)] reg2816 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2813 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2809 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2812 = (1'h0);
  reg [(5'h13):(1'h0)] reg2808 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2805 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2802 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2801 = (1'h0);
  reg [(4'hb):(1'h0)] reg2800 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2798 = (1'h0);
  reg [(4'h9):(1'h0)] reg2797 = (1'h0);
  reg [(5'h14):(1'h0)] reg2796 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2794 = (1'h0);
  reg [(5'h17):(1'h0)] reg2793 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2792 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2790 = (1'h0);
  reg [(4'ha):(1'h0)] reg2788 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2787 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2786 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2785 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2783 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2782 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2781 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2780 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2779 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2778 = (1'h0);
  reg [(5'h11):(1'h0)] reg2777 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2775 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2774 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2771 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2770 = (1'h0);
  reg [(3'h4):(1'h0)] reg2769 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2767 = (1'h0);
  reg [(5'h15):(1'h0)] reg2764 = (1'h0);
  reg [(5'h10):(1'h0)] reg2763 = (1'h0);
  reg [(5'h12):(1'h0)] reg2761 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2760 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2757 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2756 = (1'h0);
  reg [(5'h16):(1'h0)] reg2755 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2754 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2750 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2748 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2745 = (1'h0);
  reg [(5'h13):(1'h0)] reg2744 = (1'h0);
  reg [(4'ha):(1'h0)] reg2739 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2738 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2733 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2732 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2727 = (1'h0);
  reg [(5'h1c):(1'h0)] forvar2724 = (1'h0);
  reg [(3'h4):(1'h0)] reg2723 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2722 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2721 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2720 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2718 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2717 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2716 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2715 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2714 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2712 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2710 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2709 = (1'h0);
  reg [(3'h4):(1'h0)] reg2706 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2704 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2701 = (1'h0);
  reg [(3'h5):(1'h0)] reg2700 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2699 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2698 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2697 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2695 = (1'h0);
  reg [(2'h3):(1'h0)] reg2691 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2690 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2643 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2642 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2639 = (1'h0);
  reg [(4'h9):(1'h0)] reg1758 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar1744 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1757 = (1'h0);
  reg [(3'h5):(1'h0)] reg1756 = (1'h0);
  reg [(5'h16):(1'h0)] reg1753 = (1'h0);
  reg [(5'h12):(1'h0)] reg1751 = (1'h0);
  reg [(5'h16):(1'h0)] reg1750 = (1'h0);
  reg [(4'hc):(1'h0)] reg1745 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1743 = (1'h0);
  reg [(5'h10):(1'h0)] reg1742 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1741 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1740 = (1'h0);
  reg [(5'h17):(1'h0)] reg1739 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1738 = (1'h0);
  reg [(4'hd):(1'h0)] reg1737 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1732 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1731 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1733 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1732 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1730 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1727 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1726 = (1'h0);
  reg [(2'h3):(1'h0)] reg1721 = (1'h0);
  reg [(4'ha):(1'h0)] reg1719 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1717 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1716 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1715 = (1'h0);
  reg [(5'h11):(1'h0)] reg1714 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1713 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1710 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1709 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1708 = (1'h0);
  reg [(5'h15):(1'h0)] reg1706 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1705 = (1'h0);
  reg [(4'h9):(1'h0)] reg1704 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1703 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1701 = (1'h0);
  assign y = {wire2892,
                 wire2891,
                 wire2890,
                 wire2889,
                 wire2887,
                 wire2876,
                 wire2864,
                 wire2863,
                 wire2823,
                 wire2822,
                 wire2821,
                 wire2820,
                 wire2730,
                 wire2729,
                 wire2728,
                 wire2688,
                 wire2635,
                 wire1725,
                 wire1724,
                 wire1723,
                 wire1722,
                 reg2945,
                 reg2941,
                 reg2936,
                 reg2935,
                 reg2933,
                 reg2932,
                 reg2925,
                 reg2923,
                 reg2922,
                 reg2920,
                 reg2918,
                 reg2914,
                 reg2908,
                 reg2907,
                 reg2904,
                 reg2902,
                 reg2900,
                 reg1755,
                 reg1754,
                 reg1752,
                 reg1749,
                 reg1748,
                 reg1747,
                 reg1746,
                 reg1744,
                 reg1736,
                 reg1735,
                 reg1734,
                 reg1731,
                 reg1729,
                 reg1728,
                 reg1720,
                 reg1718,
                 reg1712,
                 reg1711,
                 reg1707,
                 reg1702,
                 reg1700,
                 reg2637,
                 reg2638,
                 reg2640,
                 reg2641,
                 reg2692,
                 reg2693,
                 reg2694,
                 reg2696,
                 reg2702,
                 reg2703,
                 reg2705,
                 reg2707,
                 reg2708,
                 reg2711,
                 reg2713,
                 reg2719,
                 reg2725,
                 reg2726,
                 reg2731,
                 reg2734,
                 reg2735,
                 reg2736,
                 reg2737,
                 reg2740,
                 reg2741,
                 reg2742,
                 reg2743,
                 reg2746,
                 reg2747,
                 reg2749,
                 reg2751,
                 reg2752,
                 reg2753,
                 reg2758,
                 reg2759,
                 reg2762,
                 reg2765,
                 reg2766,
                 reg2768,
                 reg2772,
                 reg2773,
                 reg2776,
                 reg2784,
                 reg2789,
                 reg2791,
                 reg2795,
                 reg2799,
                 reg2803,
                 reg2804,
                 reg2806,
                 reg2807,
                 reg2809,
                 reg2810,
                 reg2811,
                 reg2813,
                 reg2814,
                 reg2815,
                 reg2817,
                 reg2824,
                 reg2827,
                 reg2828,
                 reg2831,
                 reg2835,
                 reg2836,
                 reg2841,
                 reg2843,
                 reg2845,
                 reg2850,
                 reg2851,
                 reg2853,
                 reg2854,
                 reg2856,
                 reg2859,
                 reg2860,
                 reg2861,
                 reg2866,
                 reg2871,
                 reg2872,
                 reg2873,
                 reg2875,
                 reg2944,
                 reg2943,
                 reg2942,
                 reg2940,
                 reg2939,
                 forvar2938,
                 forvar2937,
                 reg2930,
                 reg2934,
                 reg2931,
                 forvar2930,
                 reg2929,
                 reg2928,
                 reg2927,
                 reg2926,
                 forvar2924,
                 reg2921,
                 reg2919,
                 reg2917,
                 reg2916,
                 reg2915,
                 reg2913,
                 reg2912,
                 reg2911,
                 reg2910,
                 reg2909,
                 reg2906,
                 forvar2905,
                 reg2903,
                 reg2901,
                 reg2899,
                 reg2898,
                 forvar2897,
                 reg2896,
                 forvar2895,
                 reg2894,
                 reg2893,
                 reg2874,
                 reg2870,
                 reg2869,
                 reg2868,
                 reg2867,
                 forvar2865,
                 reg2862,
                 forvar2858,
                 reg2857,
                 reg2855,
                 reg2852,
                 reg2849,
                 reg2848,
                 forvar2847,
                 reg2847,
                 reg2846,
                 reg2844,
                 forvar2838,
                 reg2842,
                 reg2840,
                 reg2839,
                 reg2838,
                 reg2837,
                 reg2834,
                 reg2833,
                 reg2832,
                 reg2830,
                 reg2829,
                 forvar2826,
                 reg2825,
                 reg2819,
                 reg2818,
                 reg2816,
                 forvar2813,
                 forvar2809,
                 reg2812,
                 reg2808,
                 forvar2805,
                 forvar2802,
                 forvar2801,
                 reg2800,
                 reg2798,
                 reg2797,
                 reg2796,
                 reg2794,
                 reg2793,
                 reg2792,
                 forvar2790,
                 reg2788,
                 reg2787,
                 reg2786,
                 forvar2785,
                 reg2783,
                 reg2782,
                 reg2781,
                 reg2780,
                 forvar2779,
                 reg2778,
                 reg2777,
                 forvar2775,
                 forvar2774,
                 reg2771,
                 reg2770,
                 reg2769,
                 forvar2767,
                 reg2764,
                 reg2763,
                 reg2761,
                 forvar2760,
                 reg2757,
                 forvar2756,
                 reg2755,
                 reg2754,
                 reg2750,
                 reg2748,
                 reg2745,
                 reg2744,
                 reg2739,
                 forvar2738,
                 forvar2733,
                 reg2732,
                 reg2727,
                 forvar2724,
                 reg2723,
                 reg2722,
                 forvar2721,
                 reg2720,
                 reg2718,
                 forvar2717,
                 reg2716,
                 reg2715,
                 reg2714,
                 reg2712,
                 reg2710,
                 reg2709,
                 reg2706,
                 reg2704,
                 reg2701,
                 reg2700,
                 reg2699,
                 reg2698,
                 reg2697,
                 forvar2695,
                 reg2691,
                 forvar2690,
                 reg2643,
                 reg2642,
                 reg2639,
                 reg1758,
                 forvar1744,
                 reg1757,
                 reg1756,
                 reg1753,
                 reg1751,
                 reg1750,
                 reg1745,
                 reg1743,
                 reg1742,
                 reg1741,
                 reg1740,
                 reg1739,
                 reg1738,
                 reg1737,
                 reg1732,
                 forvar1731,
                 reg1733,
                 forvar1732,
                 reg1730,
                 reg1727,
                 reg1726,
                 reg1721,
                 reg1719,
                 reg1717,
                 reg1716,
                 forvar1715,
                 reg1714,
                 reg1713,
                 forvar1710,
                 reg1709,
                 forvar1708,
                 reg1706,
                 reg1705,
                 reg1704,
                 reg1703,
                 reg1701,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1700 <= $unsigned($unsigned($signed(((wire1696 ? wire1698 : wire1697) ?
          (+(7'h45)) : $signed(wire1699)))));
      reg1701 = ($signed($unsigned(reg1700[(5'h19):(5'h10)])) ?
          wire1697[(3'h6):(2'h2)] : ((^$signed(wire1696[(1'h1):(1'h0)])) ?
              reg1700[(1'h1):(1'h1)] : wire1698[(5'h13):(1'h0)]));
      if ((reg1701[(4'h9):(1'h1)] ?
          $unsigned(($unsigned($unsigned((8'ha0))) ?
              ($signed(reg1700) ?
                  reg1700[(3'h6):(1'h1)] : ((7'h4e) ?
                      reg1700 : (8'hba))) : {reg1700})) : wire1697[(5'h18):(1'h0)]))
        begin
          if ((^~reg1701[(4'h9):(3'h7)]))
            begin
              reg1702 <= (wire1696 > wire1698[(4'hf):(4'ha)]);
              reg1703 = $unsigned(({(-(wire1699 ? (7'h50) : reg1702)),
                  wire1698[(5'h13):(4'h9)]} != $signed(($unsigned(reg1702) ?
                  (-wire1697) : wire1698))));
              reg1704 = $unsigned((~^$unsigned(($signed(reg1702) && reg1700[(4'h8):(3'h7)]))));
              reg1705 = (reg1700 ?
                  ((reg1703 ?
                          ((wire1697 * reg1700) ~^ (wire1698 ^ reg1704)) : wire1699[(3'h7):(2'h2)]) ?
                      (+(~|(|wire1697))) : {reg1702,
                          reg1702[(3'h7):(2'h2)],
                          (7'h4c)}) : wire1697);
              reg1706 = (^(wire1699 ?
                  $unsigned($signed(reg1703[(5'h13):(5'h10)])) : (wire1696 ?
                      (reg1700 < ((8'haa) >>> reg1701)) : (!$unsigned(wire1698)))));
            end
          else
            begin
              reg1702 <= ((reg1705 >= $unsigned(((wire1698 <= (8'hb7)) == (wire1699 == reg1703)))) ?
                  {(reg1700 ? $unsigned((-(8'hac))) : (8'hba)),
                      reg1702[(4'hb):(2'h3)]} : $signed($signed($unsigned((wire1699 ?
                      reg1701 : reg1703)))));
            end
          reg1707 <= reg1706;
        end
      else
        begin
          reg1702 <= ((({$unsigned(reg1702),
                          (reg1703 ? (8'hb8) : wire1697),
                          (reg1707 >= (8'ha6))} ?
                      reg1700[(4'ha):(4'h8)] : (~{reg1703, (7'h46), reg1702})) ?
                  ({{reg1707, reg1704}, reg1707[(3'h7):(2'h3)]} ?
                      ($signed(reg1701) - {reg1706,
                          reg1704}) : ((reg1702 <<< (7'h55)) * (reg1701 ?
                          wire1696 : (8'hb6)))) : {({(8'hb6)} >= (&(8'h9e))),
                      $unsigned((reg1705 > wire1699)),
                      (~$unsigned(reg1701))}) ?
              $signed((((~wire1697) == (reg1701 ? (7'h58) : wire1699)) ?
                  $signed((reg1705 > reg1707)) : $signed($unsigned(reg1707)))) : $signed(($signed((7'h50)) << $signed((wire1697 ?
                  (8'ha2) : wire1697)))));
        end
      for (forvar1708 = (1'h0); (forvar1708 < (1'h0)); forvar1708 = (forvar1708 + (1'h1)))
        begin
          reg1709 = $unsigned(forvar1708);
          for (forvar1710 = (1'h0); (forvar1710 < (1'h0)); forvar1710 = (forvar1710 + (1'h1)))
            begin
              reg1711 <= $unsigned(wire1696[(2'h2):(2'h2)]);
              reg1712 <= ($unsigned($unsigned({(^wire1699)})) ?
                  $unsigned((7'h47)) : ($unsigned($signed((wire1697 < forvar1710))) || $signed(($unsigned(reg1705) + $signed(reg1706)))));
              reg1713 = $signed((^~(reg1711 ^ $unsigned($signed(reg1712)))));
              reg1714 = (reg1711[(3'h7):(3'h7)] ?
                  {forvar1708[(2'h2):(1'h0)]} : (7'h46));
            end
          for (forvar1715 = (1'h0); (forvar1715 < (1'h1)); forvar1715 = (forvar1715 + (1'h1)))
            begin
              reg1716 = (8'hbd);
              reg1717 = $unsigned($unsigned((+$signed(reg1704))));
              reg1718 <= $unsigned({reg1701, reg1705});
              reg1719 = $signed($signed($unsigned(forvar1715[(3'h7):(2'h3)])));
              reg1720 <= (^reg1712[(1'h1):(1'h0)]);
              reg1721 = ($unsigned($unsigned($unsigned(forvar1708))) ?
                  (reg1713[(2'h3):(2'h2)] ?
                      $unsigned($unsigned({wire1697,
                          reg1711,
                          reg1711})) : ($unsigned((~&(7'h50))) >> (reg1706 ?
                          forvar1710 : {reg1719,
                              reg1702}))) : {$unsigned((-$unsigned(forvar1715)))});
            end
        end
    end
  assign wire1722 = reg1700[(5'h17):(2'h2)];
  assign wire1723 = reg1700;
  assign wire1724 = ($unsigned($signed($signed((wire1696 ?
                            reg1720 : wire1698)))) ?
                        (8'ha7) : (reg1707 && wire1723[(1'h0):(1'h0)]));
  assign wire1725 = ((wire1697[(5'h13):(5'h11)] ?
                        wire1722 : wire1723[(3'h7):(2'h2)]) > ($unsigned($signed(reg1707[(4'hf):(3'h6)])) == {($signed(reg1711) ?
                            $unsigned(reg1700) : {reg1702, wire1723}),
                        reg1711[(4'ha):(4'ha)],
                        (~|((8'ha9) ? reg1702 : wire1696))}));
  always
    @(posedge clk) begin
      reg1726 = wire1723[(5'h18):(4'h9)];
      reg1727 = $signed({$unsigned(wire1725)});
      reg1728 <= ((reg1700[(4'hb):(4'hb)] ^~ $signed(({wire1698} == wire1699[(3'h6):(3'h5)]))) >= (wire1699 ~^ {(+(wire1696 ?
              wire1725 : reg1727)),
          ((~|wire1722) + $signed(wire1723))}));
    end
  always
    @(posedge clk) begin
      reg1729 <= wire1724[(4'hb):(2'h2)];
      reg1730 = $unsigned(wire1723[(5'h12):(4'hd)]);
      if ($signed(reg1718))
        begin
          reg1731 <= wire1725[(2'h2):(1'h0)];
          for (forvar1732 = (1'h0); (forvar1732 < (1'h0)); forvar1732 = (forvar1732 + (1'h1)))
            begin
              reg1733 = $signed($signed($unsigned($signed((reg1728 >>> (8'hbe))))));
              reg1734 <= ((-(reg1730[(2'h2):(2'h2)] ~^ {$signed(reg1720),
                      (wire1723 | (8'hba))})) ?
                  (8'ha4) : wire1697[(3'h4):(1'h0)]);
              reg1735 <= ($signed(({(~wire1724)} + wire1723)) ?
                  (+(8'ha7)) : (~^(7'h4c)));
              reg1736 <= $unsigned((7'h40));
            end
        end
      else
        begin
          for (forvar1731 = (1'h0); (forvar1731 < (2'h3)); forvar1731 = (forvar1731 + (1'h1)))
            begin
              reg1732 = ($signed(reg1729) && $unsigned(wire1724));
              reg1733 = wire1724[(5'h19):(1'h0)];
              reg1737 = (($unsigned(forvar1732) ?
                  $unsigned(((-forvar1731) ?
                      wire1723 : (~wire1725))) : $unsigned(reg1707[(5'h17):(5'h17)])) << ($unsigned({$unsigned(reg1734)}) ^ (+(8'hbe))));
              reg1738 = $signed(($unsigned((((7'h41) <= reg1718) ?
                      $unsigned((7'h4c)) : reg1720)) ?
                  ($unsigned($signed(wire1724)) & forvar1731) : (reg1731[(1'h1):(1'h0)] ?
                      $signed(wire1722) : ($signed(reg1737) ?
                          {reg1736} : ((8'hb8) ? (8'hab) : reg1729)))));
              reg1739 = $signed(((8'ha7) & wire1698));
              reg1740 = $signed($unsigned((|wire1697)));
              reg1741 = reg1733;
            end
        end
      reg1742 = {$signed((~|$signed((wire1697 ? (7'h46) : reg1741)))),
          {$unsigned($signed($unsigned(forvar1732)))},
          ($signed(reg1729[(3'h4):(2'h2)]) ~^ (8'hb9))};
      reg1743 = $unsigned($unsigned(wire1725[(2'h2):(1'h0)]));
      if ((!(({(wire1699 ? wire1697 : reg1728),
              $signed((8'haa))} ~^ $signed(wire1724)) ?
          $signed(reg1737[(3'h4):(3'h4)]) : $signed(((~^reg1720) != reg1738)))))
        begin
          reg1744 <= $signed(reg1707[(5'h16):(4'h8)]);
          reg1745 = $signed($unsigned((($signed((7'h57)) >> (reg1729 >>> reg1740)) << (~&reg1718))));
          reg1746 <= ({wire1696[(1'h0):(1'h0)],
                  {wire1723[(4'h8):(3'h5)],
                      (7'h4b),
                      ({reg1741} <= $unsigned(wire1697))}} ?
              (!reg1743) : ($signed((7'h54)) | ((7'h4d) | {{reg1711},
                  reg1732[(2'h3):(1'h1)],
                  $signed(reg1737)})));
          reg1747 <= (~&(-(((reg1742 ? reg1732 : (8'hb8)) ?
              reg1731[(1'h0):(1'h0)] : (-reg1700)) > reg1737[(3'h7):(3'h4)])));
          if ((reg1711[(4'he):(4'he)] ?
              ($unsigned((^(wire1723 + reg1730))) ?
                  (&reg1728) : wire1699) : (~($unsigned($unsigned((8'ha1))) ?
                  wire1722[(2'h2):(2'h2)] : ($unsigned(reg1746) ?
                      reg1740 : (reg1737 ? reg1734 : reg1702))))))
            begin
              reg1748 <= $signed(reg1738);
              reg1749 <= (reg1737 * $unsigned((+{(reg1718 <= (8'ha7)),
                  wire1697[(4'hd):(2'h2)],
                  $signed(reg1732)})));
              reg1750 = ((!(($signed(reg1712) == (reg1749 ^ reg1747)) ?
                  $unsigned((reg1740 | wire1722)) : $unsigned((^reg1700)))) || $unsigned(reg1745));
              reg1751 = $unsigned($signed(($unsigned((wire1697 ?
                      reg1702 : (8'ha7))) ?
                  $signed({reg1733}) : {reg1734, $signed(wire1724)})));
              reg1752 <= wire1697[(4'hd):(3'h7)];
              reg1753 = (~$unsigned($unsigned((~^$unsigned(reg1730)))));
            end
          else
            begin
              reg1750 = {reg1711[(4'he):(4'he)], reg1738[(4'h8):(4'h8)]};
              reg1752 <= $unsigned((+(reg1734[(1'h1):(1'h0)] - (&$signed(wire1698)))));
              reg1754 <= $unsigned(reg1734);
              reg1755 <= (~$signed((({reg1712,
                      reg1737} ^~ reg1751[(4'hc):(3'h6)]) ?
                  $signed((^~reg1746)) : reg1753)));
              reg1756 = $signed(($unsigned(((+(8'hbb)) == $unsigned((8'hae)))) - reg1718[(3'h4):(1'h0)]));
              reg1757 = $signed($unsigned(($unsigned($unsigned(forvar1732)) ?
                  {reg1753,
                      $signed(reg1747),
                      (reg1700 ?
                          wire1696 : wire1722)} : $unsigned(((8'h9e) + reg1746)))));
            end
        end
      else
        begin
          for (forvar1744 = (1'h0); (forvar1744 < (1'h0)); forvar1744 = (forvar1744 + (1'h1)))
            begin
              reg1746 <= ($unsigned({$unsigned((|reg1733))}) ?
                  $unsigned(reg1747[(3'h5):(3'h5)]) : $unsigned({(reg1728[(5'h10):(1'h0)] ~^ $unsigned(reg1712))}));
              reg1750 = (wire1696[(2'h3):(1'h1)] ?
                  ((reg1750 ^ (~^(7'h41))) ?
                      (&(reg1737[(1'h0):(1'h0)] ?
                          {(8'hb8)} : reg1732)) : {(reg1702 ?
                              (reg1751 ?
                                  reg1732 : wire1697) : reg1754[(4'h9):(1'h1)]),
                          ((^~reg1729) ?
                              reg1757 : $unsigned(wire1722))}) : $unsigned({reg1731[(1'h1):(1'h1)]}));
              reg1752 <= $signed(($unsigned(reg1735[(4'he):(2'h3)]) <<< reg1743[(5'h10):(2'h2)]));
              reg1754 <= reg1752;
            end
          reg1755 <= reg1744[(2'h2):(1'h1)];
          reg1756 = (|wire1698);
          reg1757 = (~(~(reg1737[(2'h3):(2'h3)] ?
              reg1732 : ((~|(8'hb8)) ? (reg1751 || wire1724) : (&(7'h50))))));
        end
      reg1758 = ((~^reg1728) ? reg1730 : (~&(|reg1735)));
    end
  module1759 #() modinst2636 (.wire1764(reg1707), .wire1761(reg1749), .clk(clk), .wire1760(wire1722), .wire1763(reg1702), .wire1762(wire1723), .y(wire2635));
  always
    @(posedge clk) begin
      reg2637 <= $unsigned(reg1736);
      if (($signed(reg1749[(5'h11):(3'h4)]) ?
          ($signed(((reg1711 ^~ reg1747) ?
                  {wire1722, wire1696, reg1744} : reg1700)) ?
              ((reg1728 ? (~^reg1707) : wire1725) ?
                  {$unsigned((7'h42)),
                      wire1725,
                      $unsigned(reg1735)} : $signed((reg1746 != reg1729))) : $signed(reg1711)) : (((^~(~^wire1722)) ?
                  ((reg1707 ? reg1744 : reg1749) ?
                      (7'h47) : $signed((8'hb2))) : (~|$unsigned(wire1723))) ?
              {$signed($signed(reg1736)),
                  $unsigned(wire1696)} : (-($unsigned(wire1696) && wire1724)))))
        begin
          if (($signed($signed($signed((!wire2635)))) * reg1729[(4'h8):(3'h7)]))
            begin
              reg2638 <= reg2637;
              reg2639 = $signed(reg1707);
              reg2640 <= (~&(wire1696 & {($unsigned(wire1697) >= {reg1754,
                      reg1711}),
                  wire2635,
                  $unsigned((|reg1718))}));
              reg2641 <= (~|$unsigned(wire1724[(2'h3):(2'h3)]));
              reg2642 = (~$signed((($signed(wire1696) ?
                      $signed(wire1696) : $unsigned(reg2638)) ?
                  (wire1722[(4'hf):(4'hb)] ~^ (+reg2639)) : $unsigned((|reg1734)))));
              reg2643 = reg1711;
            end
          else
            begin
              reg2639 = $unsigned($unsigned($unsigned($signed($unsigned(wire1698)))));
              reg2640 <= (reg1728[(3'h4):(1'h0)] ^~ {{(+(wire1722 >= reg1711))},
                  (reg1747 ?
                      (reg1731[(2'h3):(2'h2)] | (reg1744 ?
                          reg1754 : reg1711)) : reg1749)});
            end
        end
      else
        begin
          if (((~^((reg1712 > $signed(wire1699)) ?
                  ((~&reg1712) >= (wire1696 | reg1754)) : (-wire1697))) ?
              (wire1725 <= {wire1722[(4'ha):(3'h7)],
                  $signed($unsigned(reg1702))}) : (wire1699 == $signed((~$unsigned((7'h4e)))))))
            begin
              reg2638 <= (+($signed(reg1718[(4'hb):(1'h0)]) ?
                  wire1724 : $unsigned(wire1724)));
              reg2639 = reg1728[(3'h5):(1'h1)];
            end
          else
            begin
              reg2639 = $signed({$signed($unsigned($unsigned(reg2637)))});
            end
          reg2642 = (^reg1735);
        end
    end
  module2644 #() modinst2689 (wire2688, clk, reg1749, reg1720, reg2640, reg1731);
  always
    @(posedge clk) begin
      for (forvar2690 = (1'h0); (forvar2690 < (2'h2)); forvar2690 = (forvar2690 + (1'h1)))
        begin
          reg2691 = $signed(($unsigned((~|((8'hb8) <= reg1746))) | $signed(wire1723)));
          reg2692 <= ((^reg2640) ?
              (reg1718[(5'h12):(3'h7)] > {reg1736[(2'h3):(2'h3)]}) : {($signed((+wire2688)) ?
                      (&(8'hb5)) : (8'had)),
                  reg1736[(3'h6):(2'h3)]});
          reg2693 <= (-reg1736[(4'ha):(1'h0)]);
          reg2694 <= {(reg1718 << $unsigned((wire2688 & (reg1746 && reg1754))))};
          for (forvar2695 = (1'h0); (forvar2695 < (3'h6)); forvar2695 = (forvar2695 + (1'h1)))
            begin
              reg2696 <= (($signed((-$unsigned((8'hba)))) | (!(!$unsigned((7'h51))))) <= $signed($signed((!$signed(reg1748)))));
              reg2697 = forvar2695;
            end
        end
      if ({(&reg1734[(1'h0):(1'h0)]),
          $unsigned(reg1748),
          {reg1735[(5'h16):(3'h4)]}})
        begin
          reg2698 = $unsigned($signed($signed(reg1735[(5'h11):(4'h8)])));
          reg2699 = ($signed(reg1707[(2'h3):(1'h0)]) ^ reg1718);
          reg2700 = (-$unsigned(reg1712[(1'h0):(1'h0)]));
          reg2701 = $unsigned($signed($unsigned(({wire1723, reg2692, reg2696} ?
              $unsigned(reg1734) : (!reg1728)))));
          reg2702 <= $signed($signed($signed($signed(reg2694))));
          reg2703 <= (~|$unsigned($signed((8'ha4))));
        end
      else
        begin
          if ((((~&reg1728[(1'h1):(1'h1)]) ?
                  (!wire1722) : $signed((^(reg1749 ? wire1725 : (7'h52))))) ?
              (&$signed((^~{reg1735,
                  (7'h57),
                  (7'h4b)}))) : ($unsigned((7'h4d)) | ($unsigned(wire1724[(5'h1d):(5'h11)]) ?
                  $unsigned((reg1748 >>> reg1752)) : (reg1729[(1'h0):(1'h0)] ~^ (reg1728 ?
                      (8'hab) : wire1724))))))
            begin
              reg2702 <= ((+reg2693[(1'h0):(1'h0)]) >= reg1734[(2'h2):(2'h2)]);
              reg2704 = $unsigned(wire1699[(4'h8):(1'h1)]);
              reg2705 <= {$signed((~&{((8'hae) ^~ reg2637),
                      (reg2699 && reg1728)})),
                  (|reg1755),
                  (~|$signed($signed((forvar2690 ? reg1728 : reg1700))))};
              reg2706 = $unsigned((reg1720[(5'h17):(4'h9)] ?
                  $unsigned(($signed(reg2703) - (reg1718 ?
                      reg1734 : (7'h46)))) : $signed($unsigned(reg2705))));
              reg2707 <= $signed(reg1729[(3'h7):(3'h4)]);
              reg2708 <= reg1748[(1'h0):(1'h0)];
            end
          else
            begin
              reg2698 = (8'ha9);
              reg2699 = (($signed(({(7'h46), reg1720} ?
                          $signed((7'h42)) : $unsigned(wire1722))) ?
                      $signed(reg1754) : $signed(reg1754[(4'ha):(4'h8)])) ?
                  $signed(((reg1754[(3'h6):(3'h5)] ?
                      $unsigned(reg2699) : reg1707) & ($signed(wire1725) || $signed(reg2701)))) : reg1744[(2'h3):(2'h3)]);
              reg2702 <= (reg1712 ?
                  wire1696[(3'h5):(1'h0)] : $signed(wire2688[(4'hd):(4'hd)]));
            end
          reg2709 = {$unsigned(({(wire1725 ? reg2637 : reg1707),
                      (forvar2695 ? reg2641 : (8'ha5))} ?
                  {$unsigned(reg2641), (-reg1748), (7'h47)} : ((7'h40) ?
                      {reg2706, reg2702} : reg2692))),
              (~^($signed($signed(reg1702)) ? (^~reg2698) : reg1720))};
          reg2710 = ($unsigned(reg2696[(4'h8):(3'h4)]) ^ (~(~&reg2709[(5'h1c):(5'h1c)])));
          reg2711 <= {$signed((|reg1755)),
              (|reg2691),
              $signed((&$unsigned($unsigned(reg1700))))};
          if ((reg1754[(3'h5):(2'h2)] * (7'h4d)))
            begin
              reg2712 = (7'h52);
              reg2713 <= reg2707;
              reg2714 = ($unsigned($signed(wire1699)) ? wire1698 : (7'h44));
              reg2715 = $unsigned(((~|($unsigned(reg1754) ?
                      reg2707[(4'hb):(4'hb)] : reg1754)) ?
                  $signed(((7'h43) ?
                      $unsigned((8'ha4)) : $signed(reg2691))) : $signed(((~&reg2711) * (reg1720 ?
                      reg2696 : reg2698)))));
              reg2716 = ((({$signed(wire1725), $signed(reg1728)} ?
                  $signed((reg2691 << reg1734)) : reg2638[(1'h0):(1'h0)]) >> $unsigned(wire1724[(4'hc):(4'ha)])) >= (~^((((7'h4e) && reg1747) ?
                      $signed(wire1697) : $unsigned(reg2637)) ?
                  $unsigned(reg1754[(3'h7):(3'h6)]) : (~|(+wire1723)))));
            end
          else
            begin
              reg2713 <= reg1711[(1'h1):(1'h1)];
            end
          for (forvar2717 = (1'h0); (forvar2717 < (3'h6)); forvar2717 = (forvar2717 + (1'h1)))
            begin
              reg2718 = {{$unsigned(wire1725[(2'h3):(1'h0)])}, (7'h43)};
            end
        end
      if ($unsigned(((reg1729 ?
              ((forvar2690 ? wire1697 : reg2693) ?
                  $unsigned(reg1744) : reg2638[(3'h4):(1'h1)]) : {(reg2699 ^ reg1748),
                  (reg2705 ? reg2705 : reg2696)}) ?
          reg2710[(3'h7):(3'h5)] : $unsigned($unsigned((reg1728 < (8'hbd)))))))
        begin
          reg2719 <= $unsigned($signed((!(~^(reg1752 && reg2693)))));
        end
      else
        begin
          reg2720 = reg1728;
          for (forvar2721 = (1'h0); (forvar2721 < (2'h3)); forvar2721 = (forvar2721 + (1'h1)))
            begin
              reg2722 = reg2713[(5'h18):(4'h8)];
              reg2723 = reg2692;
            end
          for (forvar2724 = (1'h0); (forvar2724 < (3'h6)); forvar2724 = (forvar2724 + (1'h1)))
            begin
              reg2725 <= reg2707;
              reg2726 <= {$unsigned((&$unsigned($unsigned(reg2712))))};
            end
          reg2727 = {reg2693[(5'h12):(3'h5)],
              (-{reg2698,
                  ($signed(reg2692) != (8'ha7)),
                  ($unsigned(wire1699) << {reg1746})}),
              reg1748};
        end
    end
  assign wire2728 = reg1729;
  assign wire2729 = $signed(($signed(reg2702) ?
                        reg2708 : (~&$signed($signed(reg1707)))));
  assign wire2730 = ((7'h53) ?
                        (((wire1724 - reg1736[(3'h7):(3'h6)]) ?
                            {(reg1729 ?
                                    reg1707 : (8'h9e))} : (~(reg1702 - (7'h4b)))) < (-{(reg1718 ?
                                reg2713 : reg1720),
                            {reg1700, wire1696, reg1755},
                            (wire1696 ? reg1711 : (8'ha7))})) : reg2708);
  always
    @(posedge clk) begin
      if ($unsigned((~^(reg2640[(1'h0):(1'h0)] ?
          {(reg1749 ~^ reg2637)} : $unsigned(reg2694)))))
        begin
          reg2731 <= wire1725[(2'h3):(1'h1)];
        end
      else
        begin
          reg2732 = (reg1735 - (($unsigned(reg2640) ?
                  (^~$unsigned(wire1723)) : ($unsigned(wire1722) >>> reg1731)) ?
              {$signed(wire2635[(4'hc):(4'hb)]),
                  reg1731,
                  reg2703} : (&((8'ha9) && (8'hb3)))));
          for (forvar2733 = (1'h0); (forvar2733 < (1'h0)); forvar2733 = (forvar2733 + (1'h1)))
            begin
              reg2734 <= {(7'h53),
                  (reg2702[(4'hf):(4'hc)] ?
                      ($unsigned(reg1747) && (reg1711 ?
                          wire1724[(2'h2):(1'h0)] : (8'ha8))) : $unsigned(($unsigned(reg1729) > {reg1718,
                          reg1754,
                          (8'ha3)}))),
                  $unsigned($unsigned(($signed(wire1722) && (~wire1724))))};
              reg2735 <= {$signed(({{reg2696,
                          reg1752,
                          reg1746}} | reg1707[(2'h2):(1'h1)]))};
              reg2736 <= (^{reg2702[(5'h11):(4'hc)], wire1698[(3'h6):(3'h4)]});
              reg2737 <= (7'h57);
            end
          for (forvar2738 = (1'h0); (forvar2738 < (1'h1)); forvar2738 = (forvar2738 + (1'h1)))
            begin
              reg2739 = ((($signed($signed(reg1734)) ?
                      ((wire1724 << reg2719) >> (7'h4d)) : $unsigned($unsigned(reg2702))) ?
                  reg2696 : $signed(((7'h4d) == (forvar2733 ?
                      reg1700 : reg1720)))) ~^ wire1722[(4'hc):(4'ha)]);
              reg2740 <= (($signed((~|reg2702)) | {$signed((-reg1735))}) || ((^reg1720) ?
                  wire2729 : (~reg2719)));
              reg2741 <= $unsigned(wire2688);
              reg2742 <= ({(^$signed($unsigned(reg1755)))} <<< (reg2737[(4'h9):(3'h6)] ?
                  reg2741 : reg2719[(4'hb):(3'h6)]));
              reg2743 <= reg2739;
              reg2744 = $signed(wire1723[(3'h4):(1'h1)]);
            end
          reg2745 = (reg2696 == $unsigned($unsigned((8'h9e))));
        end
      reg2746 <= $unsigned(((7'h51) && reg2705[(1'h0):(1'h0)]));
      if (($signed((reg2725 || $unsigned(reg1711))) ?
          $unsigned(($unsigned({(8'hb5), reg1712}) ?
              reg2703[(4'h8):(3'h4)] : (^~$unsigned(reg1729)))) : (-reg1720[(3'h4):(2'h3)])))
        begin
          reg2747 <= $signed(reg2746);
          reg2748 = $signed(wire2729[(2'h2):(1'h0)]);
          reg2749 <= reg1734[(1'h1):(1'h0)];
          if ({$unsigned(((reg1747[(1'h0):(1'h0)] * (wire2688 ?
                      wire1697 : (8'hb2))) ?
                  (+(reg1707 ? reg2693 : reg2693)) : (^(reg1728 ^~ reg1735))))})
            begin
              reg2750 = ((&$signed((~^$signed(reg2735)))) >> $unsigned((|$signed((^~reg2640)))));
              reg2751 <= $signed(($unsigned((!{reg2705,
                  reg2641})) ^ reg2705[(4'he):(4'h8)]));
              reg2752 <= reg1749;
              reg2753 <= $unsigned($signed($signed($unsigned(reg1752[(5'h11):(4'hc)]))));
            end
          else
            begin
              reg2751 <= $unsigned((reg2726[(4'h8):(3'h6)] ?
                  (~$unsigned(reg2713)) : (reg2746[(4'h8):(3'h4)] << $unsigned((reg2732 * reg2744)))));
              reg2754 = $unsigned(reg2743);
            end
        end
      else
        begin
          reg2748 = ($signed(((~|wire1698[(4'hd):(4'h8)]) ?
                  (~$signed(reg2742)) : $signed($unsigned(wire1696)))) ?
              $signed(((^~(reg2713 + wire1723)) && (~^(wire1724 ?
                  wire2730 : wire2728)))) : reg1735[(5'h18):(4'hd)]);
        end
      reg2755 = forvar2733[(1'h0):(1'h0)];
      for (forvar2756 = (1'h0); (forvar2756 < (1'h1)); forvar2756 = (forvar2756 + (1'h1)))
        begin
          reg2757 = ($unsigned((|(reg2752 & {reg2707}))) ?
              (($signed(reg2741) ?
                  $unsigned(((8'hb2) <= reg1720)) : reg2640[(5'h13):(1'h1)]) == $signed($unsigned($unsigned(reg1729)))) : $unsigned(reg2753[(5'h10):(3'h4)]));
          reg2758 <= $unsigned((reg2741 ?
              (wire2729[(1'h1):(1'h0)] ?
                  $signed((reg2736 ?
                      reg1746 : wire2688)) : wire1696) : (reg2702[(5'h12):(3'h5)] ?
                  reg2641[(2'h3):(2'h2)] : ({(8'hbf)} <<< (~&wire2728)))));
          reg2759 <= reg2726;
          for (forvar2760 = (1'h0); (forvar2760 < (2'h3)); forvar2760 = (forvar2760 + (1'h1)))
            begin
              reg2761 = wire1696[(1'h0):(1'h0)];
            end
          if (reg2753)
            begin
              reg2762 <= ((~^(8'h9c)) ?
                  ((forvar2738 <= (wire2728 ?
                      ((8'ha9) ^~ reg2746) : $signed(reg1720))) <= (forvar2760 ^~ ((!(7'h4d)) ?
                      (reg2755 >>> reg2746) : $signed(wire2728)))) : {reg1731[(2'h2):(1'h0)],
                      ((~^(!reg2744)) ?
                          reg2755 : ((reg1720 == wire1696) ?
                              reg1747[(2'h2):(1'h1)] : (~&reg2732)))});
              reg2763 = (&reg2702);
              reg2764 = $unsigned(wire2728);
              reg2765 <= wire1698;
              reg2766 <= (^~$signed({$signed((~^reg1748)),
                  reg1755[(4'h8):(3'h6)]}));
            end
          else
            begin
              reg2763 = reg2739[(4'h8):(2'h3)];
              reg2764 = $signed($unsigned(reg1754));
              reg2765 <= reg2758[(2'h3):(2'h2)];
            end
          for (forvar2767 = (1'h0); (forvar2767 < (2'h2)); forvar2767 = (forvar2767 + (1'h1)))
            begin
              reg2768 <= {reg2758,
                  ($unsigned($unsigned(reg1734[(1'h1):(1'h1)])) ?
                      reg1755[(1'h0):(1'h0)] : $signed(($unsigned(wire1722) ?
                          (8'hb9) : $unsigned(reg2637))))};
              reg2769 = wire1697[(1'h0):(1'h0)];
              reg2770 = $signed(((|((reg2736 <= (8'hb9)) ?
                  reg1752[(4'h8):(1'h1)] : reg2766[(1'h0):(1'h0)])) != $unsigned($signed(reg2702[(3'h6):(2'h3)]))));
              reg2771 = $signed(((wire2635 < ({reg1747,
                      reg2753,
                      reg2705} - $signed(reg2762))) ?
                  {(+reg2741[(2'h2):(1'h1)]),
                      ($unsigned(reg2768) == (reg2747 ?
                          reg2705 : reg1747))} : (reg2713[(5'h18):(4'he)] ?
                      ((reg2745 ? (7'h53) : reg2731) ?
                          (7'h44) : (reg2768 ?
                              (8'ha9) : reg2637)) : (reg1748[(5'h15):(5'h15)] != reg2746[(1'h1):(1'h0)]))));
              reg2772 <= (reg1720[(4'ha):(4'h8)] + reg2749);
            end
        end
    end
  always
    @(posedge clk) begin
      reg2773 <= (~&($unsigned((8'ha2)) ?
          reg1749[(5'h17):(3'h6)] : {$unsigned((reg2740 ? reg1747 : wire1723)),
              $signed($unsigned(reg2753))}));
      for (forvar2774 = (1'h0); (forvar2774 < (1'h0)); forvar2774 = (forvar2774 + (1'h1)))
        begin
          for (forvar2775 = (1'h0); (forvar2775 < (3'h4)); forvar2775 = (forvar2775 + (1'h1)))
            begin
              reg2776 <= wire1723[(5'h15):(4'ha)];
              reg2777 = ((reg2694 ?
                      reg1718[(4'hd):(4'h9)] : ($unsigned((wire1698 ?
                          (8'ha6) : reg2751)) ^~ reg2640)) ?
                  (reg1700 <= (reg2713[(5'h17):(2'h3)] - $unsigned($signed(reg2751)))) : (~reg2693[(2'h3):(1'h0)]));
              reg2778 = ($unsigned($unsigned(reg1736[(3'h5):(1'h1)])) == $unsigned(reg1711[(4'hb):(2'h3)]));
            end
          for (forvar2779 = (1'h0); (forvar2779 < (3'h4)); forvar2779 = (forvar2779 + (1'h1)))
            begin
              reg2780 = {(^$unsigned((reg1749 != reg2747))),
                  ((8'hae) ? reg1736 : $unsigned($signed((+(8'ha8))))),
                  reg2762};
              reg2781 = reg2640;
              reg2782 = $signed($unsigned({wire1697[(4'h8):(2'h2)],
                  reg1744,
                  (|$unsigned(wire1722))}));
              reg2783 = $signed($unsigned({$unsigned(reg1744[(2'h2):(1'h0)]),
                  (reg2743[(3'h7):(3'h5)] << (reg2766 ? reg2782 : wire1699)),
                  reg2766[(1'h0):(1'h0)]}));
              reg2784 <= {($signed((reg2773[(3'h7):(3'h6)] ?
                      (reg2705 <= (7'h4b)) : $signed(reg2749))) >>> reg2778)};
            end
          for (forvar2785 = (1'h0); (forvar2785 < (3'h6)); forvar2785 = (forvar2785 + (1'h1)))
            begin
              reg2786 = ((reg1736 ?
                      (reg2702[(5'h11):(3'h5)] + reg1749) : (~|wire1699[(5'h15):(5'h13)])) ?
                  forvar2779 : reg1729[(3'h4):(2'h3)]);
              reg2787 = ((^~$signed((((7'h44) + (8'hbf)) << reg2713[(3'h4):(3'h4)]))) ?
                  (7'h42) : wire2729);
              reg2788 = {(reg2776[(2'h3):(1'h1)] + (reg2638 ?
                      reg2736 : reg2719[(3'h4):(1'h1)])),
                  reg2637};
              reg2789 <= (&$signed({(wire2730 < reg1718)}));
            end
          for (forvar2790 = (1'h0); (forvar2790 < (3'h4)); forvar2790 = (forvar2790 + (1'h1)))
            begin
              reg2791 <= reg2786[(4'he):(4'hb)];
              reg2792 = (^((reg2702[(4'hc):(3'h5)] < {forvar2774[(5'h1a):(3'h5)],
                  reg1728,
                  (reg2781 ? reg1707 : reg2791)}) < (reg1712 && (-reg1731))));
              reg2793 = {$unsigned({reg2768,
                      reg2707,
                      $signed(wire2635[(5'h15):(5'h10)])})};
              reg2794 = wire2728[(3'h7):(1'h1)];
              reg2795 <= {reg2734[(2'h3):(1'h0)],
                  $unsigned((~^$signed((reg2713 ? reg2694 : reg2758))))};
            end
          reg2796 = ({$signed({(~^reg2776), (reg2758 * (7'h50))}),
                  $unsigned($unsigned(reg2743[(3'h4):(1'h0)]))} ?
              (~&reg2731) : {(({reg2789, reg2793} ?
                          $signed(reg2692) : reg2702[(1'h1):(1'h0)]) ?
                      (!reg1749) : reg2694),
                  (reg1731[(2'h2):(2'h2)] ?
                      $unsigned({reg2762,
                          reg2759}) : (wire1697[(3'h4):(1'h1)] >> (reg2789 ?
                          (7'h49) : reg2794))),
                  (reg2778 >= forvar2785)});
        end
      if ((!reg2743))
        begin
          reg2797 = $signed(reg2719);
          reg2798 = reg2782;
          reg2799 <= ($signed((~|$signed(reg2742))) <<< $unsigned(reg2696[(4'hf):(4'hb)]));
        end
      else
        begin
          reg2797 = (8'hb2);
        end
    end
  always
    @(posedge clk) begin
      reg2800 = ((+$unsigned({$unsigned(reg1731)})) ?
          ((^~reg2707[(4'h8):(3'h6)]) ?
              $unsigned(($signed((7'h40)) ?
                  $signed((8'hb3)) : reg2731)) : $unsigned(reg1720[(2'h3):(1'h1)])) : {({reg2703,
                  (reg2749 ? reg2743 : wire2728)} || wire1696),
              $unsigned((8'hb7))});
      for (forvar2801 = (1'h0); (forvar2801 < (1'h1)); forvar2801 = (forvar2801 + (1'h1)))
        begin
          for (forvar2802 = (1'h0); (forvar2802 < (2'h2)); forvar2802 = (forvar2802 + (1'h1)))
            begin
              reg2803 <= ({reg1747,
                      reg1711[(3'h4):(3'h4)],
                      reg1754[(1'h0):(1'h0)]} ?
                  (!(((reg2799 ?
                      reg2703 : (8'ha1)) ^ wire2728) + wire1724[(4'ha):(4'ha)])) : (-(wire1696[(2'h2):(1'h1)] <<< ((~^reg1735) >> $unsigned(reg2725)))));
              reg2804 <= $unsigned(wire1699[(4'ha):(2'h3)]);
            end
          for (forvar2805 = (1'h0); (forvar2805 < (3'h4)); forvar2805 = (forvar2805 + (1'h1)))
            begin
              reg2806 <= $unsigned((~(8'ha9)));
              reg2807 <= $unsigned($unsigned($unsigned((-$unsigned(wire2688)))));
              reg2808 = $signed(reg1752[(3'h7):(3'h5)]);
            end
        end
      if ((&(~&{((reg2752 - (7'h51)) == (reg2702 ? wire1723 : reg2752)),
          $unsigned($signed(reg2725))})))
        begin
          reg2809 <= wire2729[(5'h16):(2'h2)];
          if (wire1697[(5'h12):(3'h5)])
            begin
              reg2810 <= $unsigned((($unsigned({reg2640, reg2641, wire1699}) ?
                      $unsigned((reg1752 ?
                          reg1702 : (7'h4d))) : ($signed((8'hb2)) & $unsigned(wire2688))) ?
                  (((~|wire1698) ?
                      (~|wire1723) : $signed((8'ha4))) + reg2784) : reg2806));
            end
          else
            begin
              reg2810 <= $signed($unsigned((reg2703 ?
                  $signed(((7'h55) ^ (7'h43))) : ((reg2708 != wire1697) || reg2742[(5'h10):(4'hc)]))));
              reg2811 <= reg1754[(3'h7):(1'h1)];
              reg2812 = (-(reg2719[(4'he):(4'ha)] & $signed(({reg2800} <= (^~reg2735)))));
              reg2813 <= reg2737[(3'h5):(3'h5)];
              reg2814 <= $signed($unsigned(reg1734));
            end
          reg2815 <= reg2693;
        end
      else
        begin
          for (forvar2809 = (1'h0); (forvar2809 < (2'h3)); forvar2809 = (forvar2809 + (1'h1)))
            begin
              reg2812 = ((-reg1707) << (~^(+(~^$signed(reg2800)))));
            end
          for (forvar2813 = (1'h0); (forvar2813 < (3'h6)); forvar2813 = (forvar2813 + (1'h1)))
            begin
              reg2814 <= reg2641;
              reg2815 <= $unsigned($unsigned((^$signed($signed(reg1718)))));
              reg2816 = reg1734[(2'h3):(1'h0)];
              reg2817 <= (+$unsigned(($signed((reg2753 || reg2765)) ?
                  wire2635[(5'h13):(4'hb)] : (^reg2772[(5'h13):(1'h1)]))));
              reg2818 = reg2813[(5'h1b):(5'h19)];
              reg2819 = (^((((forvar2802 * reg2816) >= reg2696) ?
                      reg1747[(3'h5):(2'h3)] : (7'h42)) ?
                  $signed(((reg1702 ? reg1702 : forvar2801) == (reg2817 ?
                      wire1696 : (7'h49)))) : reg2640));
            end
        end
    end
  assign wire2820 = (^~$unsigned({$signed((wire1723 ? reg1735 : reg2705)),
                        $signed($unsigned(wire2635)),
                        $signed((reg2703 > wire2729))}));
  assign wire2821 = ({$unsigned($signed((reg1754 << reg2768))), (7'h4d)} ?
                        reg2749 : $unsigned((^(-reg2731[(3'h5):(3'h5)]))));
  assign wire2822 = (7'h43);
  assign wire2823 = $unsigned(($signed($unsigned((!(7'h55)))) & (-(+(reg1734 ?
                        reg2741 : wire1698)))));
  always
    @(posedge clk) begin
      reg2824 <= ($unsigned($signed((&(~reg2762)))) > ((~|((~^reg2784) ?
              $signed(reg2776) : reg2719)) ?
          wire2823[(2'h3):(1'h0)] : (($unsigned(reg1720) ^ (reg2696 * wire2729)) || $signed(reg2741))));
      reg2825 = (^$signed((~^(reg2814[(1'h1):(1'h1)] & reg2711))));
      if ((({$signed(reg2809)} ?
              $signed(($signed(wire1698) <= (reg2640 ?
                  wire1696 : (8'hb0)))) : (~^$signed($signed(reg2762)))) ?
          {$unsigned((~|(wire2635 != reg2734)))} : (~^reg2806)))
        begin
          for (forvar2826 = (1'h0); (forvar2826 < (2'h2)); forvar2826 = (forvar2826 + (1'h1)))
            begin
              reg2827 <= reg1700[(3'h7):(2'h3)];
              reg2828 <= reg2804;
              reg2829 = $signed(reg1748);
              reg2830 = (~&$unsigned(((reg1729[(1'h1):(1'h1)] ?
                  reg2693 : $signed(reg1711)) == (^(8'haa)))));
              reg2831 <= $signed($signed($signed(($signed(wire2728) ?
                  $signed(reg2707) : (reg1747 >> reg2753)))));
              reg2832 = reg1711;
            end
          if (reg1735[(5'h12):(5'h11)])
            begin
              reg2833 = (reg2640 ?
                  $signed(wire2688[(5'h17):(4'hb)]) : {$signed(($unsigned(wire2635) >>> reg1736))});
              reg2834 = wire2728[(4'h8):(3'h4)];
              reg2835 <= reg2832;
              reg2836 <= ((reg2765 || ($unsigned((reg2707 ?
                  reg2638 : reg2829)) + $unsigned({reg2741,
                  wire1722}))) >>> (-$unsigned($signed({(8'hbb), wire1697}))));
            end
          else
            begin
              reg2835 <= ((!((8'haa) << (-wire1725[(1'h0):(1'h0)]))) ~^ $unsigned((~$unsigned((wire2730 ?
                  reg1748 : reg2813)))));
              reg2836 <= $signed($signed(reg1712[(2'h2):(1'h1)]));
              reg2837 = $unsigned(reg2741);
              reg2838 = $unsigned($unsigned((~^(+reg2811))));
            end
          reg2839 = wire1696;
          reg2840 = wire2822[(2'h2):(1'h1)];
          reg2841 <= (&reg2832);
          reg2842 = reg2726;
        end
      else
        begin
          for (forvar2826 = (1'h0); (forvar2826 < (1'h0)); forvar2826 = (forvar2826 + (1'h1)))
            begin
              reg2827 <= {{$signed(($signed(reg2804) ?
                          (reg1700 && wire1698) : $unsigned(reg2825))),
                      (~^$signed((&reg2809))),
                      ($signed($signed(reg2740)) ?
                          reg2795[(4'h8):(3'h5)] : wire2728)},
                  (8'ha7),
                  $unsigned((wire2821 ?
                      $unsigned(reg2707) : ((reg2759 << reg2751) >= reg2830)))};
              reg2828 <= $unsigned(($signed(reg2803[(3'h7):(3'h5)]) ?
                  (reg2736 + {(^reg2707)}) : (~|$signed((reg2827 >> (8'ha7))))));
              reg2831 <= reg2791[(2'h2):(2'h2)];
              reg2832 = $unsigned((reg2813[(3'h7):(3'h4)] && $unsigned($unsigned((reg2799 <= reg2835)))));
              reg2833 = (7'h4c);
              reg2835 <= (^~reg1746[(2'h3):(1'h0)]);
              reg2836 <= reg1711;
            end
          reg2837 = {$unsigned(reg2640), $signed(reg2830)};
          for (forvar2838 = (1'h0); (forvar2838 < (1'h1)); forvar2838 = (forvar2838 + (1'h1)))
            begin
              reg2839 = ($unsigned(((-(reg2705 != (8'hb2))) & ($signed(wire2822) ?
                  (wire2688 ?
                      reg2841 : reg2713) : $unsigned(reg2753)))) ^ reg2837[(4'hd):(4'hb)]);
              reg2841 <= (~^$signed(({{reg2836, (7'h56), reg2836},
                      (reg2824 == reg2830)} ?
                  (~(reg2824 ?
                      wire1699 : reg2736)) : $signed(reg2746[(4'hb):(4'h8)]))));
              reg2842 = $unsigned(reg2803);
              reg2843 <= (-({(|(reg2791 ? reg2835 : reg1731)),
                  (~^{reg1749})} <= reg1744[(1'h0):(1'h0)]));
              reg2844 = {{(~&reg2825)}};
              reg2845 <= reg2815[(1'h1):(1'h1)];
              reg2846 = $unsigned($signed((reg2694 << $unsigned({reg1707,
                  reg2825,
                  reg2840}))));
            end
        end
      if (($unsigned((($signed(reg2791) ?
              (&reg2827) : (reg1744 >> (8'hac))) <= reg2641)) ?
          $signed(wire1698) : (($unsigned($signed(reg2734)) >> $signed({reg1700})) && (&$signed(reg2758)))))
        begin
          reg2847 = (((~$signed($signed(reg2726))) ?
                  {($signed(reg2749) ?
                          $unsigned(reg2829) : $signed(reg1731))} : $unsigned(((reg2810 ?
                      reg2828 : reg2772) || (-reg2803)))) ?
              $unsigned((!$unsigned((wire1697 >> wire2728)))) : reg2765[(4'h9):(2'h2)]);
        end
      else
        begin
          for (forvar2847 = (1'h0); (forvar2847 < (3'h6)); forvar2847 = (forvar2847 + (1'h1)))
            begin
              reg2848 = reg2847;
              reg2849 = ($signed((~((reg2702 ^ (8'had)) ?
                  {wire2728} : reg2824))) >= $unsigned($signed($signed(reg2834[(3'h4):(1'h1)]))));
            end
          if ($signed($signed($signed(($signed(reg2713) <= (&reg2752))))))
            begin
              reg2850 <= $unsigned((~^(|reg1736[(2'h2):(1'h0)])));
              reg2851 <= (((reg2776 || reg2640[(5'h12):(3'h4)]) - $signed(((~&reg2753) ?
                      (reg2832 ? reg2766 : wire1697) : (reg2813 ?
                          (8'ha3) : reg1707)))) ?
                  $unsigned(wire1698[(3'h6):(3'h4)]) : $unsigned($signed(reg1744[(1'h1):(1'h0)])));
            end
          else
            begin
              reg2850 <= (~$signed($signed($unsigned(reg2830[(4'h8):(3'h7)]))));
              reg2852 = $unsigned($unsigned((^((reg1749 ?
                  reg2827 : wire2823) <<< $signed(reg2827)))));
              reg2853 <= $signed((^~(reg2713[(4'hc):(2'h3)] ?
                  $signed((-reg2707)) : reg2746[(4'h8):(1'h1)])));
              reg2854 <= $signed(reg1752[(3'h5):(3'h5)]);
              reg2855 = (reg1712[(1'h1):(1'h1)] != reg1718);
              reg2856 <= {$signed($unsigned(((reg2703 <<< reg1700) * reg1734))),
                  $signed((((wire2728 ? forvar2826 : reg1702) ?
                          $unsigned((7'h49)) : (!reg2837)) ?
                      (~&$signed(reg2746)) : ((8'hb7) ?
                          (reg1728 ? reg2828 : reg2840) : (~&(8'hb7))))),
                  {(reg2703[(4'hb):(1'h1)] ? reg2766 : $signed(reg2843))}};
            end
          reg2857 = (~|reg2731[(4'ha):(4'h9)]);
          for (forvar2858 = (1'h0); (forvar2858 < (2'h3)); forvar2858 = (forvar2858 + (1'h1)))
            begin
              reg2859 <= $unsigned((reg2828 >= reg1735[(4'hb):(3'h4)]));
              reg2860 <= (+$signed($signed(wire2688[(4'hf):(4'h8)])));
            end
          reg2861 <= (~&reg2839[(2'h3):(1'h0)]);
          reg2862 = {((reg2735[(2'h3):(2'h2)] ?
                      $unsigned({wire1722,
                          wire1698,
                          reg2703}) : reg2803[(5'h15):(1'h0)]) ?
                  reg2740[(5'h10):(4'hd)] : reg2765[(3'h6):(1'h0)]),
              ({reg1736[(1'h0):(1'h0)]} != $signed((^~((8'hae) ?
                  reg2737 : (8'ha0))))),
              (~$signed(reg2734))};
        end
    end
  assign wire2863 = (^{reg1734[(1'h0):(1'h0)],
                        (wire1722[(5'h13):(5'h11)] != $unsigned($signed(reg2856)))});
  assign wire2864 = $unsigned((((~|(reg1718 ? wire1722 : (8'had))) ?
                            ($unsigned(reg2843) & $unsigned(reg1700)) : ($unsigned(wire1725) ?
                                (reg2703 + reg2726) : reg2640)) ?
                        reg2734[(5'h11):(5'h10)] : reg2799[(4'he):(4'ha)]));
  always
    @(posedge clk) begin
      for (forvar2865 = (1'h0); (forvar2865 < (3'h5)); forvar2865 = (forvar2865 + (1'h1)))
        begin
          reg2866 <= reg2841[(5'h13):(2'h3)];
          if (((&{$signed(reg2753[(4'hd):(4'hc)])}) + {($signed(reg2742[(4'he):(4'hb)]) ?
                  reg1749[(1'h0):(1'h0)] : ({reg1731} ?
                      (reg2749 ?
                          reg2734 : reg1754) : reg2851[(4'hf):(4'hf)]))}))
            begin
              reg2867 = $signed((($signed((reg2693 ?
                      wire2823 : reg2804)) + $unsigned((reg2827 ?
                      wire1697 : reg2762))) ?
                  $unsigned(reg2850) : {($unsigned(reg1711) | ((8'hb3) ~^ reg2831)),
                      (&(reg2751 == reg2850))}));
              reg2868 = {$signed($unsigned({(reg2859 ? (8'hbe) : reg2813),
                      $signed(reg1746)}))};
              reg2869 = reg1752[(5'h14):(2'h2)];
              reg2870 = (-(~&reg2831));
            end
          else
            begin
              reg2871 <= $signed(reg2811[(3'h7):(2'h2)]);
              reg2872 <= {$signed(((wire2820 ?
                          (wire2822 ? (8'had) : wire2635) : (!reg1747)) ?
                      $unsigned(wire2730) : reg1746[(1'h0):(1'h0)])),
                  (reg2694 ?
                      $signed($unsigned(reg1702[(3'h7):(2'h2)])) : $signed(reg2866))};
              reg2873 <= reg2707;
            end
          reg2874 = reg2836;
        end
      reg2875 <= ((^(($signed(reg1718) ? (8'ha0) : (~&reg2870)) ?
          $signed(reg2795) : $signed({wire1725}))) > (reg2713 ?
          (~|(|reg2870)) : ((wire2863[(2'h2):(1'h0)] ?
                  {wire1698, reg2751, reg2758} : forvar2865) ?
              wire2729[(5'h16):(5'h11)] : reg2742[(4'h9):(3'h6)])));
    end
  assign wire2876 = $unsigned(wire2823[(2'h2):(1'h1)]);
  module2877 #() modinst2888 (.wire2878(reg2814), .wire2881(reg2746), .wire2882(reg1720), .wire2879(reg2776), .clk(clk), .wire2880(reg2845), .y(wire2887));
  assign wire2889 = reg2807[(4'hf):(4'hf)];
  assign wire2890 = {(($unsigned($signed(wire1724)) >> wire2887) ?
                            reg2813 : $unsigned($signed(wire2820[(3'h7):(2'h2)]))),
                        reg2766};
  assign wire2891 = ((!(reg2765 & ($unsigned((7'h41)) ?
                        $signed(wire1725) : $unsigned(reg2694)))) < (((+(reg2843 ?
                        reg1700 : wire2876)) <= $signed(wire2730)) > $signed($unsigned({wire2890}))));
  assign wire2892 = (7'h4a);
  always
    @(posedge clk) begin
      reg2893 = ($unsigned((~&{(^reg2731)})) > reg1711);
      reg2894 = (reg2850[(4'hd):(3'h7)] ?
          reg2861 : ($unsigned(reg2817[(5'h12):(4'h8)]) ~^ $signed(reg2696[(3'h7):(1'h0)])));
      for (forvar2895 = (1'h0); (forvar2895 < (3'h5)); forvar2895 = (forvar2895 + (1'h1)))
        begin
          reg2896 = reg1736;
          for (forvar2897 = (1'h0); (forvar2897 < (2'h3)); forvar2897 = (forvar2897 + (1'h1)))
            begin
              reg2898 = reg1754[(3'h5):(2'h3)];
              reg2899 = (~&(|reg2853));
              reg2900 <= $signed(wire2864);
              reg2901 = $unsigned($signed((7'h43)));
              reg2902 <= reg2873[(4'hf):(2'h2)];
              reg2903 = ($unsigned($unsigned({reg2799[(5'h1b):(4'ha)],
                      $signed(reg2693)})) ?
                  {$unsigned({{(8'hbd), (8'hb8), wire1722},
                          $signed(wire2730)})} : (((((8'hba) == reg2811) >> (reg2696 ?
                          wire1725 : reg2734)) <<< reg2811) ?
                      (&reg1718) : ($unsigned(((8'ha6) ? reg2806 : reg2789)) ?
                          reg2747 : $unsigned({reg2735}))));
              reg2904 <= (^~((reg2742[(3'h5):(3'h4)] ?
                  reg2806 : $unsigned((wire1724 ?
                      reg2703 : reg2853))) ^~ $unsigned(reg1744)));
            end
          for (forvar2905 = (1'h0); (forvar2905 < (2'h2)); forvar2905 = (forvar2905 + (1'h1)))
            begin
              reg2906 = $signed($unsigned(reg2866[(3'h6):(1'h1)]));
              reg2907 <= reg1711;
              reg2908 <= $signed($signed(reg2873[(2'h2):(1'h1)]));
              reg2909 = $unsigned(($signed((7'h4d)) != reg2708));
            end
          if ($signed(reg2743[(4'ha):(3'h4)]))
            begin
              reg2910 = reg2731;
              reg2911 = (~(&reg2900[(5'h10):(4'ha)]));
              reg2912 = $unsigned($unsigned(($unsigned($unsigned(reg2810)) + reg2772[(5'h13):(4'h9)])));
              reg2913 = ($unsigned(($unsigned((~|reg2807)) ?
                  (reg1747 << {reg2894}) : (8'hb5))) != forvar2905);
            end
          else
            begin
              reg2914 <= {(reg2638 ?
                      wire1699[(4'ha):(3'h6)] : ($unsigned(wire2891[(2'h3):(1'h0)]) ?
                          (~|((7'h41) ?
                              reg2711 : reg2859)) : wire1724[(5'h1c):(3'h6)])),
                  forvar2905[(5'h16):(4'hc)]};
              reg2915 = {reg2860[(3'h6):(3'h4)],
                  ($signed($unsigned((-reg1702))) & (|($unsigned(reg2789) | (reg1707 * reg2866))))};
            end
          if ($signed(((~^$unsigned((-(7'h53)))) != $unsigned((+$signed(wire2864))))))
            begin
              reg2916 = ($unsigned(reg2753[(4'hd):(3'h6)]) ?
                  $signed($signed($signed(((8'ha2) ?
                      reg2707 : reg2707)))) : (($signed($unsigned(wire2635)) ?
                      $unsigned((~(8'hb1))) : $signed($signed(reg2768))) && (&(7'h54))));
              reg2917 = {(reg2807 * $unsigned(wire2823[(1'h0):(1'h0)]))};
            end
          else
            begin
              reg2918 <= (~&(~|$signed((reg2872[(3'h5):(3'h5)] <<< {reg2856}))));
              reg2919 = (+(+(!({reg2762, wire1724} ?
                  reg2694[(1'h0):(1'h0)] : (reg2694 <<< reg1728)))));
              reg2920 <= reg2856;
              reg2921 = reg2919;
              reg2922 <= ($signed($signed((~&$signed(reg2762)))) > (7'h44));
              reg2923 <= ((($signed(reg2922) ?
                      wire1696[(1'h0):(1'h0)] : (-$unsigned(reg2919))) + reg1728) ?
                  (reg2766 ?
                      (~&(wire2688 ?
                          {wire2823} : {reg2705,
                              reg2910})) : ($signed(reg2899) >>> reg2803)) : reg2784);
            end
          for (forvar2924 = (1'h0); (forvar2924 < (2'h2)); forvar2924 = (forvar2924 + (1'h1)))
            begin
              reg2925 <= reg2828[(3'h6):(2'h3)];
              reg2926 = wire2863;
              reg2927 = {$signed((((wire1699 <<< reg2746) ?
                          (~&(7'h55)) : forvar2924) ?
                      reg2705 : ((reg2926 ? reg2784 : wire2728) ?
                          (wire1723 ? reg2705 : reg2913) : {reg2711})))};
              reg2928 = {wire2822[(2'h3):(1'h1)],
                  (($unsigned((reg2708 == reg2809)) ?
                      $unsigned(((8'hb6) - wire1698)) : (-(reg2836 + reg2742))) <<< wire2688[(5'h10):(4'ha)]),
                  {(reg1747 ?
                          ((reg2696 ? reg2854 : reg2740) ?
                              reg2799 : $unsigned(reg2740)) : reg2696),
                      reg2807}};
              reg2929 = (!$signed(((reg2725 ^ reg2637[(1'h1):(1'h1)]) ?
                  ($signed(reg2854) ?
                      {(7'h50),
                          (8'had)} : wire1725[(2'h2):(1'h0)]) : (reg2795[(3'h7):(2'h3)] | $unsigned(reg2893)))));
            end
        end
      if ((wire1696 ?
          (((8'hb4) ? reg2696 : reg1749[(4'hd):(1'h0)]) ?
              ((reg1702[(5'h16):(5'h13)] ?
                      $unsigned(reg2731) : (reg2917 ? reg2841 : wire1696)) ?
                  $unsigned((^reg2641)) : {(reg2746 ? (7'h46) : wire1724),
                      ((8'hb1) - (7'h49))}) : reg2806) : $signed(reg2641)))
        begin
          for (forvar2930 = (1'h0); (forvar2930 < (2'h3)); forvar2930 = (forvar2930 + (1'h1)))
            begin
              reg2931 = reg2911;
              reg2932 <= (reg2831 ?
                  $unsigned($signed($signed((8'hb3)))) : (((!((7'h58) ?
                          (8'hb9) : reg2916)) ?
                      $unsigned(reg2900) : (((8'ha6) ? reg1720 : reg2836) ?
                          {(8'hbb)} : ((8'hb2) ?
                              reg2918 : reg2914))) * ((&reg2836) >>> $signed(reg2894[(4'ha):(3'h7)]))));
            end
          reg2933 <= reg2911[(1'h0):(1'h0)];
          reg2934 = $signed((~|{(&reg1755), $unsigned((reg2736 <= reg2817))}));
          if ($unsigned((~((reg2856 ?
              (reg1749 ? reg2866 : reg2747) : reg1712) || ((reg2932 ?
              reg2856 : reg2784) && (reg1747 < reg2725))))))
            begin
              reg2935 <= reg2693[(3'h7):(2'h3)];
            end
          else
            begin
              reg2935 <= $unsigned((8'h9e));
              reg2936 <= wire2729;
            end
        end
      else
        begin
          if (({{((-wire2889) * (reg2933 ^~ (7'h4c)))},
                  reg2898[(5'h11):(3'h4)]} ?
              (|(reg2725[(5'h10):(3'h6)] ?
                  (^((8'h9e) <= wire2822)) : (~^(~reg2799)))) : (^reg1711[(4'hb):(3'h5)])))
            begin
              reg2930 = $unsigned(((reg2933 ?
                      (((8'haf) << reg2907) ?
                          $signed(reg2920) : reg2734) : $unsigned($unsigned(reg2817))) ?
                  ({(reg2831 + reg2725), (&reg2726)} ?
                      wire2887 : reg2811[(3'h5):(1'h0)]) : $signed(((+reg2759) + (|reg1736)))));
            end
          else
            begin
              reg2930 = (reg2904 ~^ (~|reg1718));
              reg2931 = ((^~reg1735) ?
                  reg2893 : (~$signed(reg2926[(5'h18):(4'ha)])));
              reg2932 <= (wire2729 ? reg2922[(3'h4):(2'h2)] : $signed((8'ha7)));
              reg2933 <= ((reg2904[(3'h6):(1'h1)] < reg1700) ?
                  (^~($signed($signed(wire2823)) ?
                      {$unsigned(reg2931)} : (reg1752 <<< reg2638))) : ((^~reg1752) + (7'h53)));
              reg2934 = $signed((reg2713[(5'h18):(4'hf)] ?
                  (-((!reg2827) ?
                      (reg2910 <= reg2854) : $signed(reg2759))) : {(((8'hbd) ?
                              reg2827 : reg2831) ?
                          (~wire1696) : (reg2933 + wire2891))}));
            end
        end
      for (forvar2937 = (1'h0); (forvar2937 < (1'h1)); forvar2937 = (forvar2937 + (1'h1)))
        begin
          for (forvar2938 = (1'h0); (forvar2938 < (3'h6)); forvar2938 = (forvar2938 + (1'h1)))
            begin
              reg2939 = reg2827;
              reg2940 = forvar2905;
              reg2941 <= reg1744[(1'h0):(1'h0)];
              reg2942 = ({(!$signed((reg2835 ?
                      reg2923 : (8'hae))))} < wire2864);
              reg2943 = (((reg1735 ~^ reg2789) ?
                  reg1736 : (8'ha1)) <<< $signed($unsigned((~&(wire2892 ?
                  reg2789 : wire2891)))));
            end
        end
      reg2944 = (~{reg2804[(5'h14):(3'h7)],
          {$signed($unsigned(reg2904)),
              $unsigned(((8'hbc) ? (8'hae) : reg2827))}});
      reg2945 <= reg2931;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2877  (y, clk, wire2882, wire2881, wire2880, wire2879, wire2878);
  output wire [(32'h56):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire2882;
  input wire signed [(5'h1d):(1'h0)] wire2881;
  input wire [(5'h15):(1'h0)] wire2880;
  input wire [(5'h1a):(1'h0)] wire2879;
  input wire signed [(5'h14):(1'h0)] wire2878;
  wire [(5'h18):(1'h0)] wire2886;
  wire [(5'h15):(1'h0)] wire2885;
  wire signed [(5'h10):(1'h0)] wire2884;
  wire signed [(5'h18):(1'h0)] wire2883;
  assign y = {wire2886, wire2885, wire2884, wire2883, (1'h0)};
  assign wire2883 = $signed(wire2879);
  assign wire2884 = $signed((-$signed(wire2879[(1'h1):(1'h0)])));
  assign wire2885 = ((($signed(((8'had) ? wire2880 : wire2881)) ?
                            wire2883 : wire2883[(1'h1):(1'h1)]) ?
                        (8'h9e) : wire2882[(3'h7):(2'h2)]) ~^ (($unsigned((^wire2881)) >= $signed($signed(wire2882))) == (((!wire2880) + $signed((8'hb1))) & (((8'hae) ?
                            wire2882 : wire2880) ?
                        $signed(wire2882) : {(8'hb5)}))));
  assign wire2886 = wire2883;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2644  (y, clk, wire2648, wire2647, wire2646, wire2645);
  output wire [(32'h271):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h18):(1'h0)] wire2648;
  input wire signed [(3'h4):(1'h0)] wire2647;
  input wire signed [(5'h18):(1'h0)] wire2646;
  input wire [(3'h7):(1'h0)] wire2645;
  wire signed [(3'h4):(1'h0)] wire2687;
  wire signed [(4'h8):(1'h0)] wire2670;
  wire signed [(5'h1b):(1'h0)] wire2649;
  reg [(2'h2):(1'h0)] reg2685 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2676 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2680 = (1'h0);
  reg [(5'h19):(1'h0)] reg2678 = (1'h0);
  reg [(4'hf):(1'h0)] reg2674 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2673 = (1'h0);
  reg [(2'h3):(1'h0)] reg2671 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2668 = (1'h0);
  reg [(4'he):(1'h0)] reg2666 = (1'h0);
  reg [(5'h14):(1'h0)] reg2664 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2659 = (1'h0);
  reg [(2'h3):(1'h0)] reg2658 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2656 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2655 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2654 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2652 = (1'h0);
  reg [(3'h7):(1'h0)] reg2650 = (1'h0);
  reg [(3'h5):(1'h0)] reg2686 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2681 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2674 = (1'h0);
  reg [(4'hf):(1'h0)] reg2684 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2683 = (1'h0);
  reg [(5'h10):(1'h0)] reg2682 = (1'h0);
  reg [(4'h9):(1'h0)] reg2681 = (1'h0);
  reg [(3'h6):(1'h0)] reg2679 = (1'h0);
  reg [(4'hc):(1'h0)] reg2677 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2676 = (1'h0);
  reg [(2'h2):(1'h0)] reg2675 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2672 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2669 = (1'h0);
  reg [(5'h18):(1'h0)] reg2667 = (1'h0);
  reg [(4'hd):(1'h0)] reg2665 = (1'h0);
  reg [(5'h16):(1'h0)] reg2663 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2662 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2661 = (1'h0);
  reg [(5'h10):(1'h0)] reg2660 = (1'h0);
  reg [(4'ha):(1'h0)] reg2657 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2653 = (1'h0);
  reg [(5'h17):(1'h0)] reg2651 = (1'h0);
  assign y = {wire2687,
                 wire2670,
                 wire2649,
                 reg2685,
                 reg2676,
                 reg2680,
                 reg2678,
                 reg2674,
                 reg2673,
                 reg2671,
                 reg2668,
                 reg2666,
                 reg2664,
                 reg2659,
                 reg2658,
                 reg2656,
                 reg2655,
                 reg2654,
                 reg2652,
                 reg2650,
                 reg2686,
                 forvar2681,
                 forvar2674,
                 reg2684,
                 reg2683,
                 reg2682,
                 reg2681,
                 reg2679,
                 reg2677,
                 forvar2676,
                 reg2675,
                 reg2672,
                 reg2669,
                 reg2667,
                 reg2665,
                 reg2663,
                 reg2662,
                 forvar2661,
                 reg2660,
                 reg2657,
                 forvar2653,
                 reg2651,
                 (1'h0)};
  assign wire2649 = (wire2647 >= ($unsigned(({wire2645,
                        wire2645,
                        wire2647} >> ((7'h56) | wire2648))) <= {wire2646}));
  always
    @(posedge clk) begin
      reg2650 <= ($unsigned((-($signed((8'ha2)) ?
          wire2649[(5'h14):(4'hd)] : $unsigned(wire2648)))) ^~ wire2646[(5'h17):(5'h17)]);
      reg2651 = ($signed($unsigned((wire2646 ?
              wire2647[(2'h3):(1'h0)] : (wire2645 ? wire2646 : wire2647)))) ?
          ({(!(wire2647 | wire2647))} ?
              (7'h40) : wire2648[(1'h1):(1'h0)]) : $signed($unsigned((~^$unsigned(reg2650)))));
      reg2652 <= ($unsigned(wire2649) > reg2650[(3'h5):(2'h2)]);
      for (forvar2653 = (1'h0); (forvar2653 < (3'h5)); forvar2653 = (forvar2653 + (1'h1)))
        begin
          if (($signed($unsigned($unsigned({reg2650, reg2650}))) | (~|reg2650)))
            begin
              reg2654 <= (|reg2651);
              reg2655 <= $signed($unsigned(reg2650));
              reg2656 <= {{(-((forvar2653 <<< reg2650) ?
                          $signed((8'hb7)) : $unsigned(wire2647))),
                      $signed((wire2649 != forvar2653[(2'h2):(1'h0)]))},
                  $unsigned({{reg2654, (wire2647 ? (7'h4b) : reg2655)},
                      {wire2645}})};
            end
          else
            begin
              reg2654 <= wire2646;
            end
          if ((+wire2646))
            begin
              reg2657 = reg2655;
              reg2658 <= $unsigned((!$signed(($signed((7'h53)) ?
                  wire2649 : reg2655))));
              reg2659 <= $signed(reg2652[(5'h11):(3'h5)]);
            end
          else
            begin
              reg2657 = $signed($signed(($unsigned((^~reg2651)) | reg2656)));
              reg2658 <= $signed($signed(wire2645));
              reg2660 = (^$signed($unsigned(((reg2654 != forvar2653) < wire2647[(3'h4):(2'h2)]))));
            end
          for (forvar2661 = (1'h0); (forvar2661 < (2'h3)); forvar2661 = (forvar2661 + (1'h1)))
            begin
              reg2662 = $unsigned($unsigned((($unsigned((8'h9e)) ?
                      wire2647 : {reg2654}) ?
                  (~wire2646) : (^~reg2651[(1'h0):(1'h0)]))));
              reg2663 = (~^reg2655[(5'h12):(3'h7)]);
              reg2664 <= ($signed(((((8'hbd) - wire2646) >> (&reg2655)) | ({reg2659} ?
                  (reg2650 ?
                      reg2660 : reg2662) : (forvar2653 < reg2663)))) > $signed($unsigned((-reg2652[(4'h9):(2'h2)]))));
              reg2665 = {(forvar2653 ?
                      (~&wire2649) : (^(forvar2661[(2'h2):(2'h2)] || $signed(wire2647)))),
                  (^reg2664[(3'h7):(1'h0)]),
                  $signed((($signed(reg2654) ?
                          $signed(wire2645) : (reg2663 > reg2655)) ?
                      (forvar2653 ?
                          ((7'h50) | wire2646) : $signed(reg2657)) : $unsigned((reg2658 ?
                          reg2659 : forvar2653))))};
              reg2666 <= reg2660;
            end
          reg2667 = (-reg2654);
        end
      reg2668 <= reg2662[(1'h0):(1'h0)];
      reg2669 = ($signed((&{(reg2662 ? reg2662 : (8'hbb)),
          $signed(reg2663)})) ^~ {({$signed(reg2663), reg2650[(1'h1):(1'h0)]} ?
              $signed({reg2655,
                  reg2660,
                  reg2656}) : ($signed(forvar2653) ^ (reg2666 ^ reg2654))),
          ((!(^~forvar2653)) ?
              (!(&(7'h4c))) : ({reg2664, (8'hb3)} * {reg2658,
                  reg2656,
                  reg2655})),
          (reg2655 || {(!reg2650)})});
    end
  assign wire2670 = ({$unsigned(reg2659),
                        reg2656[(4'ha):(2'h2)]} - {$signed(reg2658[(1'h1):(1'h0)]),
                        {reg2658, {(~^reg2654), ((7'h55) - wire2646)}},
                        $unsigned($unsigned($unsigned(wire2646)))});
  always
    @(posedge clk) begin
      reg2671 <= (((((wire2647 ? reg2658 : reg2650) ?
          (reg2656 >> reg2656) : wire2646) && (7'h4b)) - $unsigned($signed((reg2656 | reg2652)))) ^~ $signed(((wire2649[(1'h0):(1'h0)] ?
              (reg2668 ? reg2659 : reg2659) : ((7'h41) >= reg2654)) ?
          wire2670[(4'h8):(1'h0)] : ({reg2652} >= (reg2652 ~^ reg2654)))));
      if (reg2668[(5'h10):(4'hc)])
        begin
          reg2672 = reg2664;
          reg2673 <= $signed(reg2656);
          reg2674 <= $unsigned($unsigned(($unsigned((reg2655 == reg2664)) != (reg2650[(2'h2):(2'h2)] != reg2668[(4'ha):(2'h2)]))));
          reg2675 = $signed((reg2659 & $signed({{reg2650}, (^reg2664)})));
          for (forvar2676 = (1'h0); (forvar2676 < (1'h1)); forvar2676 = (forvar2676 + (1'h1)))
            begin
              reg2677 = $signed($unsigned(($signed((reg2658 * (8'ha1))) ~^ $signed(reg2671[(1'h1):(1'h0)]))));
              reg2678 <= reg2666[(2'h2):(1'h0)];
              reg2679 = reg2674;
              reg2680 <= $signed({(((wire2647 & reg2678) + {wire2647,
                      reg2659,
                      (8'hbc)}) < reg2654),
                  ($unsigned((~&reg2679)) ?
                      ((wire2670 ^~ reg2664) - (~^reg2678)) : $unsigned($signed((8'haf)))),
                  (~(7'h55))});
              reg2681 = {(~($signed((^~reg2654)) ?
                      (8'ha1) : ((reg2650 < reg2677) == (7'h4b)))),
                  (8'haa)};
              reg2682 = (&$unsigned((7'h42)));
            end
          if ($signed(reg2680))
            begin
              reg2683 = $unsigned(reg2671[(2'h3):(1'h0)]);
              reg2684 = (~|(^(8'h9f)));
            end
          else
            begin
              reg2683 = (reg2680 ? reg2658[(2'h2):(1'h0)] : reg2668);
            end
        end
      else
        begin
          reg2673 <= $signed(reg2668[(1'h1):(1'h0)]);
          for (forvar2674 = (1'h0); (forvar2674 < (3'h5)); forvar2674 = (forvar2674 + (1'h1)))
            begin
              reg2676 <= reg2666;
              reg2677 = ({(reg2664[(4'hb):(4'h8)] || (!reg2673[(5'h16):(3'h7)])),
                  reg2676[(4'hf):(1'h1)]} | $signed(wire2646[(5'h14):(5'h11)]));
              reg2679 = ($unsigned(reg2671[(2'h3):(1'h0)]) ?
                  (reg2673 > (reg2666[(1'h1):(1'h1)] <= $unsigned($unsigned(reg2656)))) : ({$unsigned($signed((7'h4c))),
                          ($unsigned(reg2675) <<< reg2683),
                          $signed((wire2646 | forvar2676))} ?
                      $unsigned($signed((-(8'hb7)))) : reg2658[(2'h3):(1'h1)]));
              reg2680 <= reg2658[(2'h3):(1'h1)];
            end
          for (forvar2681 = (1'h0); (forvar2681 < (3'h4)); forvar2681 = (forvar2681 + (1'h1)))
            begin
              reg2682 = (7'h4c);
              reg2685 <= {reg2679};
              reg2686 = $signed({$unsigned((|reg2677)),
                  $signed($unsigned((+(7'h4b))))});
            end
        end
    end
  assign wire2687 = (($unsigned((&((7'h58) + reg2678))) != reg2666[(3'h4):(2'h2)]) && reg2678[(2'h3):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1759  (y, clk, wire1764, wire1763, wire1762, wire1761, wire1760);
  output wire [(32'h37b2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h17):(1'h0)] wire1764;
  input wire signed [(2'h3):(1'h0)] wire1763;
  input wire [(4'hb):(1'h0)] wire1762;
  input wire signed [(5'h1e):(1'h0)] wire1761;
  input wire [(5'h10):(1'h0)] wire1760;
  wire signed [(4'hf):(1'h0)] wire2568;
  wire [(3'h5):(1'h0)] wire2453;
  wire signed [(5'h1b):(1'h0)] wire2208;
  wire [(5'h18):(1'h0)] wire2207;
  wire signed [(3'h4):(1'h0)] wire2043;
  wire [(3'h6):(1'h0)] wire1896;
  wire signed [(3'h5):(1'h0)] wire1765;
  reg [(4'he):(1'h0)] reg2634 = (1'h0);
  reg [(3'h4):(1'h0)] reg2633 = (1'h0);
  reg [(5'h19):(1'h0)] reg2631 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2628 = (1'h0);
  reg [(5'h10):(1'h0)] reg2626 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2625 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2624 = (1'h0);
  reg [(2'h2):(1'h0)] reg2623 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2622 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2620 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2618 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2616 = (1'h0);
  reg [(5'h14):(1'h0)] reg2613 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2612 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2610 = (1'h0);
  reg [(5'h15):(1'h0)] reg2607 = (1'h0);
  reg [(5'h12):(1'h0)] reg2606 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2604 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2603 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2601 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2595 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2592 = (1'h0);
  reg [(3'h6):(1'h0)] reg2591 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2589 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2582 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2578 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2573 = (1'h0);
  reg [(5'h12):(1'h0)] reg2570 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2569 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2567 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2564 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2562 = (1'h0);
  reg [(4'h8):(1'h0)] reg2560 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2558 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2556 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2553 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2552 = (1'h0);
  reg [(4'hd):(1'h0)] reg2551 = (1'h0);
  reg [(3'h7):(1'h0)] reg2548 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2547 = (1'h0);
  reg [(3'h4):(1'h0)] reg2546 = (1'h0);
  reg [(4'hc):(1'h0)] reg2544 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2538 = (1'h0);
  reg [(4'hb):(1'h0)] reg2536 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2535 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2534 = (1'h0);
  reg [(4'h8):(1'h0)] reg2531 = (1'h0);
  reg [(2'h2):(1'h0)] reg2528 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2527 = (1'h0);
  reg [(4'hc):(1'h0)] reg2525 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2523 = (1'h0);
  reg [(4'hb):(1'h0)] reg2518 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2516 = (1'h0);
  reg [(4'hc):(1'h0)] reg2514 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2510 = (1'h0);
  reg [(5'h19):(1'h0)] reg2508 = (1'h0);
  reg [(4'h9):(1'h0)] reg2505 = (1'h0);
  reg [(4'ha):(1'h0)] reg2502 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2501 = (1'h0);
  reg [(4'hb):(1'h0)] reg2500 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2499 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2498 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2496 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2493 = (1'h0);
  reg [(4'h8):(1'h0)] reg2487 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2484 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2482 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2480 = (1'h0);
  reg [(5'h11):(1'h0)] reg2479 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2478 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2477 = (1'h0);
  reg [(2'h2):(1'h0)] reg2476 = (1'h0);
  reg [(4'h8):(1'h0)] reg2471 = (1'h0);
  reg [(3'h4):(1'h0)] reg2470 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2466 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2464 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2461 = (1'h0);
  reg [(2'h2):(1'h0)] reg2454 = (1'h0);
  reg [(5'h10):(1'h0)] reg2450 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2449 = (1'h0);
  reg [(5'h10):(1'h0)] reg2447 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2446 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2444 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2440 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2437 = (1'h0);
  reg [(2'h2):(1'h0)] reg2436 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2433 = (1'h0);
  reg [(3'h7):(1'h0)] reg2422 = (1'h0);
  reg [(5'h15):(1'h0)] reg2420 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2418 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2417 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2414 = (1'h0);
  reg [(4'hb):(1'h0)] reg2413 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2410 = (1'h0);
  reg [(4'hc):(1'h0)] reg2409 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2408 = (1'h0);
  reg [(2'h3):(1'h0)] reg2407 = (1'h0);
  reg [(4'h8):(1'h0)] reg2404 = (1'h0);
  reg [(5'h17):(1'h0)] reg2403 = (1'h0);
  reg [(5'h19):(1'h0)] reg2383 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2401 = (1'h0);
  reg [(4'he):(1'h0)] reg2400 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2396 = (1'h0);
  reg [(5'h17):(1'h0)] reg2395 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2393 = (1'h0);
  reg [(4'hc):(1'h0)] reg2391 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2390 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2388 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2385 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2384 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2370 = (1'h0);
  reg [(5'h14):(1'h0)] reg2380 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2376 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2368 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2363 = (1'h0);
  reg [(5'h12):(1'h0)] reg2360 = (1'h0);
  reg [(5'h16):(1'h0)] reg2359 = (1'h0);
  reg [(5'h13):(1'h0)] reg2356 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2355 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2351 = (1'h0);
  reg [(4'hb):(1'h0)] reg2344 = (1'h0);
  reg [(5'h11):(1'h0)] reg2342 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2341 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2340 = (1'h0);
  reg [(3'h5):(1'h0)] reg2336 = (1'h0);
  reg [(5'h14):(1'h0)] reg2335 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2334 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2333 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2332 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2329 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2325 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2324 = (1'h0);
  reg [(4'hf):(1'h0)] reg2322 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2321 = (1'h0);
  reg [(4'he):(1'h0)] reg2320 = (1'h0);
  reg [(4'ha):(1'h0)] reg2318 = (1'h0);
  reg [(4'hb):(1'h0)] reg2316 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2311 = (1'h0);
  reg [(4'hf):(1'h0)] reg2308 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2307 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2305 = (1'h0);
  reg [(4'hd):(1'h0)] reg2304 = (1'h0);
  reg [(2'h3):(1'h0)] reg2302 = (1'h0);
  reg [(2'h3):(1'h0)] reg2301 = (1'h0);
  reg [(3'h4):(1'h0)] reg2299 = (1'h0);
  reg [(4'hb):(1'h0)] reg2297 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2295 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2293 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2289 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2287 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2286 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2285 = (1'h0);
  reg [(5'h14):(1'h0)] reg2284 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2279 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2275 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2260 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2271 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2270 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2268 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2265 = (1'h0);
  reg [(5'h17):(1'h0)] reg2264 = (1'h0);
  reg [(3'h5):(1'h0)] reg2263 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2262 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2258 = (1'h0);
  reg [(5'h10):(1'h0)] reg2255 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2252 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2250 = (1'h0);
  reg [(5'h12):(1'h0)] reg2249 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2248 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2244 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2243 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2242 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2241 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2240 = (1'h0);
  reg [(5'h13):(1'h0)] reg2238 = (1'h0);
  reg [(4'he):(1'h0)] reg2234 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2209 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2231 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2229 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2226 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2224 = (1'h0);
  reg [(5'h18):(1'h0)] reg2223 = (1'h0);
  reg [(4'hd):(1'h0)] reg2221 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2220 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2218 = (1'h0);
  reg [(5'h12):(1'h0)] reg2217 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2216 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2215 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2214 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2210 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2200 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2198 = (1'h0);
  reg [(3'h7):(1'h0)] reg2196 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2195 = (1'h0);
  reg [(3'h4):(1'h0)] reg2194 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2187 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2180 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2177 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2176 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2175 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2171 = (1'h0);
  reg [(5'h18):(1'h0)] reg2169 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2168 = (1'h0);
  reg [(4'ha):(1'h0)] reg2165 = (1'h0);
  reg [(5'h16):(1'h0)] reg2161 = (1'h0);
  reg [(3'h7):(1'h0)] reg2160 = (1'h0);
  reg [(4'hc):(1'h0)] reg2153 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2152 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2151 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2150 = (1'h0);
  reg [(5'h18):(1'h0)] reg2149 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2148 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2143 = (1'h0);
  reg [(2'h3):(1'h0)] reg2142 = (1'h0);
  reg [(3'h7):(1'h0)] reg2136 = (1'h0);
  reg [(5'h18):(1'h0)] reg2135 = (1'h0);
  reg [(5'h11):(1'h0)] reg2131 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2132 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2124 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2121 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2118 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2117 = (1'h0);
  reg [(3'h4):(1'h0)] reg2116 = (1'h0);
  reg [(5'h16):(1'h0)] reg2115 = (1'h0);
  reg [(3'h7):(1'h0)] reg2114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2111 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2110 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2109 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2108 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2107 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2104 = (1'h0);
  reg [(5'h18):(1'h0)] reg2098 = (1'h0);
  reg [(5'h19):(1'h0)] reg2097 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2095 = (1'h0);
  reg [(5'h10):(1'h0)] reg2094 = (1'h0);
  reg [(3'h5):(1'h0)] reg2093 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2091 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2088 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2082 = (1'h0);
  reg [(5'h17):(1'h0)] reg2075 = (1'h0);
  reg [(5'h15):(1'h0)] reg2078 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2073 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2071 = (1'h0);
  reg [(5'h14):(1'h0)] reg2070 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2067 = (1'h0);
  reg [(2'h2):(1'h0)] reg2066 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2065 = (1'h0);
  reg [(5'h11):(1'h0)] reg2064 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2063 = (1'h0);
  reg [(3'h7):(1'h0)] reg2062 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2060 = (1'h0);
  reg [(5'h10):(1'h0)] reg2057 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2056 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2054 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2053 = (1'h0);
  reg [(4'hd):(1'h0)] reg2052 = (1'h0);
  reg [(4'he):(1'h0)] reg2049 = (1'h0);
  reg [(4'h8):(1'h0)] reg2048 = (1'h0);
  reg [(4'hc):(1'h0)] reg2047 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2046 = (1'h0);
  reg [(5'h14):(1'h0)] reg2042 = (1'h0);
  reg [(4'h8):(1'h0)] reg2039 = (1'h0);
  reg [(4'hf):(1'h0)] reg2038 = (1'h0);
  reg [(4'hb):(1'h0)] reg2037 = (1'h0);
  reg [(5'h14):(1'h0)] reg2030 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2029 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2028 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2027 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2023 = (1'h0);
  reg [(5'h12):(1'h0)] reg2021 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2020 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2010 = (1'h0);
  reg [(4'hb):(1'h0)] reg2018 = (1'h0);
  reg [(4'ha):(1'h0)] reg2017 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2016 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2015 = (1'h0);
  reg [(5'h19):(1'h0)] reg2014 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2009 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2007 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2006 = (1'h0);
  reg [(5'h11):(1'h0)] reg2004 = (1'h0);
  reg [(2'h3):(1'h0)] reg2002 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2001 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2000 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1999 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1998 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1995 = (1'h0);
  reg [(5'h11):(1'h0)] reg1993 = (1'h0);
  reg [(5'h17):(1'h0)] reg1991 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1990 = (1'h0);
  reg [(4'ha):(1'h0)] reg1987 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1985 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1982 = (1'h0);
  reg [(5'h10):(1'h0)] reg1981 = (1'h0);
  reg [(5'h11):(1'h0)] reg1979 = (1'h0);
  reg [(3'h5):(1'h0)] reg1978 = (1'h0);
  reg [(4'h9):(1'h0)] reg1977 = (1'h0);
  reg [(5'h15):(1'h0)] reg1973 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1967 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1966 = (1'h0);
  reg [(5'h10):(1'h0)] reg1962 = (1'h0);
  reg [(5'h11):(1'h0)] reg1961 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1956 = (1'h0);
  reg [(2'h3):(1'h0)] reg1954 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1950 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1948 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1946 = (1'h0);
  reg [(4'hc):(1'h0)] reg1932 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1943 = (1'h0);
  reg [(5'h14):(1'h0)] reg1942 = (1'h0);
  reg [(5'h17):(1'h0)] reg1940 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1936 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1935 = (1'h0);
  reg [(4'hf):(1'h0)] reg1933 = (1'h0);
  reg [(5'h18):(1'h0)] reg1928 = (1'h0);
  reg [(4'hd):(1'h0)] reg1926 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1923 = (1'h0);
  reg [(4'hf):(1'h0)] reg1917 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1915 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1914 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1912 = (1'h0);
  reg [(5'h12):(1'h0)] reg1911 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1908 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1906 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1905 = (1'h0);
  reg [(3'h7):(1'h0)] reg1904 = (1'h0);
  reg [(5'h16):(1'h0)] reg1903 = (1'h0);
  reg [(4'hb):(1'h0)] reg1902 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1900 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1897 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1894 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1893 = (1'h0);
  reg [(4'hb):(1'h0)] reg1892 = (1'h0);
  reg [(5'h15):(1'h0)] reg1891 = (1'h0);
  reg [(5'h19):(1'h0)] reg1886 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1885 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1884 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1883 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1880 = (1'h0);
  reg [(4'hf):(1'h0)] reg1878 = (1'h0);
  reg [(3'h5):(1'h0)] reg1877 = (1'h0);
  reg [(4'h9):(1'h0)] reg1875 = (1'h0);
  reg [(3'h5):(1'h0)] reg1869 = (1'h0);
  reg [(2'h2):(1'h0)] reg1868 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1864 = (1'h0);
  reg [(4'h8):(1'h0)] reg1861 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1860 = (1'h0);
  reg [(3'h6):(1'h0)] reg1858 = (1'h0);
  reg [(4'h8):(1'h0)] reg1857 = (1'h0);
  reg [(3'h7):(1'h0)] reg1855 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1853 = (1'h0);
  reg [(5'h10):(1'h0)] reg1848 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1847 = (1'h0);
  reg [(5'h18):(1'h0)] reg1846 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1833 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1843 = (1'h0);
  reg [(4'h8):(1'h0)] reg1840 = (1'h0);
  reg [(4'hf):(1'h0)] reg1839 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1838 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1836 = (1'h0);
  reg [(2'h2):(1'h0)] reg1832 = (1'h0);
  reg [(5'h16):(1'h0)] reg1829 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1828 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg1826 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1825 = (1'h0);
  reg [(4'ha):(1'h0)] reg1824 = (1'h0);
  reg [(4'h9):(1'h0)] reg1822 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1819 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1818 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1816 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1814 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1811 = (1'h0);
  reg [(5'h12):(1'h0)] reg1808 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1806 = (1'h0);
  reg [(5'h11):(1'h0)] reg1804 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1803 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1800 = (1'h0);
  reg [(5'h1e):(1'h0)] reg1799 = (1'h0);
  reg [(5'h11):(1'h0)] reg1797 = (1'h0);
  reg [(3'h4):(1'h0)] reg1796 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1794 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1791 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1790 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1788 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1785 = (1'h0);
  reg [(4'hc):(1'h0)] reg1783 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1782 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1766 = (1'h0);
  reg [(5'h15):(1'h0)] reg1777 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1775 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1774 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1771 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1769 = (1'h0);
  reg [(4'hf):(1'h0)] reg1768 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2632 = (1'h0);
  reg [(2'h2):(1'h0)] reg2630 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2629 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2627 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2621 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2619 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2617 = (1'h0);
  reg [(4'h8):(1'h0)] reg2615 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2614 = (1'h0);
  reg [(5'h19):(1'h0)] reg2611 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2609 = (1'h0);
  reg [(5'h11):(1'h0)] reg2608 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2605 = (1'h0);
  reg [(5'h19):(1'h0)] reg2602 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2600 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2599 = (1'h0);
  reg [(4'hf):(1'h0)] reg2598 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2597 = (1'h0);
  reg [(4'h9):(1'h0)] reg2596 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2594 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2593 = (1'h0);
  reg [(5'h10):(1'h0)] reg2586 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2590 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2588 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2587 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2586 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2585 = (1'h0);
  reg [(5'h16):(1'h0)] reg2584 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2583 = (1'h0);
  reg [(2'h3):(1'h0)] reg2581 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2580 = (1'h0);
  reg [(2'h2):(1'h0)] reg2579 = (1'h0);
  reg [(5'h10):(1'h0)] reg2577 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2576 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2575 = (1'h0);
  reg [(5'h16):(1'h0)] reg2574 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2572 = (1'h0);
  reg [(4'hd):(1'h0)] reg2571 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2566 = (1'h0);
  reg [(4'hb):(1'h0)] reg2565 = (1'h0);
  reg [(3'h7):(1'h0)] reg2563 = (1'h0);
  reg [(5'h17):(1'h0)] reg2561 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2559 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2557 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2555 = (1'h0);
  reg [(3'h4):(1'h0)] reg2554 = (1'h0);
  reg [(5'h13):(1'h0)] reg2550 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2549 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2537 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2531 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2545 = (1'h0);
  reg [(2'h3):(1'h0)] reg2543 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2542 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2541 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2540 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2539 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2537 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2533 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2532 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2530 = (1'h0);
  reg [(2'h2):(1'h0)] reg2529 = (1'h0);
  reg [(2'h2):(1'h0)] reg2526 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2524 = (1'h0);
  reg [(5'h13):(1'h0)] reg2522 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2521 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2520 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2519 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2517 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2515 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2513 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2512 = (1'h0);
  reg [(4'ha):(1'h0)] reg2511 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2509 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2507 = (1'h0);
  reg [(5'h11):(1'h0)] reg2506 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2496 = (1'h0);
  reg [(3'h4):(1'h0)] reg2492 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2504 = (1'h0);
  reg [(5'h16):(1'h0)] reg2503 = (1'h0);
  reg [(3'h7):(1'h0)] reg2497 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2495 = (1'h0);
  reg [(4'ha):(1'h0)] reg2494 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2492 = (1'h0);
  reg [(5'h13):(1'h0)] reg2491 = (1'h0);
  reg [(4'h9):(1'h0)] reg2490 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2489 = (1'h0);
  reg [(5'h15):(1'h0)] reg2488 = (1'h0);
  reg [(4'h8):(1'h0)] reg2486 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2485 = (1'h0);
  reg [(3'h4):(1'h0)] reg2483 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2481 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2475 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2474 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2473 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2472 = (1'h0);
  reg [(5'h14):(1'h0)] reg2469 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2468 = (1'h0);
  reg [(5'h10):(1'h0)] reg2467 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2465 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2463 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2462 = (1'h0);
  reg [(5'h12):(1'h0)] reg2460 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2459 = (1'h0);
  reg [(4'ha):(1'h0)] reg2458 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2457 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2456 = (1'h0);
  reg [(5'h13):(1'h0)] reg2455 = (1'h0);
  reg [(4'hc):(1'h0)] reg2452 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2451 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2448 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2445 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2443 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2442 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2441 = (1'h0);
  reg [(4'h9):(1'h0)] reg2439 = (1'h0);
  reg [(5'h19):(1'h0)] reg2438 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar2435 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2434 = (1'h0);
  reg [(4'hc):(1'h0)] reg2432 = (1'h0);
  reg [(5'h17):(1'h0)] reg2431 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2430 = (1'h0);
  reg [(5'h14):(1'h0)] reg2429 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2428 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2427 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2426 = (1'h0);
  reg [(5'h10):(1'h0)] reg2425 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2424 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2423 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2421 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2419 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2416 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2415 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2412 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2411 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2406 = (1'h0);
  reg [(4'hb):(1'h0)] reg2405 = (1'h0);
  reg [(5'h13):(1'h0)] reg2394 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2402 = (1'h0);
  reg [(4'h9):(1'h0)] reg2399 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2398 = (1'h0);
  reg [(3'h4):(1'h0)] reg2397 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2394 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2392 = (1'h0);
  reg [(4'h8):(1'h0)] reg2389 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2387 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2386 = (1'h0);
  reg signed [(5'h1d):(1'h0)] forvar2383 = (1'h0);
  reg [(4'h9):(1'h0)] reg2382 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2365 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar2362 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2355 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2381 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2379 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2378 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2377 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2375 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2374 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2373 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2372 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2371 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2370 = (1'h0);
  reg [(5'h10):(1'h0)] reg2369 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2367 = (1'h0);
  reg [(5'h12):(1'h0)] reg2366 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar2365 = (1'h0);
  reg [(5'h17):(1'h0)] reg2364 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2362 = (1'h0);
  reg [(4'ha):(1'h0)] reg2361 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2357 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2354 = (1'h0);
  reg [(5'h18):(1'h0)] reg2353 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2352 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2350 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2349 = (1'h0);
  reg [(4'he):(1'h0)] reg2348 = (1'h0);
  reg [(5'h12):(1'h0)] reg2347 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2346 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2345 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2343 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2339 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2338 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2337 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2331 = (1'h0);
  reg [(5'h19):(1'h0)] reg2330 = (1'h0);
  reg [(5'h17):(1'h0)] reg2328 = (1'h0);
  reg [(4'hd):(1'h0)] reg2327 = (1'h0);
  reg [(3'h6):(1'h0)] reg2326 = (1'h0);
  reg [(4'ha):(1'h0)] reg2323 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2317 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2309 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2319 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2317 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2315 = (1'h0);
  reg [(4'hc):(1'h0)] reg2314 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2313 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2312 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2310 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar2309 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2306 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2303 = (1'h0);
  reg signed [(5'h1e):(1'h0)] forvar2300 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2298 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2296 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2294 = (1'h0);
  reg [(4'hd):(1'h0)] reg2292 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2291 = (1'h0);
  reg [(2'h2):(1'h0)] reg2290 = (1'h0);
  reg [(4'hd):(1'h0)] reg2288 = (1'h0);
  reg [(4'hf):(1'h0)] reg2283 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2282 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2281 = (1'h0);
  reg [(2'h2):(1'h0)] reg2280 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2278 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2277 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2276 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2274 = (1'h0);
  reg [(5'h17):(1'h0)] reg2273 = (1'h0);
  reg [(5'h17):(1'h0)] reg2272 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2269 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2267 = (1'h0);
  reg [(5'h14):(1'h0)] reg2266 = (1'h0);
  reg [(4'hd):(1'h0)] reg2261 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2260 = (1'h0);
  reg [(4'hc):(1'h0)] reg2259 = (1'h0);
  reg [(5'h14):(1'h0)] reg2257 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg2256 = (1'h0);
  reg [(5'h16):(1'h0)] forvar2254 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2253 = (1'h0);
  reg [(3'h7):(1'h0)] reg2251 = (1'h0);
  reg [(2'h3):(1'h0)] reg2247 = (1'h0);
  reg [(5'h14):(1'h0)] reg2246 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2245 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2239 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2237 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2236 = (1'h0);
  reg [(3'h5):(1'h0)] reg2235 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2223 = (1'h0);
  reg [(3'h7):(1'h0)] reg2233 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2232 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2230 = (1'h0);
  reg [(3'h5):(1'h0)] reg2228 = (1'h0);
  reg [(5'h16):(1'h0)] reg2227 = (1'h0);
  reg [(5'h1d):(1'h0)] reg2225 = (1'h0);
  reg [(2'h3):(1'h0)] reg2222 = (1'h0);
  reg [(4'hf):(1'h0)] reg2219 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2213 = (1'h0);
  reg [(3'h7):(1'h0)] reg2212 = (1'h0);
  reg [(5'h16):(1'h0)] reg2211 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2209 = (1'h0);
  reg [(4'ha):(1'h0)] reg2206 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2205 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2204 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2203 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2202 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2201 = (1'h0);
  reg [(5'h11):(1'h0)] reg2199 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar2197 = (1'h0);
  reg [(5'h14):(1'h0)] reg2193 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2192 = (1'h0);
  reg [(3'h4):(1'h0)] reg2191 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2190 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2189 = (1'h0);
  reg [(4'ha):(1'h0)] reg2188 = (1'h0);
  reg [(5'h15):(1'h0)] reg2186 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2185 = (1'h0);
  reg [(5'h1e):(1'h0)] reg2184 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2183 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2182 = (1'h0);
  reg [(4'he):(1'h0)] reg2181 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2179 = (1'h0);
  reg [(4'h8):(1'h0)] reg2178 = (1'h0);
  reg [(4'h9):(1'h0)] reg2174 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2173 = (1'h0);
  reg [(4'h8):(1'h0)] reg2172 = (1'h0);
  reg [(4'he):(1'h0)] reg2170 = (1'h0);
  reg [(4'hc):(1'h0)] reg2167 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar2166 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2164 = (1'h0);
  reg [(4'ha):(1'h0)] reg2163 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2162 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2159 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2158 = (1'h0);
  reg signed [(5'h1f):(1'h0)] reg2157 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2156 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2155 = (1'h0);
  reg [(4'hb):(1'h0)] reg2154 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2147 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2146 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2145 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2144 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2141 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2140 = (1'h0);
  reg [(3'h7):(1'h0)] reg2139 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg2138 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2137 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg2134 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2133 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2131 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2130 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2129 = (1'h0);
  reg [(4'hc):(1'h0)] reg2128 = (1'h0);
  reg [(4'hc):(1'h0)] reg2127 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2126 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2125 = (1'h0);
  reg [(5'h19):(1'h0)] reg2123 = (1'h0);
  reg [(5'h13):(1'h0)] reg2122 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2120 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2119 = (1'h0);
  reg [(5'h11):(1'h0)] reg2113 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2112 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2106 = (1'h0);
  reg [(5'h13):(1'h0)] reg2105 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2103 = (1'h0);
  reg [(5'h13):(1'h0)] reg2102 = (1'h0);
  reg [(4'hd):(1'h0)] reg2101 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2100 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2099 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2096 = (1'h0);
  reg [(5'h13):(1'h0)] reg2092 = (1'h0);
  reg [(5'h15):(1'h0)] reg2090 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2089 = (1'h0);
  reg [(5'h18):(1'h0)] reg2087 = (1'h0);
  reg [(5'h11):(1'h0)] reg2086 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2085 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2084 = (1'h0);
  reg [(3'h7):(1'h0)] reg2083 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar2073 = (1'h0);
  reg [(3'h5):(1'h0)] reg2072 = (1'h0);
  reg [(5'h1b):(1'h0)] reg2081 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2080 = (1'h0);
  reg [(5'h1c):(1'h0)] reg2079 = (1'h0);
  reg [(4'hf):(1'h0)] reg2077 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2076 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2075 = (1'h0);
  reg [(4'h9):(1'h0)] reg2074 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2072 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2069 = (1'h0);
  reg [(5'h19):(1'h0)] reg2068 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2061 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2059 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2058 = (1'h0);
  reg [(5'h16):(1'h0)] reg2055 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2051 = (1'h0);
  reg [(2'h3):(1'h0)] reg2050 = (1'h0);
  reg [(4'h9):(1'h0)] reg2045 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2044 = (1'h0);
  reg [(4'hd):(1'h0)] reg2041 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2040 = (1'h0);
  reg [(4'hc):(1'h0)] reg2036 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2035 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2034 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2033 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2032 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg2031 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2026 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2025 = (1'h0);
  reg [(5'h17):(1'h0)] reg2024 = (1'h0);
  reg [(4'hc):(1'h0)] reg2022 = (1'h0);
  reg [(5'h1f):(1'h0)] reg2019 = (1'h0);
  reg signed [(5'h1f):(1'h0)] forvar2015 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2005 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2013 = (1'h0);
  reg [(3'h4):(1'h0)] reg2012 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2011 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2010 = (1'h0);
  reg [(4'ha):(1'h0)] reg2008 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2005 = (1'h0);
  reg [(4'h9):(1'h0)] reg2003 = (1'h0);
  reg [(5'h19):(1'h0)] reg1997 = (1'h0);
  reg [(3'h6):(1'h0)] reg1996 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg1994 = (1'h0);
  reg [(5'h13):(1'h0)] reg1992 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1989 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1988 = (1'h0);
  reg [(3'h4):(1'h0)] reg1986 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1984 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1983 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1980 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1976 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1975 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1974 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1972 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1971 = (1'h0);
  reg [(4'h8):(1'h0)] reg1970 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1969 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1968 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1965 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1964 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1963 = (1'h0);
  reg [(4'ha):(1'h0)] reg1960 = (1'h0);
  reg [(5'h14):(1'h0)] reg1959 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1958 = (1'h0);
  reg [(5'h11):(1'h0)] reg1957 = (1'h0);
  reg [(4'h8):(1'h0)] reg1955 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1953 = (1'h0);
  reg [(4'h9):(1'h0)] reg1952 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1951 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1949 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1947 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1937 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1945 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1944 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1941 = (1'h0);
  reg [(5'h15):(1'h0)] reg1939 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1938 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1937 = (1'h0);
  reg [(3'h5):(1'h0)] reg1934 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1932 = (1'h0);
  reg [(4'hd):(1'h0)] reg1931 = (1'h0);
  reg [(4'ha):(1'h0)] reg1930 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1929 = (1'h0);
  reg [(3'h4):(1'h0)] reg1927 = (1'h0);
  reg [(3'h6):(1'h0)] reg1925 = (1'h0);
  reg signed [(5'h1d):(1'h0)] reg1924 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1922 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1921 = (1'h0);
  reg [(5'h13):(1'h0)] reg1920 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1919 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1918 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1916 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1913 = (1'h0);
  reg [(5'h11):(1'h0)] reg1910 = (1'h0);
  reg [(5'h1b):(1'h0)] reg1909 = (1'h0);
  reg [(5'h11):(1'h0)] reg1907 = (1'h0);
  reg [(4'hd):(1'h0)] reg1901 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1899 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1898 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1895 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1890 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1889 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1888 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1887 = (1'h0);
  reg [(5'h1f):(1'h0)] reg1882 = (1'h0);
  reg [(4'h9):(1'h0)] reg1881 = (1'h0);
  reg [(3'h4):(1'h0)] reg1879 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1876 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1874 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1873 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1872 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1871 = (1'h0);
  reg [(4'hc):(1'h0)] reg1870 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1867 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1866 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1865 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1863 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1859 = (1'h0);
  reg [(5'h10):(1'h0)] reg1856 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1853 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1862 = (1'h0);
  reg [(5'h1e):(1'h0)] forvar1859 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1856 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1854 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1852 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1851 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1850 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1849 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1847 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1826 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1845 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1844 = (1'h0);
  reg signed [(5'h1e):(1'h0)] reg1842 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1841 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1837 = (1'h0);
  reg [(3'h6):(1'h0)] reg1835 = (1'h0);
  reg [(5'h10):(1'h0)] reg1834 = (1'h0);
  reg [(4'he):(1'h0)] forvar1833 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1831 = (1'h0);
  reg [(2'h2):(1'h0)] reg1830 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1827 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1823 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1821 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1820 = (1'h0);
  reg signed [(5'h1c):(1'h0)] reg1817 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1815 = (1'h0);
  reg [(5'h1c):(1'h0)] reg1813 = (1'h0);
  reg [(3'h6):(1'h0)] reg1812 = (1'h0);
  reg [(5'h1d):(1'h0)] forvar1810 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1809 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1807 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1805 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1802 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1801 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1798 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1795 = (1'h0);
  reg [(5'h16):(1'h0)] reg1793 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1792 = (1'h0);
  reg [(5'h1d):(1'h0)] reg1789 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1787 = (1'h0);
  reg [(5'h10):(1'h0)] reg1786 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1784 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1781 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1780 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1779 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1770 = (1'h0);
  reg signed [(5'h1c):(1'h0)] forvar1767 = (1'h0);
  reg [(5'h18):(1'h0)] reg1778 = (1'h0);
  reg [(3'h6):(1'h0)] reg1776 = (1'h0);
  reg [(3'h4):(1'h0)] reg1773 = (1'h0);
  reg [(5'h12):(1'h0)] reg1772 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1770 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1767 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1766 = (1'h0);
  assign y = {wire2568,
                 wire2453,
                 wire2208,
                 wire2207,
                 wire2043,
                 wire1896,
                 wire1765,
                 reg2634,
                 reg2633,
                 reg2631,
                 reg2628,
                 reg2626,
                 reg2625,
                 reg2624,
                 reg2623,
                 reg2622,
                 reg2620,
                 reg2618,
                 reg2616,
                 reg2613,
                 reg2612,
                 reg2610,
                 reg2607,
                 reg2606,
                 reg2604,
                 reg2603,
                 reg2601,
                 reg2595,
                 reg2592,
                 reg2591,
                 reg2589,
                 reg2582,
                 reg2578,
                 reg2573,
                 reg2570,
                 reg2569,
                 reg2567,
                 reg2564,
                 reg2562,
                 reg2560,
                 reg2558,
                 reg2556,
                 reg2553,
                 reg2552,
                 reg2551,
                 reg2548,
                 reg2547,
                 reg2546,
                 reg2544,
                 reg2538,
                 reg2536,
                 reg2535,
                 reg2534,
                 reg2531,
                 reg2528,
                 reg2527,
                 reg2525,
                 reg2523,
                 reg2518,
                 reg2516,
                 reg2514,
                 reg2510,
                 reg2508,
                 reg2505,
                 reg2502,
                 reg2501,
                 reg2500,
                 reg2499,
                 reg2498,
                 reg2496,
                 reg2493,
                 reg2487,
                 reg2484,
                 reg2482,
                 reg2480,
                 reg2479,
                 reg2478,
                 reg2477,
                 reg2476,
                 reg2471,
                 reg2470,
                 reg2466,
                 reg2464,
                 reg2461,
                 reg2454,
                 reg2450,
                 reg2449,
                 reg2447,
                 reg2446,
                 reg2444,
                 reg2440,
                 reg2437,
                 reg2436,
                 reg2433,
                 reg2422,
                 reg2420,
                 reg2418,
                 reg2417,
                 reg2414,
                 reg2413,
                 reg2410,
                 reg2409,
                 reg2408,
                 reg2407,
                 reg2404,
                 reg2403,
                 reg2383,
                 reg2401,
                 reg2400,
                 reg2396,
                 reg2395,
                 reg2393,
                 reg2391,
                 reg2390,
                 reg2388,
                 reg2385,
                 reg2384,
                 reg2370,
                 reg2380,
                 reg2376,
                 reg2368,
                 reg2363,
                 reg2360,
                 reg2359,
                 reg2356,
                 reg2355,
                 reg2351,
                 reg2344,
                 reg2342,
                 reg2341,
                 reg2340,
                 reg2336,
                 reg2335,
                 reg2334,
                 reg2333,
                 reg2332,
                 reg2329,
                 reg2325,
                 reg2324,
                 reg2322,
                 reg2321,
                 reg2320,
                 reg2318,
                 reg2316,
                 reg2311,
                 reg2308,
                 reg2307,
                 reg2305,
                 reg2304,
                 reg2302,
                 reg2301,
                 reg2299,
                 reg2297,
                 reg2295,
                 reg2293,
                 reg2289,
                 reg2287,
                 reg2286,
                 reg2285,
                 reg2284,
                 reg2279,
                 reg2275,
                 reg2260,
                 reg2271,
                 reg2270,
                 reg2268,
                 reg2265,
                 reg2264,
                 reg2263,
                 reg2262,
                 reg2258,
                 reg2255,
                 reg2252,
                 reg2250,
                 reg2249,
                 reg2248,
                 reg2244,
                 reg2243,
                 reg2242,
                 reg2241,
                 reg2240,
                 reg2238,
                 reg2234,
                 reg2209,
                 reg2231,
                 reg2229,
                 reg2226,
                 reg2224,
                 reg2223,
                 reg2221,
                 reg2220,
                 reg2218,
                 reg2217,
                 reg2216,
                 reg2215,
                 reg2214,
                 reg2210,
                 reg2200,
                 reg2198,
                 reg2196,
                 reg2195,
                 reg2194,
                 reg2187,
                 reg2180,
                 reg2177,
                 reg2176,
                 reg2175,
                 reg2171,
                 reg2169,
                 reg2168,
                 reg2165,
                 reg2161,
                 reg2160,
                 reg2153,
                 reg2152,
                 reg2151,
                 reg2150,
                 reg2149,
                 reg2148,
                 reg2143,
                 reg2142,
                 reg2136,
                 reg2135,
                 reg2131,
                 reg2132,
                 reg2124,
                 reg2121,
                 reg2118,
                 reg2117,
                 reg2116,
                 reg2115,
                 reg2114,
                 reg2111,
                 reg2110,
                 reg2109,
                 reg2108,
                 reg2107,
                 reg2104,
                 reg2098,
                 reg2097,
                 reg2095,
                 reg2094,
                 reg2093,
                 reg2091,
                 reg2088,
                 reg2082,
                 reg2075,
                 reg2078,
                 reg2073,
                 reg2071,
                 reg2070,
                 reg2067,
                 reg2066,
                 reg2065,
                 reg2064,
                 reg2063,
                 reg2062,
                 reg2060,
                 reg2057,
                 reg2056,
                 reg2054,
                 reg2053,
                 reg2052,
                 reg2049,
                 reg2048,
                 reg2047,
                 reg2046,
                 reg2042,
                 reg2039,
                 reg2038,
                 reg2037,
                 reg2030,
                 reg2029,
                 reg2028,
                 reg2027,
                 reg2023,
                 reg2021,
                 reg2020,
                 reg2010,
                 reg2018,
                 reg2017,
                 reg2016,
                 reg2015,
                 reg2014,
                 reg2009,
                 reg2007,
                 reg2006,
                 reg2004,
                 reg2002,
                 reg2001,
                 reg2000,
                 reg1999,
                 reg1998,
                 reg1995,
                 reg1993,
                 reg1991,
                 reg1990,
                 reg1987,
                 reg1985,
                 reg1982,
                 reg1981,
                 reg1979,
                 reg1978,
                 reg1977,
                 reg1973,
                 reg1967,
                 reg1966,
                 reg1962,
                 reg1961,
                 reg1956,
                 reg1954,
                 reg1950,
                 reg1948,
                 reg1946,
                 reg1932,
                 reg1943,
                 reg1942,
                 reg1940,
                 reg1936,
                 reg1935,
                 reg1933,
                 reg1928,
                 reg1926,
                 reg1923,
                 reg1917,
                 reg1915,
                 reg1914,
                 reg1912,
                 reg1911,
                 reg1908,
                 reg1906,
                 reg1905,
                 reg1904,
                 reg1903,
                 reg1902,
                 reg1900,
                 reg1897,
                 reg1894,
                 reg1893,
                 reg1892,
                 reg1891,
                 reg1886,
                 reg1885,
                 reg1884,
                 reg1883,
                 reg1880,
                 reg1878,
                 reg1877,
                 reg1875,
                 reg1869,
                 reg1868,
                 reg1864,
                 reg1861,
                 reg1860,
                 reg1858,
                 reg1857,
                 reg1855,
                 reg1853,
                 reg1848,
                 reg1847,
                 reg1846,
                 reg1833,
                 reg1843,
                 reg1840,
                 reg1839,
                 reg1838,
                 reg1836,
                 reg1832,
                 reg1829,
                 reg1828,
                 reg1826,
                 reg1825,
                 reg1824,
                 reg1822,
                 reg1819,
                 reg1818,
                 reg1816,
                 reg1814,
                 reg1811,
                 reg1808,
                 reg1806,
                 reg1804,
                 reg1803,
                 reg1800,
                 reg1799,
                 reg1797,
                 reg1796,
                 reg1794,
                 reg1791,
                 reg1790,
                 reg1788,
                 reg1785,
                 reg1783,
                 reg1782,
                 reg1766,
                 reg1777,
                 reg1775,
                 reg1774,
                 reg1771,
                 reg1769,
                 reg1768,
                 reg2632,
                 reg2630,
                 reg2629,
                 reg2627,
                 reg2621,
                 reg2619,
                 reg2617,
                 reg2615,
                 reg2614,
                 reg2611,
                 reg2609,
                 reg2608,
                 forvar2605,
                 reg2602,
                 reg2600,
                 reg2599,
                 reg2598,
                 reg2597,
                 reg2596,
                 reg2594,
                 reg2593,
                 reg2586,
                 reg2590,
                 reg2588,
                 reg2587,
                 forvar2586,
                 reg2585,
                 reg2584,
                 reg2583,
                 reg2581,
                 reg2580,
                 reg2579,
                 reg2577,
                 reg2576,
                 reg2575,
                 reg2574,
                 forvar2572,
                 reg2571,
                 reg2566,
                 reg2565,
                 reg2563,
                 reg2561,
                 forvar2559,
                 reg2557,
                 reg2555,
                 reg2554,
                 reg2550,
                 reg2549,
                 reg2537,
                 forvar2531,
                 reg2545,
                 reg2543,
                 reg2542,
                 reg2541,
                 reg2540,
                 reg2539,
                 forvar2537,
                 reg2533,
                 reg2532,
                 reg2530,
                 reg2529,
                 reg2526,
                 reg2524,
                 reg2522,
                 reg2521,
                 forvar2520,
                 reg2519,
                 reg2517,
                 reg2515,
                 forvar2513,
                 forvar2512,
                 reg2511,
                 reg2509,
                 reg2507,
                 reg2506,
                 forvar2496,
                 reg2492,
                 reg2504,
                 reg2503,
                 reg2497,
                 reg2495,
                 reg2494,
                 forvar2492,
                 reg2491,
                 reg2490,
                 reg2489,
                 reg2488,
                 reg2486,
                 reg2485,
                 reg2483,
                 reg2481,
                 reg2475,
                 forvar2474,
                 reg2473,
                 reg2472,
                 reg2469,
                 reg2468,
                 reg2467,
                 forvar2465,
                 forvar2463,
                 reg2462,
                 reg2460,
                 reg2459,
                 reg2458,
                 forvar2457,
                 forvar2456,
                 reg2455,
                 reg2452,
                 reg2451,
                 reg2448,
                 reg2445,
                 reg2443,
                 reg2442,
                 reg2441,
                 reg2439,
                 reg2438,
                 forvar2435,
                 reg2434,
                 reg2432,
                 reg2431,
                 reg2430,
                 reg2429,
                 reg2428,
                 reg2427,
                 reg2426,
                 reg2425,
                 forvar2424,
                 reg2423,
                 reg2421,
                 reg2419,
                 reg2416,
                 reg2415,
                 reg2412,
                 forvar2411,
                 reg2406,
                 reg2405,
                 reg2394,
                 reg2402,
                 reg2399,
                 reg2398,
                 reg2397,
                 forvar2394,
                 reg2392,
                 reg2389,
                 reg2387,
                 reg2386,
                 forvar2383,
                 reg2382,
                 reg2365,
                 forvar2362,
                 forvar2355,
                 reg2381,
                 forvar2379,
                 reg2378,
                 forvar2377,
                 reg2375,
                 reg2374,
                 reg2373,
                 reg2372,
                 reg2371,
                 forvar2370,
                 reg2369,
                 reg2367,
                 reg2366,
                 forvar2365,
                 reg2364,
                 reg2362,
                 reg2361,
                 reg2358,
                 reg2357,
                 reg2354,
                 reg2353,
                 reg2352,
                 reg2350,
                 forvar2349,
                 reg2348,
                 reg2347,
                 reg2346,
                 reg2345,
                 forvar2343,
                 reg2339,
                 reg2338,
                 forvar2337,
                 forvar2331,
                 reg2330,
                 reg2328,
                 reg2327,
                 reg2326,
                 reg2323,
                 reg2317,
                 reg2309,
                 reg2319,
                 forvar2317,
                 reg2315,
                 reg2314,
                 reg2313,
                 reg2312,
                 reg2310,
                 forvar2309,
                 reg2306,
                 forvar2303,
                 forvar2300,
                 reg2298,
                 reg2296,
                 reg2294,
                 reg2292,
                 reg2291,
                 reg2290,
                 reg2288,
                 reg2283,
                 forvar2282,
                 reg2281,
                 reg2280,
                 reg2278,
                 reg2277,
                 reg2276,
                 forvar2274,
                 reg2273,
                 reg2272,
                 reg2269,
                 reg2267,
                 reg2266,
                 reg2261,
                 forvar2260,
                 reg2259,
                 reg2257,
                 reg2256,
                 forvar2254,
                 reg2253,
                 reg2251,
                 reg2247,
                 reg2246,
                 reg2245,
                 reg2239,
                 reg2237,
                 reg2236,
                 reg2235,
                 forvar2223,
                 reg2233,
                 reg2232,
                 reg2230,
                 reg2228,
                 reg2227,
                 reg2225,
                 reg2222,
                 reg2219,
                 reg2213,
                 reg2212,
                 reg2211,
                 forvar2209,
                 reg2206,
                 forvar2205,
                 forvar2204,
                 reg2203,
                 reg2202,
                 reg2201,
                 reg2199,
                 forvar2197,
                 reg2193,
                 reg2192,
                 reg2191,
                 forvar2190,
                 reg2189,
                 reg2188,
                 reg2186,
                 reg2185,
                 reg2184,
                 reg2183,
                 forvar2182,
                 reg2181,
                 reg2179,
                 reg2178,
                 reg2174,
                 reg2173,
                 reg2172,
                 reg2170,
                 reg2167,
                 forvar2166,
                 reg2164,
                 reg2163,
                 reg2162,
                 reg2159,
                 forvar2158,
                 reg2157,
                 reg2156,
                 reg2155,
                 reg2154,
                 forvar2147,
                 reg2146,
                 forvar2145,
                 reg2144,
                 reg2141,
                 reg2140,
                 reg2139,
                 reg2138,
                 reg2137,
                 reg2134,
                 reg2133,
                 forvar2131,
                 reg2130,
                 reg2129,
                 reg2128,
                 reg2127,
                 reg2126,
                 reg2125,
                 reg2123,
                 reg2122,
                 reg2120,
                 reg2119,
                 reg2113,
                 reg2112,
                 reg2106,
                 reg2105,
                 forvar2103,
                 reg2102,
                 reg2101,
                 reg2100,
                 forvar2099,
                 forvar2096,
                 reg2092,
                 reg2090,
                 reg2089,
                 reg2087,
                 reg2086,
                 forvar2085,
                 forvar2084,
                 reg2083,
                 forvar2073,
                 reg2072,
                 reg2081,
                 reg2080,
                 reg2079,
                 reg2077,
                 reg2076,
                 forvar2075,
                 reg2074,
                 forvar2072,
                 reg2069,
                 reg2068,
                 reg2061,
                 reg2059,
                 forvar2058,
                 reg2055,
                 forvar2051,
                 reg2050,
                 reg2045,
                 forvar2044,
                 reg2041,
                 reg2040,
                 reg2036,
                 forvar2035,
                 reg2034,
                 reg2033,
                 forvar2032,
                 reg2031,
                 reg2026,
                 reg2025,
                 reg2024,
                 reg2022,
                 reg2019,
                 forvar2015,
                 reg2005,
                 reg2013,
                 reg2012,
                 reg2011,
                 forvar2010,
                 reg2008,
                 forvar2005,
                 reg2003,
                 reg1997,
                 reg1996,
                 reg1994,
                 reg1992,
                 reg1989,
                 reg1988,
                 reg1986,
                 forvar1984,
                 forvar1983,
                 reg1980,
                 reg1976,
                 reg1975,
                 reg1974,
                 reg1972,
                 reg1971,
                 reg1970,
                 reg1969,
                 forvar1968,
                 forvar1965,
                 reg1964,
                 reg1963,
                 reg1960,
                 reg1959,
                 reg1958,
                 reg1957,
                 reg1955,
                 reg1953,
                 reg1952,
                 forvar1951,
                 reg1949,
                 forvar1947,
                 reg1937,
                 reg1945,
                 reg1944,
                 reg1941,
                 reg1939,
                 reg1938,
                 forvar1937,
                 reg1934,
                 forvar1932,
                 reg1931,
                 reg1930,
                 reg1929,
                 reg1927,
                 reg1925,
                 reg1924,
                 forvar1922,
                 reg1921,
                 reg1920,
                 reg1919,
                 reg1918,
                 reg1916,
                 forvar1913,
                 reg1910,
                 reg1909,
                 reg1907,
                 reg1901,
                 forvar1899,
                 forvar1898,
                 reg1895,
                 reg1890,
                 forvar1889,
                 reg1888,
                 reg1887,
                 reg1882,
                 reg1881,
                 reg1879,
                 reg1876,
                 reg1874,
                 reg1873,
                 reg1872,
                 reg1871,
                 reg1870,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1863,
                 reg1859,
                 reg1856,
                 forvar1853,
                 reg1862,
                 forvar1859,
                 forvar1856,
                 reg1854,
                 reg1852,
                 reg1851,
                 reg1850,
                 reg1849,
                 forvar1847,
                 forvar1826,
                 reg1845,
                 reg1844,
                 reg1842,
                 reg1841,
                 reg1837,
                 reg1835,
                 reg1834,
                 forvar1833,
                 reg1831,
                 reg1830,
                 reg1827,
                 reg1823,
                 reg1821,
                 reg1820,
                 reg1817,
                 reg1815,
                 reg1813,
                 reg1812,
                 forvar1810,
                 reg1809,
                 reg1807,
                 reg1805,
                 reg1802,
                 reg1801,
                 reg1798,
                 forvar1795,
                 reg1793,
                 forvar1792,
                 reg1789,
                 reg1787,
                 reg1786,
                 forvar1784,
                 reg1781,
                 forvar1780,
                 forvar1779,
                 reg1770,
                 forvar1767,
                 reg1778,
                 reg1776,
                 reg1773,
                 reg1772,
                 forvar1770,
                 reg1767,
                 forvar1766,
                 (1'h0)};
  assign wire1765 = ((~(($signed((8'hb2)) != wire1760[(4'h8):(4'h8)]) ^~ $signed($unsigned(wire1760)))) - $unsigned((!$signed({wire1762,
                        (8'hbc),
                        wire1763}))));
  always
    @(posedge clk) begin
      if ((wire1765[(2'h2):(1'h1)] >> wire1762))
        begin
          for (forvar1766 = (1'h0); (forvar1766 < (3'h6)); forvar1766 = (forvar1766 + (1'h1)))
            begin
              reg1767 = $unsigned(wire1763[(1'h0):(1'h0)]);
              reg1768 <= {(wire1764[(3'h4):(2'h3)] << $signed(reg1767)),
                  forvar1766,
                  ((~&$unsigned(wire1763)) ? (8'hb4) : (8'ha3))};
              reg1769 <= {(wire1760[(4'ha):(3'h6)] ~^ $unsigned(((wire1761 ?
                      wire1760 : forvar1766) * $signed((8'ha5))))),
                  (-$signed((^~(~wire1763)))),
                  (~$unsigned((reg1768[(2'h3):(1'h1)] ?
                      wire1761[(4'hf):(4'hf)] : (^wire1764))))};
            end
          for (forvar1770 = (1'h0); (forvar1770 < (3'h4)); forvar1770 = (forvar1770 + (1'h1)))
            begin
              reg1771 <= (-forvar1766[(5'h16):(3'h5)]);
              reg1772 = ((7'h52) ?
                  (({((7'h4e) ? reg1768 : wire1762)} && ($unsigned(wire1762) ?
                      (reg1769 & forvar1770) : $unsigned(wire1761))) ^~ reg1769[(1'h1):(1'h1)]) : {(reg1771[(1'h0):(1'h0)] ?
                          (~^$unsigned((7'h51))) : ((reg1769 == wire1761) < wire1764[(5'h13):(4'hb)]))});
              reg1773 = $signed($signed($unsigned(($unsigned(forvar1766) | $unsigned(reg1768)))));
              reg1774 <= $signed(reg1768);
            end
          reg1775 <= $signed((((reg1767 == $signed((7'h57))) || reg1774[(4'h8):(1'h1)]) ?
              (8'ha7) : ((+reg1769[(4'hd):(2'h3)]) ?
                  $signed((wire1763 ?
                      reg1772 : wire1764)) : $signed((reg1773 - wire1763)))));
          if ($signed((((7'h44) ? $unsigned($unsigned(forvar1766)) : wire1764) ?
              wire1762[(3'h7):(3'h6)] : $unsigned((~^reg1771[(2'h3):(1'h1)])))))
            begin
              reg1776 = (~($unsigned($unsigned((8'hbe))) >>> (^($unsigned(reg1775) + (reg1769 == wire1760)))));
              reg1777 <= (+(($signed(reg1767) > (+$signed(reg1769))) >> wire1760[(1'h0):(1'h0)]));
            end
          else
            begin
              reg1777 <= (~|(8'hb1));
              reg1778 = $signed((~&reg1771[(1'h0):(1'h0)]));
            end
        end
      else
        begin
          reg1766 <= (!((^~{(+wire1762),
              reg1775[(2'h3):(1'h1)]}) ^ $signed(((^wire1763) ?
              reg1778 : wire1765))));
          for (forvar1767 = (1'h0); (forvar1767 < (3'h4)); forvar1767 = (forvar1767 + (1'h1)))
            begin
              reg1768 <= $unsigned({(!(((7'h40) ^ reg1767) ?
                      ((8'hbd) & forvar1770) : (wire1763 <= wire1764)))});
              reg1770 = reg1773[(1'h1):(1'h1)];
              reg1771 <= $unsigned(wire1764);
              reg1774 <= $signed(reg1766);
              reg1776 = wire1763[(1'h0):(1'h0)];
            end
        end
      for (forvar1779 = (1'h0); (forvar1779 < (2'h2)); forvar1779 = (forvar1779 + (1'h1)))
        begin
          for (forvar1780 = (1'h0); (forvar1780 < (2'h3)); forvar1780 = (forvar1780 + (1'h1)))
            begin
              reg1781 = {wire1765};
              reg1782 <= $signed((~$signed({$unsigned(reg1776),
                  $signed((8'hba))})));
              reg1783 <= wire1760[(4'hc):(2'h2)];
            end
          for (forvar1784 = (1'h0); (forvar1784 < (2'h3)); forvar1784 = (forvar1784 + (1'h1)))
            begin
              reg1785 <= ($unsigned($signed($unsigned((+reg1769)))) == (+$signed({$signed(forvar1779),
                  reg1775[(1'h1):(1'h0)],
                  $unsigned(wire1762)})));
              reg1786 = (wire1764[(5'h14):(5'h11)] != (forvar1766[(4'hc):(3'h4)] <= ({(wire1763 ?
                      (7'h4d) : (8'had))} >= $unsigned($signed(reg1768)))));
              reg1787 = (~|forvar1766[(5'h1a):(4'ha)]);
              reg1788 <= $signed((($unsigned({reg1768}) ?
                  reg1785 : wire1764) ~^ $signed(wire1765[(1'h1):(1'h0)])));
              reg1789 = reg1782;
            end
          reg1790 <= $unsigned(($signed({(~wire1765),
                  (reg1766 ? reg1767 : forvar1779)}) ?
              $signed(reg1768[(3'h4):(1'h1)]) : (|((wire1765 && forvar1779) ?
                  (wire1760 * (8'ha9)) : {reg1770, wire1760, wire1761}))));
          reg1791 <= ($signed($signed(reg1782)) ?
              (((|$signed(reg1785)) ?
                  reg1775[(1'h1):(1'h0)] : $signed(reg1790)) | $signed($unsigned($unsigned(reg1770)))) : reg1776[(2'h3):(1'h1)]);
          for (forvar1792 = (1'h0); (forvar1792 < (1'h0)); forvar1792 = (forvar1792 + (1'h1)))
            begin
              reg1793 = $unsigned(((~((~^reg1787) >> wire1760[(4'hd):(3'h7)])) ?
                  reg1770 : $unsigned((reg1771 <= reg1778[(3'h6):(3'h5)]))));
            end
          reg1794 <= $unsigned(reg1777[(2'h3):(2'h3)]);
          for (forvar1795 = (1'h0); (forvar1795 < (3'h4)); forvar1795 = (forvar1795 + (1'h1)))
            begin
              reg1796 <= reg1794;
              reg1797 <= (reg1781 >> $signed(reg1789));
            end
        end
      reg1798 = (7'h4e);
      reg1799 <= ({(8'hac),
              {reg1781, reg1766[(1'h0):(1'h0)], reg1788[(5'h19):(3'h4)]},
              reg1794[(5'h12):(3'h4)]} ?
          (($signed((7'h4a)) > (reg1798 * (~&forvar1770))) | reg1774) : reg1773);
      if ((reg1774[(1'h0):(1'h0)] | reg1775))
        begin
          reg1800 <= {$signed($unsigned(((reg1786 | reg1770) ?
                  (reg1777 << reg1793) : (reg1769 ? forvar1770 : reg1772)))),
              ((!$unsigned(((7'h58) & reg1791))) > wire1760[(4'h8):(4'h8)]),
              {(~$signed(reg1799))}};
        end
      else
        begin
          if ($unsigned(({($unsigned((8'hbd)) ? reg1786 : (~&reg1772)),
              $signed({reg1776, reg1771}),
              ((~^reg1769) ?
                  (reg1790 >>> reg1790) : forvar1784)} <<< reg1797[(3'h5):(1'h0)])))
            begin
              reg1801 = (($signed((forvar1795 ?
                  $unsigned(reg1796) : (^~reg1781))) && {(reg1768 ?
                      forvar1792[(4'he):(3'h4)] : reg1769[(1'h0):(1'h0)]),
                  reg1771[(1'h1):(1'h1)]}) ~^ $unsigned((-$signed(reg1794))));
              reg1802 = wire1764[(3'h5):(2'h3)];
              reg1803 <= $signed((^~$signed((|reg1783[(3'h6):(1'h1)]))));
              reg1804 <= ($signed((7'h47)) && {reg1771[(3'h7):(3'h5)],
                  (((~wire1762) ? {reg1782, reg1796, reg1788} : (~&reg1769)) ?
                      (!reg1799[(5'h1e):(4'he)]) : {reg1797[(3'h7):(3'h6)],
                          $unsigned((8'hb7))})});
              reg1805 = $unsigned((reg1800 ?
                  ((reg1781[(1'h0):(1'h0)] ?
                          ((7'h52) ? reg1785 : reg1772) : wire1762) ?
                      (~&{(8'ha0),
                          reg1798,
                          forvar1770}) : reg1775) : (+$signed(reg1773))));
            end
          else
            begin
              reg1801 = (|reg1801[(5'h12):(4'ha)]);
              reg1803 <= reg1788;
              reg1805 = reg1775;
              reg1806 <= (~|{((((8'ha6) ? reg1799 : reg1776) ?
                          {wire1760} : forvar1779[(3'h6):(2'h3)]) ?
                      {(~^reg1775)} : (8'hbe)),
                  ((+reg1773[(1'h1):(1'h1)]) ?
                      (~&$unsigned((8'hb4))) : reg1767)});
              reg1807 = forvar1795;
              reg1808 <= $signed({$signed((^(reg1801 >> reg1796))), reg1800});
            end
          reg1809 = reg1783[(4'h8):(2'h3)];
          for (forvar1810 = (1'h0); (forvar1810 < (1'h0)); forvar1810 = (forvar1810 + (1'h1)))
            begin
              reg1811 <= reg1773[(2'h3):(2'h3)];
              reg1812 = $signed(((^($signed((8'hb0)) ?
                      $signed(reg1794) : (!(8'hbd)))) ?
                  reg1781 : (reg1767[(3'h4):(1'h0)] <= $unsigned(reg1788))));
              reg1813 = {((($signed(reg1774) ?
                          $signed((7'h53)) : (reg1783 | reg1800)) ?
                      $signed(reg1766) : reg1768) >>> (~^(reg1798[(4'he):(4'h8)] || $signed(reg1778)))),
                  $signed(reg1772[(4'he):(3'h6)]),
                  (reg1808 >> (!(~&wire1760)))};
              reg1814 <= (reg1807 * $unsigned(({(reg1777 ? (7'h4c) : wire1762),
                      reg1804} ?
                  forvar1779[(5'h13):(5'h12)] : ($unsigned(reg1766) ?
                      reg1812 : {reg1802, reg1775}))));
              reg1815 = $unsigned((reg1814[(4'hb):(4'ha)] ?
                  forvar1810 : forvar1766));
              reg1816 <= ($signed(({(^~forvar1810), forvar1792, (^~reg1773)} ?
                  (+(~|reg1768)) : reg1793[(4'he):(3'h5)])) && ($signed(((+reg1808) ?
                      {reg1799} : $unsigned(reg1766))) ?
                  {{$signed(wire1765)}} : $unsigned($signed((reg1766 ?
                      reg1797 : reg1768)))));
              reg1817 = (reg1789[(3'h6):(3'h6)] ?
                  (~reg1813[(4'he):(4'hd)]) : reg1789);
            end
          reg1818 <= (($unsigned($signed(reg1791)) <<< ((+wire1765[(2'h2):(1'h0)]) | (wire1764[(5'h14):(5'h14)] ?
              reg1787[(5'h16):(5'h12)] : (reg1793 ?
                  reg1774 : reg1788)))) - $unsigned(reg1783[(2'h2):(2'h2)]));
          reg1819 <= (~|((wire1764[(4'hd):(1'h0)] ?
              (reg1768 + reg1800[(5'h13):(3'h7)]) : (forvar1792[(4'hc):(3'h7)] * (reg1774 + forvar1767))) < $signed((~^reg1803))));
          reg1820 = $signed($unsigned((($signed(reg1785) <= (forvar1779 ?
                  reg1802 : reg1813)) ?
              (|(-(8'h9e))) : $signed(forvar1795))));
        end
      reg1821 = $signed(($signed($unsigned((reg1815 ~^ reg1799))) ?
          wire1762 : $unsigned(reg1796)));
    end
  always
    @(posedge clk) begin
      reg1822 <= reg1788[(5'h19):(3'h7)];
      reg1823 = (({(!(&wire1760)),
              reg1785[(1'h1):(1'h0)],
              (reg1808[(4'he):(2'h3)] ?
                  $unsigned(reg1797) : $unsigned(reg1785))} ~^ (&reg1791[(2'h3):(1'h0)])) ?
          wire1761[(4'h8):(4'h8)] : $signed(($unsigned($unsigned(wire1765)) ?
              {$unsigned(reg1816),
                  $unsigned(reg1769),
                  wire1764} : {(wire1762 | wire1765),
                  $unsigned(reg1799),
                  (reg1766 | wire1765)})));
      reg1824 <= ($signed((((wire1764 < reg1771) <<< (reg1797 ?
          reg1822 : reg1816)) < $unsigned(wire1760[(2'h3):(2'h2)]))) + (!$unsigned((wire1764 >= $unsigned(wire1763)))));
      reg1825 <= reg1824;
      if ($signed((reg1794[(4'hd):(1'h0)] ?
          ($unsigned((reg1782 + reg1766)) ?
              (reg1800[(5'h1a):(5'h17)] == $unsigned(wire1765)) : ((reg1796 ?
                  wire1764 : reg1818) ~^ $unsigned(reg1824))) : ($unsigned($unsigned(reg1799)) ?
              (^{reg1799, reg1808, reg1774}) : $unsigned(wire1763)))))
        begin
          reg1826 <= $signed(reg1811[(4'hc):(2'h3)]);
          if (reg1796[(3'h4):(1'h1)])
            begin
              reg1827 = $unsigned(wire1765);
              reg1828 <= reg1783;
              reg1829 <= ((~^((reg1769 ? $unsigned((8'hac)) : (7'h55)) ?
                      (reg1771[(1'h1):(1'h1)] ^~ (reg1794 <= reg1803)) : $unsigned(reg1808[(4'h8):(2'h2)]))) ?
                  $unsigned((reg1814[(4'hb):(2'h3)] ?
                      $signed(reg1825) : wire1765[(1'h1):(1'h0)])) : reg1775[(2'h2):(1'h1)]);
              reg1830 = $signed($unsigned($signed((+$signed(reg1829)))));
              reg1831 = $signed($signed($unsigned(((+wire1762) ?
                  reg1785 : {reg1788, reg1829}))));
              reg1832 <= reg1823[(3'h4):(1'h0)];
            end
          else
            begin
              reg1828 <= (|($unsigned({$unsigned(reg1811),
                  $signed((8'hb1))}) < reg1766));
            end
          for (forvar1833 = (1'h0); (forvar1833 < (3'h6)); forvar1833 = (forvar1833 + (1'h1)))
            begin
              reg1834 = wire1761;
              reg1835 = reg1814;
              reg1836 <= (!(+(reg1782 ?
                  $signed(reg1808[(4'hb):(4'hb)]) : ({reg1803, wire1764} ?
                      $signed(reg1835) : {reg1775, reg1799, reg1826}))));
              reg1837 = reg1797[(2'h3):(1'h1)];
              reg1838 <= reg1794;
            end
          if ((~&($signed(($unsigned(reg1790) ?
                  (reg1836 <<< (8'hac)) : $signed(reg1777))) ?
              (-$unsigned((reg1834 ?
                  reg1783 : reg1808))) : (!((~|reg1768) - $signed(reg1785))))))
            begin
              reg1839 <= {$signed(wire1765[(1'h0):(1'h0)]),
                  reg1774[(3'h4):(2'h2)],
                  reg1825[(3'h5):(1'h1)]};
              reg1840 <= reg1785[(2'h2):(1'h1)];
              reg1841 = ({reg1808[(4'hd):(1'h0)]} ?
                  ($unsigned(reg1839[(4'hb):(3'h6)]) > (|(!reg1797[(4'hd):(3'h6)]))) : reg1838[(5'h17):(5'h12)]);
              reg1842 = {reg1814[(1'h1):(1'h1)],
                  (reg1806 ^ (&($unsigned(reg1814) ?
                      reg1837[(3'h6):(1'h0)] : (reg1819 | reg1769)))),
                  $signed($unsigned({(7'h40), $unsigned(reg1794), (8'ha8)}))};
              reg1843 <= $unsigned(reg1790[(2'h3):(2'h3)]);
            end
          else
            begin
              reg1841 = reg1791[(1'h0):(1'h0)];
              reg1842 = {$signed(reg1837[(3'h6):(3'h4)]),
                  (((+reg1808) ?
                      (~|(~^reg1799)) : reg1816[(4'hb):(2'h3)]) != reg1768)};
              reg1844 = $signed($unsigned(({$signed(reg1788)} ?
                  $unsigned((reg1790 ~^ reg1842)) : ((~reg1774) ?
                      {(8'hbe)} : reg1804[(3'h7):(3'h5)]))));
              reg1845 = reg1843[(4'ha):(2'h2)];
            end
        end
      else
        begin
          for (forvar1826 = (1'h0); (forvar1826 < (2'h2)); forvar1826 = (forvar1826 + (1'h1)))
            begin
              reg1827 = reg1806;
            end
          if (((~$unsigned({((7'h44) >>> reg1788)})) ?
              (8'had) : {(wire1761[(5'h1d):(4'hf)] ^~ ($unsigned((8'hb8)) ?
                      $signed(reg1838) : reg1826))}))
            begin
              reg1830 = (~|reg1803);
              reg1832 <= (($signed(((~^reg1799) <<< (reg1832 ?
                          reg1826 : wire1762))) ?
                      reg1829[(3'h7):(3'h5)] : (($unsigned(reg1790) ?
                              reg1840[(3'h5):(1'h1)] : (reg1843 >>> reg1790)) ?
                          ((~^reg1831) ?
                              (reg1838 + wire1765) : reg1791[(2'h2):(2'h2)]) : (7'h55))) ?
                  reg1838[(1'h0):(1'h0)] : reg1822[(3'h5):(3'h4)]);
            end
          else
            begin
              reg1828 <= reg1806[(5'h18):(2'h2)];
              reg1829 <= (^~(($unsigned(reg1841[(4'ha):(2'h2)]) == ((reg1803 <= reg1814) ?
                  $unsigned(reg1841) : ((8'hb6) ?
                      reg1774 : reg1804))) + (8'hb0)));
            end
          reg1833 <= reg1816[(5'h1b):(5'h14)];
          reg1836 <= (|(~^(reg1829 ?
              (~$signed((8'ha2))) : (reg1768 ?
                  reg1768[(4'he):(1'h0)] : $unsigned(reg1804)))));
        end
      if ((reg1836[(3'h6):(3'h4)] ?
          ((~&$signed($signed(wire1764))) ~^ $signed($unsigned($unsigned((7'h56))))) : reg1845))
        begin
          reg1846 <= $unsigned(($signed($unsigned((reg1804 ^ reg1814))) ?
              $unsigned(reg1766[(3'h4):(1'h1)]) : (wire1762[(3'h7):(2'h3)] && $unsigned((^~reg1844)))));
          reg1847 <= reg1790;
        end
      else
        begin
          reg1846 <= $unsigned(($signed($unsigned((8'hbf))) ?
              {((wire1760 ? reg1783 : (8'h9d)) ?
                      $unsigned(reg1800) : $unsigned(reg1823)),
                  {reg1818, $unsigned(reg1844), (reg1835 <= (7'h58))},
                  ($unsigned(wire1765) << (~&reg1790))} : (^reg1846)));
          for (forvar1847 = (1'h0); (forvar1847 < (1'h0)); forvar1847 = (forvar1847 + (1'h1)))
            begin
              reg1848 <= $unsigned($unsigned($signed(($unsigned(reg1791) < (-reg1804)))));
              reg1849 = $unsigned({$unsigned(reg1777),
                  (((reg1844 ?
                      reg1811 : wire1762) >= $unsigned(reg1814)) || $signed((8'hb2)))});
              reg1850 = reg1831[(4'ha):(4'ha)];
              reg1851 = reg1832[(1'h1):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg1852 = $signed(reg1811[(3'h4):(2'h3)]);
      if ((reg1822[(1'h0):(1'h0)] ?
          ($unsigned(((wire1761 <<< reg1852) || (reg1847 ?
              (8'hb3) : reg1766))) * reg1782[(5'h16):(3'h5)]) : reg1777[(4'he):(1'h0)]))
        begin
          reg1853 <= ($unsigned((($unsigned(reg1847) ?
                  $signed(reg1839) : $signed(reg1799)) ?
              ($signed(reg1852) ?
                  (reg1803 ?
                      reg1796 : reg1804) : (~|reg1822)) : reg1852)) ^ ($signed({$unsigned(reg1808),
                  reg1782,
                  (reg1822 ? reg1832 : reg1840)}) ?
              (8'ha8) : reg1804[(4'h9):(2'h2)]));
          reg1854 = $signed(reg1782[(4'hc):(3'h5)]);
          reg1855 <= $signed($signed(($signed(reg1811[(3'h6):(1'h1)]) ?
              reg1782[(5'h13):(4'hc)] : $signed(((7'h41) ?
                  reg1796 : reg1783)))));
          for (forvar1856 = (1'h0); (forvar1856 < (1'h1)); forvar1856 = (forvar1856 + (1'h1)))
            begin
              reg1857 <= reg1803;
              reg1858 <= (~^(reg1846 ?
                  (~$unsigned((reg1790 ?
                      reg1818 : reg1825))) : $unsigned(reg1797)));
            end
          for (forvar1859 = (1'h0); (forvar1859 < (3'h4)); forvar1859 = (forvar1859 + (1'h1)))
            begin
              reg1860 <= $unsigned((&$unsigned(($unsigned(reg1843) <<< reg1769))));
              reg1861 <= {(8'h9f),
                  ($signed($signed($unsigned(reg1833))) ?
                      (^~(!((7'h4e) ?
                          reg1822 : reg1833))) : reg1816[(5'h16):(4'hf)]),
                  $signed({(^$signed(reg1771)),
                      $unsigned({reg1843, reg1836, wire1764})})};
              reg1862 = (~^((((7'h58) > {reg1768, reg1769, reg1814}) ?
                  $unsigned((wire1760 | reg1800)) : $signed((^reg1858))) & (reg1768[(2'h2):(1'h0)] ?
                  $signed(reg1800) : ($unsigned(wire1763) <<< (!reg1843)))));
            end
        end
      else
        begin
          for (forvar1853 = (1'h0); (forvar1853 < (3'h6)); forvar1853 = (forvar1853 + (1'h1)))
            begin
              reg1854 = reg1803;
              reg1855 <= reg1829[(5'h14):(3'h7)];
              reg1856 = (~(reg1858 ?
                  (&reg1832[(2'h2):(1'h1)]) : (({reg1790, reg1768} >= reg1846) ?
                      (~&$signed(forvar1856)) : ($unsigned(forvar1853) ?
                          {reg1768} : reg1774))));
              reg1857 <= $signed($unsigned(({reg1856[(5'h10):(2'h2)]} ?
                  reg1828 : reg1826)));
            end
          if ($signed(($unsigned((^$unsigned(reg1856))) * ($signed(((8'hbe) ?
              reg1785 : reg1794)) & ((forvar1859 ?
              reg1775 : reg1816) < reg1828[(3'h6):(3'h4)])))))
            begin
              reg1858 <= $signed((~&(+((reg1858 ? reg1847 : reg1854) ?
                  $signed(reg1826) : $unsigned((7'h50))))));
              reg1859 = reg1799;
              reg1862 = (~^$unsigned(reg1833));
            end
          else
            begin
              reg1859 = $signed(reg1771);
              reg1862 = reg1769;
              reg1863 = reg1861[(3'h5):(1'h0)];
            end
          reg1864 <= ({(reg1846[(4'hf):(1'h1)] < (((7'h41) ?
                  reg1860 : reg1803) & $unsigned(reg1829))),
              (~|({wire1761, reg1857, reg1848} ?
                  (wire1762 > reg1818) : (|reg1853))),
              forvar1856} | reg1832[(2'h2):(2'h2)]);
          if ((-((reg1828 ?
              $signed((7'h58)) : reg1788[(4'hb):(1'h0)]) ^~ $signed((8'haa)))))
            begin
              reg1865 = reg1816[(1'h0):(1'h0)];
              reg1866 = $signed(($signed($signed($unsigned(reg1858))) >= reg1797[(4'h8):(3'h4)]));
              reg1867 = reg1826;
              reg1868 <= $unsigned($unsigned({reg1818[(3'h6):(2'h2)]}));
              reg1869 <= $signed(($signed($signed((|reg1818))) <<< (+reg1826)));
              reg1870 = ((((^~reg1771) | reg1853[(2'h2):(1'h1)]) & $signed($unsigned($signed(forvar1856)))) ?
                  (({reg1858[(2'h2):(1'h0)]} ?
                      reg1866 : ((-(8'hb7)) < reg1804)) || $unsigned({(reg1848 ?
                          reg1775 : reg1828)})) : (&$signed($unsigned($signed(reg1829)))));
            end
          else
            begin
              reg1868 <= reg1855[(3'h7):(3'h5)];
              reg1870 = (reg1825 >= reg1816[(5'h16):(5'h14)]);
              reg1871 = (reg1840 | (7'h56));
              reg1872 = (({({reg1794,
                          (7'h49)} >>> reg1832[(1'h0):(1'h0)])} < reg1788[(5'h11):(2'h2)]) ?
                  (~^reg1836) : $signed(forvar1856[(5'h15):(4'hb)]));
              reg1873 = wire1764;
              reg1874 = $unsigned(reg1873);
              reg1875 <= $signed($unsigned(reg1840[(3'h4):(3'h4)]));
            end
          reg1876 = ($unsigned(reg1868) ? wire1763 : reg1875);
          reg1877 <= reg1788;
          reg1878 <= $signed($signed(wire1763));
        end
      if ($unsigned((($signed(reg1814) ?
          $unsigned(((8'hb0) ? reg1868 : wire1763)) : {$signed((7'h4f)),
              (reg1856 ? reg1806 : reg1816),
              reg1797[(4'hb):(2'h2)]}) << reg1861[(2'h3):(1'h1)])))
        begin
          reg1879 = (reg1836[(3'h5):(3'h4)] & reg1769);
          reg1880 <= $unsigned($unsigned((!($unsigned(reg1775) << reg1791))));
        end
      else
        begin
          reg1880 <= reg1863[(3'h6):(1'h1)];
          reg1881 = (reg1828 ~^ $signed((reg1855[(1'h0):(1'h0)] ?
              reg1826 : reg1806[(5'h15):(4'h9)])));
          reg1882 = $unsigned(reg1797);
          reg1883 <= ((8'hb6) ?
              reg1777[(5'h14):(1'h1)] : ($signed(((reg1863 ^ reg1857) ?
                      $unsigned(reg1833) : reg1808)) ?
                  {(-(reg1796 < reg1882))} : reg1785[(3'h5):(1'h1)]));
          if ($unsigned(reg1882[(4'h9):(2'h2)]))
            begin
              reg1884 <= ($signed(reg1825[(3'h7):(3'h7)]) ?
                  reg1875 : {(8'h9c),
                      (|(reg1822[(4'h9):(3'h4)] << $unsigned(reg1788)))});
              reg1885 <= (reg1855[(1'h0):(1'h0)] ?
                  (^(((reg1882 << (7'h41)) == $signed(reg1877)) ?
                      (reg1846[(4'ha):(3'h4)] ^~ {reg1848,
                          reg1878}) : reg1859)) : $unsigned({$unsigned(((8'hbe) | (8'hbf))),
                      reg1854[(4'h8):(2'h2)]}));
              reg1886 <= ($unsigned(reg1783) ?
                  $signed((|(-$unsigned(reg1852)))) : reg1800);
              reg1887 = ((~(^(reg1785[(2'h2):(2'h2)] & (~|reg1766)))) ?
                  ((-($unsigned(reg1799) ? {reg1775} : $signed((8'hb6)))) ?
                      reg1832[(1'h1):(1'h0)] : reg1799) : ((~reg1856) >> $signed($signed($signed(reg1881)))));
              reg1888 = (8'hbe);
            end
          else
            begin
              reg1884 <= (~|$signed((8'hb5)));
              reg1885 <= ($signed((reg1867[(5'h11):(4'hb)] + reg1888[(3'h4):(2'h2)])) ?
                  (($signed((~|reg1838)) ?
                          (reg1848[(1'h0):(1'h0)] << (reg1864 ?
                              reg1832 : reg1804)) : reg1839) ?
                      {((wire1760 ? (7'h51) : reg1866) && $unsigned(reg1855)),
                          reg1825,
                          reg1847[(5'h1d):(3'h7)]} : ($signed((8'hbe)) ?
                          (^~reg1854[(5'h16):(2'h2)]) : (^wire1762[(1'h0):(1'h0)]))) : reg1854);
            end
          for (forvar1889 = (1'h0); (forvar1889 < (2'h3)); forvar1889 = (forvar1889 + (1'h1)))
            begin
              reg1890 = {((~|reg1768[(4'hb):(3'h4)]) ~^ reg1876[(2'h2):(2'h2)]),
                  {(reg1832 >>> $signed(((7'h45) && forvar1856))),
                      $unsigned($signed($unsigned(reg1799))),
                      $signed(((8'hba) ?
                          $signed(reg1814) : $unsigned(reg1847)))},
                  $unsigned(reg1766[(1'h1):(1'h0)])};
              reg1891 <= (!({reg1880[(5'h12):(1'h0)]} ?
                  ($unsigned($unsigned(reg1828)) ?
                      reg1890 : $unsigned(((7'h49) | reg1859))) : (reg1865 ?
                      $signed(wire1762[(4'h9):(3'h5)]) : $unsigned($unsigned(reg1890)))));
              reg1892 <= (|reg1882[(5'h14):(4'he)]);
              reg1893 <= $unsigned($signed(reg1796));
              reg1894 <= reg1876;
              reg1895 = $signed((reg1867 ? $signed(reg1870) : {reg1860}));
            end
        end
    end
  assign wire1896 = ($unsigned((((+reg1788) ?
                            (7'h56) : (-(8'haf))) & reg1843)) ?
                        (reg1824[(3'h5):(3'h4)] ?
                            reg1811[(4'h9):(3'h5)] : (8'hba)) : reg1804[(4'he):(1'h1)]);
  always
    @(posedge clk) begin
      reg1897 <= reg1864[(3'h4):(2'h3)];
      for (forvar1898 = (1'h0); (forvar1898 < (1'h0)); forvar1898 = (forvar1898 + (1'h1)))
        begin
          for (forvar1899 = (1'h0); (forvar1899 < (3'h5)); forvar1899 = (forvar1899 + (1'h1)))
            begin
              reg1900 <= $signed($unsigned(reg1858[(2'h3):(2'h3)]));
              reg1901 = ({({$unsigned(reg1785)} ?
                          reg1775[(1'h0):(1'h0)] : reg1883[(5'h17):(4'h9)])} ?
                  reg1885 : $unsigned(reg1775));
              reg1902 <= (8'hb9);
            end
          if ((~$signed(reg1828[(3'h4):(3'h4)])))
            begin
              reg1903 <= (7'h58);
              reg1904 <= ($unsigned($unsigned($signed((~^reg1838)))) ?
                  (($signed((&reg1861)) ?
                          {(reg1775 ? wire1760 : wire1763),
                              (reg1811 ?
                                  reg1868 : reg1788)} : ($signed(wire1762) ?
                              (reg1785 <= reg1838) : (reg1848 - reg1799))) ?
                      {($unsigned((7'h4f)) ?
                              (-reg1833) : (reg1826 ?
                                  (8'hb5) : reg1847))} : $signed((!{wire1760}))) : (($unsigned(reg1811) >= (~^(&(8'h9f)))) >= (~^reg1816[(3'h4):(2'h2)])));
              reg1905 <= $unsigned(reg1785[(1'h1):(1'h1)]);
              reg1906 <= {(({(reg1825 ? reg1864 : (7'h4e)),
                      ((8'ha0) ? wire1760 : wire1764),
                      (wire1765 ?
                          (8'hb2) : reg1891)} <= $unsigned(reg1847[(5'h14):(4'hb)])) >= $signed({(reg1791 | reg1832),
                      reg1785[(1'h1):(1'h1)],
                      reg1875})),
                  ($unsigned({{reg1783, forvar1898}, reg1891}) ?
                      $unsigned(reg1788) : reg1833[(2'h3):(1'h1)])};
            end
          else
            begin
              reg1907 = (~^reg1886);
              reg1908 <= $signed(reg1904[(1'h1):(1'h0)]);
              reg1909 = $unsigned($unsigned(($unsigned($unsigned(reg1883)) ?
                  $signed(wire1764[(4'hd):(4'h8)]) : reg1836)));
              reg1910 = ((({reg1811} & (reg1833 ?
                      reg1790 : $signed(reg1811))) - reg1907[(3'h5):(3'h4)]) ?
                  $signed($unsigned(reg1880)) : $unsigned(wire1760));
              reg1911 <= reg1819[(2'h2):(1'h0)];
              reg1912 <= reg1877;
            end
          for (forvar1913 = (1'h0); (forvar1913 < (1'h1)); forvar1913 = (forvar1913 + (1'h1)))
            begin
              reg1914 <= $signed((8'hba));
              reg1915 <= $unsigned((~^(~($signed(reg1910) >> reg1769[(4'he):(1'h1)]))));
              reg1916 = ($signed($signed($unsigned(((8'hb9) >>> (7'h56))))) <<< (&reg1893[(2'h2):(1'h0)]));
              reg1917 <= ((-$signed($unsigned(reg1816[(4'hd):(4'ha)]))) ?
                  reg1861[(4'h8):(1'h0)] : reg1897);
              reg1918 = $signed($unsigned(reg1900));
              reg1919 = ((reg1806[(5'h17):(5'h12)] < (reg1828 ?
                  ((reg1825 ?
                      reg1892 : reg1911) * $signed(reg1840)) : $unsigned($signed(wire1762)))) ^~ ($signed(wire1896) ?
                  ($signed((wire1760 ?
                      reg1843 : (8'hb2))) <<< (~^reg1900)) : (!{$unsigned(reg1826),
                      ((7'h56) ^~ reg1782)})));
            end
          reg1920 = ($unsigned(wire1761) == (-(reg1880 ^~ reg1894)));
          reg1921 = reg1771[(1'h0):(1'h0)];
          for (forvar1922 = (1'h0); (forvar1922 < (2'h3)); forvar1922 = (forvar1922 + (1'h1)))
            begin
              reg1923 <= ($signed((~reg1775)) ?
                  ((reg1836[(1'h0):(1'h0)] ?
                          ((reg1911 >>> reg1836) ^ (reg1855 ?
                              reg1775 : (8'ha9))) : (~&$unsigned(reg1918))) ?
                      (^~$unsigned($unsigned(forvar1922))) : ((|$signed(reg1826)) | (((8'h9f) ?
                              reg1811 : reg1785) ?
                          (reg1814 > reg1785) : reg1900))) : $signed(reg1900));
              reg1924 = $signed(wire1762);
              reg1925 = ($unsigned((!(reg1768 ?
                      (forvar1922 && reg1806) : reg1822))) ?
                  $unsigned(reg1816[(5'h11):(4'he)]) : reg1840[(3'h7):(1'h1)]);
            end
          reg1926 <= $unsigned($unsigned((($unsigned(reg1806) ?
                  (reg1914 + reg1796) : (reg1785 ? reg1769 : reg1811)) ?
              {(8'hbb),
                  (reg1864 ? reg1826 : reg1924),
                  (&wire1763)} : (wire1762[(4'hb):(1'h0)] ?
                  reg1794 : $signed(reg1846)))));
        end
      reg1927 = $unsigned({{((reg1796 ? (8'ha9) : reg1775) <= (reg1884 ?
                  reg1818 : (7'h4b)))},
          (reg1829 + $signed(((7'h57) > reg1910)))});
    end
  always
    @(posedge clk) begin
      if ((~&$unsigned(($signed(reg1875) ^ $signed($signed(reg1897))))))
        begin
          if ((|((((7'h4a) ^~ reg1868[(1'h0):(1'h0)]) - reg1864[(4'hc):(3'h6)]) << reg1768)))
            begin
              reg1928 <= $signed((($unsigned($unsigned(reg1790)) ?
                  $signed({reg1843}) : {reg1864,
                      (reg1897 ? reg1878 : wire1765),
                      (reg1838 >> reg1880)}) ^ reg1894[(4'hb):(1'h0)]));
              reg1929 = $signed((~^((-$unsigned(reg1915)) ?
                  reg1905[(2'h2):(1'h0)] : (~^(wire1761 & reg1819)))));
              reg1930 = (reg1897 + $unsigned(reg1838[(5'h13):(3'h6)]));
              reg1931 = (($unsigned(((reg1900 ? reg1928 : reg1825) == {reg1774,
                      wire1761,
                      reg1843})) ~^ (7'h4f)) ?
                  $unsigned($signed($signed($signed(reg1893)))) : $unsigned((|(^(-(7'h48))))));
            end
          else
            begin
              reg1928 <= (({reg1791[(1'h1):(1'h0)],
                          (~&reg1782[(5'h11):(4'h9)]),
                          ((reg1912 <<< reg1878) ?
                              ((8'h9e) ?
                                  reg1858 : reg1790) : ((8'hae) - reg1883))} ?
                      {(&(|reg1858))} : wire1763) ?
                  {(|((~|(8'ha7)) ?
                          $unsigned(reg1828) : reg1808[(4'hd):(3'h6)]))} : $signed(reg1884));
              reg1929 = reg1926[(4'h9):(3'h6)];
              reg1930 = ($unsigned((((wire1765 ?
                      reg1857 : reg1826) ^ $unsigned(reg1885)) ?
                  reg1897[(4'he):(2'h2)] : wire1760)) || $signed((~|(reg1774[(3'h4):(1'h0)] < reg1869))));
              reg1931 = ((8'ha0) ?
                  (7'h58) : {$unsigned($unsigned((reg1839 ?
                          reg1818 : wire1896))),
                      $unsigned(reg1774[(1'h0):(1'h0)])});
            end
          for (forvar1932 = (1'h0); (forvar1932 < (3'h5)); forvar1932 = (forvar1932 + (1'h1)))
            begin
              reg1933 <= $signed(reg1794);
              reg1934 = (8'ha6);
              reg1935 <= ((reg1788 <<< (~^{(reg1891 & reg1799),
                  reg1860[(2'h2):(1'h1)]})) | (reg1847[(5'h14):(4'h9)] ^ ((~&{reg1864,
                  reg1846}) ~^ (-{reg1864, reg1928, reg1788}))));
            end
          reg1936 <= $signed($unsigned((reg1838 ?
              $unsigned(reg1771[(2'h3):(1'h1)]) : reg1853)));
          for (forvar1937 = (1'h0); (forvar1937 < (3'h4)); forvar1937 = (forvar1937 + (1'h1)))
            begin
              reg1938 = reg1847;
              reg1939 = (|reg1846[(5'h14):(4'ha)]);
              reg1940 <= ((reg1788[(4'hf):(4'h9)] & reg1926[(3'h5):(3'h5)]) ^~ wire1765[(3'h4):(2'h2)]);
            end
          if (((^reg1930) ?
              $signed(((((8'ha1) ?
                  reg1906 : reg1926) && (reg1814 * reg1826)) <<< $signed($unsigned(reg1768)))) : (reg1774 || $signed(({reg1818,
                  (8'ha9)} + $unsigned(reg1769))))))
            begin
              reg1941 = $signed($signed(($signed(reg1883) ?
                  reg1775[(1'h1):(1'h1)] : (|reg1864[(3'h5):(1'h1)]))));
              reg1942 <= {(^~reg1788[(4'ha):(4'h8)]), reg1914};
              reg1943 <= (reg1905[(1'h0):(1'h0)] ?
                  (^~reg1840) : $signed($unsigned((((7'h58) * reg1768) ?
                      wire1763[(2'h3):(1'h0)] : (~|reg1839)))));
              reg1944 = {reg1935};
              reg1945 = (~^(^~(^(reg1838[(4'h8):(2'h2)] ?
                  reg1893[(3'h6):(1'h1)] : reg1902[(3'h5):(3'h5)]))));
            end
          else
            begin
              reg1941 = $signed(((~&(~&(reg1912 ?
                  reg1877 : reg1903))) == $unsigned({(reg1943 << reg1818),
                  (reg1800 & reg1832)})));
              reg1944 = ((8'ha5) * {(reg1883 ?
                      $unsigned((reg1822 ?
                          (7'h48) : reg1782)) : $unsigned($unsigned(reg1826))),
                  reg1928});
            end
        end
      else
        begin
          if ((reg1868[(2'h2):(2'h2)] <= $unsigned(reg1941)))
            begin
              reg1929 = wire1896;
              reg1932 <= ((({{(8'haf), reg1885, reg1797}, $unsigned(wire1760)} ?
                      ((8'hb0) + reg1806) : (|(~|reg1931))) <<< $unsigned($unsigned((8'had)))) ?
                  reg1885 : (($signed(reg1829[(4'hb):(2'h2)]) ?
                          (+(8'hbb)) : ($unsigned(reg1824) ?
                              $signed((8'hb3)) : reg1808)) ?
                      (($signed(reg1945) >> $signed(reg1847)) ?
                          $signed((reg1936 ?
                              reg1923 : reg1915)) : reg1824) : {reg1877,
                          ((~|reg1838) ?
                              (reg1940 || reg1769) : reg1806[(5'h18):(4'hd)]),
                          $signed({reg1864})}));
              reg1934 = ((|{((8'h9c) ~^ $signed(reg1797)),
                  (reg1915[(4'h8):(3'h5)] - (reg1860 ~^ reg1864)),
                  (reg1939 || $unsigned(reg1829))}) <= (8'hbd));
              reg1935 <= ({reg1839[(3'h5):(1'h1)], $unsigned(reg1878)} ?
                  $unsigned(reg1777) : $signed((7'h43)));
            end
          else
            begin
              reg1929 = reg1853;
              reg1932 <= $signed(($unsigned((reg1884 || {reg1848,
                  reg1928,
                  reg1796})) ^~ $signed($unsigned((reg1791 >>> reg1931)))));
              reg1934 = (!($signed((-(-reg1791))) ?
                  {(-reg1769),
                      reg1766,
                      wire1765} : (reg1908[(4'hb):(4'ha)] & (((8'ha6) ?
                      reg1769 : reg1797) <<< $unsigned((7'h41))))));
              reg1937 = (+(+({(reg1855 ? reg1877 : reg1942),
                      (reg1875 | reg1933),
                      reg1785} ?
                  reg1930 : ((7'h50) < reg1783[(4'ha):(3'h7)]))));
              reg1940 <= {reg1860[(4'ha):(3'h4)],
                  ((reg1847[(5'h15):(5'h12)] ?
                          $unsigned((reg1923 ?
                              reg1768 : reg1800)) : $unsigned(forvar1937)) ?
                      (({reg1935, wire1896} ?
                          reg1806[(4'h9):(1'h0)] : {reg1833,
                              wire1762}) >> $unsigned((reg1811 || wire1762))) : (7'h58))};
              reg1941 = (reg1768[(4'he):(1'h0)] > ((reg1904[(1'h1):(1'h0)] > (7'h4c)) ?
                  $unsigned(reg1894[(3'h7):(2'h2)]) : $unsigned(((^~(8'hb0)) && (|(7'h55))))));
              reg1942 <= $signed((~&(((reg1932 ?
                      reg1883 : reg1790) <<< (-reg1884)) ?
                  ((&reg1818) ?
                      (reg1774 ?
                          reg1904 : reg1848) : $signed(reg1904)) : $unsigned(reg1883))));
            end
          reg1944 = ((reg1806 + $unsigned(reg1791)) && (~&$unsigned(reg1797)));
          reg1945 = (reg1914 ?
              reg1796 : $unsigned((reg1892 | $signed(((8'hbe) ?
                  reg1785 : reg1897)))));
          reg1946 <= ({$signed($unsigned(reg1941)),
              ((+reg1804) ?
                  reg1885[(4'hd):(1'h0)] : ($signed(reg1860) ?
                      (reg1940 - (8'hbb)) : reg1794[(4'ha):(4'h8)])),
              (|$signed($signed(reg1885)))} ^ (reg1933 < $signed($signed(reg1880))));
          for (forvar1947 = (1'h0); (forvar1947 < (3'h4)); forvar1947 = (forvar1947 + (1'h1)))
            begin
              reg1948 <= (((~$unsigned((|reg1938))) << (reg1886 ?
                      reg1864[(4'hb):(3'h5)] : $unsigned(reg1884[(4'hb):(4'ha)]))) ?
                  reg1846[(1'h1):(1'h1)] : (~&reg1800[(4'hc):(3'h5)]));
              reg1949 = $unsigned(((-((reg1940 && reg1799) <= $signed(reg1868))) ?
                  $unsigned(reg1903) : $unsigned($unsigned((&(8'h9d))))));
              reg1950 <= (+((^~$unsigned($unsigned(reg1937))) ?
                  ((8'ha0) ?
                      $unsigned(((7'h42) ?
                          reg1839 : reg1825)) : {(reg1869 * (7'h53)),
                          (reg1948 ? reg1936 : (8'h9f)),
                          $unsigned(reg1940)}) : (($signed(reg1769) ?
                          (wire1762 ? forvar1947 : reg1936) : ((8'hb4) ?
                              reg1800 : reg1926)) ?
                      $signed((reg1948 & (7'h52))) : {{reg1788,
                              reg1799,
                              (8'ha0)}})));
            end
        end
      if (((wire1760 < (~|$unsigned(((7'h4f) ? reg1828 : (8'hb7))))) ?
          (!reg1836) : reg1799[(4'ha):(3'h7)]))
        begin
          for (forvar1951 = (1'h0); (forvar1951 < (1'h0)); forvar1951 = (forvar1951 + (1'h1)))
            begin
              reg1952 = {reg1838};
              reg1953 = {reg1936[(4'hc):(1'h0)], reg1931, reg1886};
              reg1954 <= ((8'ha2) ^ reg1839[(1'h1):(1'h0)]);
              reg1955 = (((+(&{reg1824,
                      forvar1932})) && (~reg1875[(3'h6):(3'h6)])) ?
                  reg1860[(2'h3):(2'h3)] : ($signed(((reg1832 ?
                          (7'h54) : reg1825) != (reg1884 ?
                          reg1832 : reg1948))) ?
                      (reg1803 ?
                          reg1796[(2'h3):(1'h1)] : ((reg1900 >>> reg1785) * {reg1943})) : ((~^$signed(reg1939)) > $signed(((7'h47) >>> reg1818)))));
              reg1956 <= reg1824[(4'h9):(2'h3)];
              reg1957 = reg1877;
              reg1958 = (({$signed($signed((8'hb8))),
                          reg1828[(5'h15):(1'h1)],
                          $unsigned($signed(reg1942))} ?
                      $unsigned(wire1760[(4'ha):(1'h1)]) : $signed((^$unsigned((8'hb9))))) ?
                  (((~|(forvar1932 ? reg1948 : reg1848)) ?
                      {reg1833, $unsigned((7'h55)), (|reg1775)} : ((8'h9f) ?
                          $signed(reg1932) : $unsigned(reg1853))) & reg1860) : reg1833);
            end
          reg1959 = $signed($signed($signed(reg1953[(4'h8):(2'h2)])));
          reg1960 = $unsigned(($unsigned({(reg1825 >> reg1948),
              $signed(reg1958)}) * (~&reg1934)));
          if (reg1797[(1'h0):(1'h0)])
            begin
              reg1961 <= (reg1904[(1'h0):(1'h0)] - $signed($unsigned((-$unsigned(reg1839)))));
              reg1962 <= reg1771[(1'h1):(1'h0)];
            end
          else
            begin
              reg1961 <= ((^({(~&reg1884),
                  (reg1788 == reg1768),
                  $unsigned(wire1760)} * reg1949)) != ({(^reg1912)} >> reg1935));
              reg1962 <= $signed(($unsigned($signed((reg1858 ?
                      reg1930 : reg1819))) ?
                  reg1822 : $signed((reg1932[(4'ha):(3'h6)] ?
                      (reg1940 ? reg1869 : (7'h57)) : $signed(reg1869)))));
            end
        end
      else
        begin
          for (forvar1951 = (1'h0); (forvar1951 < (3'h6)); forvar1951 = (forvar1951 + (1'h1)))
            begin
              reg1954 <= reg1766[(3'h6):(2'h2)];
              reg1955 = $unsigned((reg1791[(1'h0):(1'h0)] ?
                  $signed((~^reg1939)) : ($signed($signed((8'ha3))) ?
                      reg1957[(3'h4):(1'h1)] : $unsigned((^(7'h53))))));
              reg1957 = ((+((~^(~|reg1893)) - $signed((reg1930 >>> reg1777)))) && ($unsigned($signed((reg1788 ?
                  reg1908 : reg1911))) == (((-reg1960) < (!reg1935)) ?
                  $signed((reg1840 ?
                      reg1944 : reg1894)) : reg1838[(1'h1):(1'h0)])));
              reg1961 <= (($signed(reg1836[(1'h1):(1'h1)]) >= (~&((-reg1846) ?
                      (!(7'h41)) : (|reg1930)))) ?
                  $signed(reg1937[(3'h7):(2'h2)]) : (^~$signed($signed($signed((7'h47))))));
              reg1963 = reg1912[(1'h0):(1'h0)];
              reg1964 = $signed(reg1828);
            end
          for (forvar1965 = (1'h0); (forvar1965 < (1'h1)); forvar1965 = (forvar1965 + (1'h1)))
            begin
              reg1966 <= (reg1868[(1'h0):(1'h0)] + (~(reg1961[(3'h5):(3'h4)] ?
                  (~^reg1822) : (~&(reg1961 << reg1883)))));
            end
          reg1967 <= $unsigned(reg1875[(1'h0):(1'h0)]);
          for (forvar1968 = (1'h0); (forvar1968 < (3'h6)); forvar1968 = (forvar1968 + (1'h1)))
            begin
              reg1969 = reg1905[(2'h3):(2'h2)];
              reg1970 = (reg1788[(5'h17):(3'h4)] == (wire1763 ?
                  ((^~reg1800) ^ $signed((reg1911 | reg1822))) : ($signed(reg1905[(1'h1):(1'h1)]) ?
                      $unsigned((^reg1926)) : reg1936)));
              reg1971 = reg1937;
            end
          if (($signed($signed(reg1880)) ? reg1769 : reg1957[(4'ha):(3'h5)]))
            begin
              reg1972 = (|(~(~&($signed(reg1836) ?
                  $signed(reg1934) : reg1932))));
              reg1973 <= reg1958[(4'he):(4'hb)];
              reg1974 = $unsigned({(~^(~|$unsigned(reg1791)))});
              reg1975 = ($signed((!($unsigned(reg1948) ?
                  reg1796 : (reg1846 ? (8'hb0) : (8'ha2))))) <<< (8'hb4));
              reg1976 = (((~((reg1832 ?
                      reg1840 : reg1912) ^ reg1948)) ~^ (($signed(reg1966) ?
                      reg1877[(2'h3):(1'h0)] : (~reg1952)) ^ reg1803)) ?
                  {$unsigned((^(7'h49))),
                      reg1803[(1'h0):(1'h0)],
                      ($signed((reg1958 ?
                          reg1963 : reg1914)) << $unsigned(reg1833[(5'h11):(2'h3)]))} : (reg1950[(4'hd):(3'h6)] ?
                      ((~|(|reg1917)) ^~ (((8'ha7) ?
                          (8'hb6) : reg1822) * $unsigned(reg1829))) : $unsigned($unsigned((reg1891 ?
                          reg1936 : (7'h51))))));
              reg1977 <= (($signed(reg1769) + $unsigned(($unsigned(wire1763) ^~ $signed(reg1884)))) ?
                  ($signed(($signed(wire1762) ?
                      wire1765[(3'h4):(2'h3)] : {reg1797,
                          reg1972,
                          reg1972})) + (((~|reg1894) ?
                      (reg1933 ?
                          reg1843 : reg1911) : $signed((7'h53))) > $signed((forvar1951 ^ (8'ha4))))) : (-reg1976));
              reg1978 <= reg1860;
            end
          else
            begin
              reg1972 = ($unsigned(((~&reg1790[(2'h3):(1'h1)]) | reg1937)) ?
                  reg1855 : (~|($unsigned((^~reg1894)) >>> $signed(reg1782[(4'hf):(4'h9)]))));
              reg1974 = reg1953[(2'h3):(2'h3)];
              reg1975 = $signed(((({reg1883, reg1900} ?
                          $unsigned(reg1836) : (~&reg1822)) ?
                      {(reg1926 >= reg1814)} : $signed({reg1948})) ?
                  $signed((~|(!(8'ha1)))) : reg1858));
              reg1977 <= reg1944;
              reg1978 <= $unsigned($unsigned((!$signed({wire1896}))));
              reg1979 <= ((((&(reg1945 & reg1846)) ?
                          ({reg1956,
                              reg1794,
                              reg1893} >= (reg1788 < reg1875)) : reg1843) ?
                      $signed((reg1777[(3'h5):(2'h2)] ?
                          (reg1816 ?
                              reg1944 : reg1957) : $unsigned(reg1955))) : $signed((|(reg1955 ^~ reg1946)))) ?
                  (reg1961 >> (|$signed($unsigned(forvar1947)))) : ((~|(|(reg1864 && reg1797))) >> reg1864[(4'h9):(4'h9)]));
              reg1980 = (((-reg1962[(4'he):(4'hc)]) < reg1829[(1'h0):(1'h0)]) ?
                  reg1969[(1'h1):(1'h0)] : (7'h57));
            end
          reg1981 <= (reg1973[(3'h7):(1'h1)] <= $unsigned(reg1904[(1'h0):(1'h0)]));
          reg1982 <= ((&(reg1950 ?
              (-(reg1962 ? reg1902 : reg1976)) : {reg1943[(1'h0):(1'h0)],
                  reg1875,
                  (~|reg1804)})) * (reg1944[(1'h1):(1'h1)] ?
              $unsigned(wire1761) : reg1864[(4'hb):(2'h3)]));
        end
      for (forvar1983 = (1'h0); (forvar1983 < (3'h5)); forvar1983 = (forvar1983 + (1'h1)))
        begin
          for (forvar1984 = (1'h0); (forvar1984 < (2'h3)); forvar1984 = (forvar1984 + (1'h1)))
            begin
              reg1985 <= reg1884[(5'h10):(1'h1)];
              reg1986 = reg1858;
              reg1987 <= $signed(($signed($unsigned($unsigned((8'ha5)))) & (~&(reg1783[(2'h3):(1'h1)] >>> (&reg1964)))));
            end
          reg1988 = (((8'had) > {reg1808,
              $signed((~^reg1803)),
              (8'ha7)}) | (7'h47));
        end
      reg1989 = (({$unsigned($signed(wire1762)),
              (reg1975 ~^ $signed(reg1906)),
              (reg1945 >>> reg1847[(3'h7):(3'h5)])} < {reg1848,
              $signed((reg1986 < reg1864))}) ?
          $signed($unsigned(reg1893[(3'h5):(2'h3)])) : (reg1946[(5'h18):(4'hf)] ?
              {reg1832} : $signed(reg1796)));
    end
  always
    @(posedge clk) begin
      reg1990 <= $unsigned(({reg1774[(1'h0):(1'h0)]} ^ (-($signed(reg1926) ?
          (8'hb4) : $signed(reg1942)))));
      reg1991 <= (($unsigned(reg1908) | $unsigned(reg1981[(5'h10):(3'h4)])) ?
          $signed($signed($signed($signed(reg1928)))) : $signed(reg1926[(4'hc):(4'ha)]));
      reg1992 = {(~&($signed($signed(reg1803)) ?
              $unsigned((8'ha5)) : (+(wire1765 != reg1839))))};
      reg1993 <= ($unsigned((((~wire1764) < (wire1763 ~^ reg1917)) + reg1935[(3'h4):(1'h1)])) ?
          $unsigned($signed($signed($signed(reg1771)))) : {(8'hb6),
              $unsigned(reg1973[(5'h12):(2'h3)])});
      reg1994 = $unsigned((({(^~(8'hb5)),
          reg1914[(4'hc):(4'ha)],
          reg1804[(4'hb):(1'h1)]} > reg1894[(2'h2):(1'h1)]) >> (~&$signed($signed(reg1808)))));
      if (reg1788)
        begin
          if (reg1808)
            begin
              reg1995 <= $unsigned((^~reg1799[(5'h14):(2'h3)]));
              reg1996 = reg1967[(2'h2):(2'h2)];
              reg1997 = $signed({reg1981,
                  $signed($signed(((7'h52) ? reg1868 : reg1990)))});
              reg1998 <= $signed((^(|((~|reg1900) ?
                  $unsigned(reg1860) : reg1833[(4'hd):(4'h9)]))));
              reg1999 <= $unsigned(reg1908[(3'h7):(1'h1)]);
              reg2000 <= (~($signed((&$signed((8'haa)))) ?
                  ($unsigned((reg1777 ? wire1761 : reg1819)) ?
                      reg1912[(4'h8):(3'h7)] : (|reg1858[(3'h4):(1'h1)])) : (8'ha6)));
            end
          else
            begin
              reg1996 = (reg1932 >= ($signed(reg1993[(1'h1):(1'h0)]) ?
                  $unsigned((((8'h9f) ?
                      reg1973 : reg1883) ~^ reg1967)) : reg1946[(4'ha):(2'h3)]));
            end
          if (reg1816[(4'hf):(4'hb)])
            begin
              reg2001 <= (8'hb4);
              reg2002 <= ((reg1894 ?
                      ($unsigned($unsigned(reg1769)) ~^ $unsigned($signed((7'h4c)))) : $unsigned($unsigned($unsigned(reg1853)))) ?
                  (reg1979[(2'h3):(2'h2)] ?
                      reg1825[(4'hd):(4'hc)] : (reg1999[(4'hd):(4'h9)] && (reg1811 ^~ $signed(reg1996)))) : ((~&(~((8'hb8) & reg1824))) << $unsigned(reg1769)));
              reg2003 = $unsigned((+(-reg1782)));
            end
          else
            begin
              reg2003 = ($unsigned(reg1904) ?
                  (((8'hb8) >>> $unsigned((~|reg1868))) ^ reg1794) : reg1942[(5'h13):(4'h9)]);
            end
          reg2004 <= $signed((($unsigned((!(8'h9d))) ^ ((reg1868 ?
                  reg1903 : reg1785) || reg1904)) ?
              $signed(((reg1996 >>> reg1973) ?
                  reg1816 : reg1790[(3'h4):(2'h2)])) : $unsigned($unsigned($signed(reg1816)))));
          for (forvar2005 = (1'h0); (forvar2005 < (1'h0)); forvar2005 = (forvar2005 + (1'h1)))
            begin
              reg2006 <= (-(~(^(-(+reg1868)))));
              reg2007 <= $unsigned({{{{reg1803}}},
                  {$unsigned((reg1956 >= reg1926)),
                      $unsigned({(8'ha3)}),
                      (reg1982 & (reg1774 ? reg1993 : reg1886))},
                  reg1961});
              reg2008 = ((~&reg1914[(5'h11):(4'hb)]) << {reg1864});
            end
          reg2009 <= $unsigned((~&$signed(reg1880)));
          for (forvar2010 = (1'h0); (forvar2010 < (2'h2)); forvar2010 = (forvar2010 + (1'h1)))
            begin
              reg2011 = (($unsigned(reg1857[(3'h5):(2'h3)]) ?
                  ($signed((reg1822 ? reg1883 : (8'h9f))) ?
                      ($signed(reg1991) * reg1828[(1'h0):(1'h0)]) : ((8'hb0) && (reg1885 - reg1843))) : $unsigned((7'h40))) == $signed((^((reg1912 >> (8'ha4)) ?
                  (wire1896 ~^ reg1774) : reg1877))));
              reg2012 = {((&$signed($unsigned(reg1908))) != reg1868[(1'h1):(1'h0)]),
                  (~^({{(8'had)}, (reg1788 < reg1950), reg1766[(1'h1):(1'h0)]} ?
                      (reg1808[(1'h1):(1'h1)] ?
                          reg1911[(4'hc):(4'h9)] : reg1855) : reg1791[(1'h1):(1'h0)])),
                  $unsigned($unsigned({wire1896}))};
              reg2013 = (reg1775 >>> reg1825[(5'h15):(1'h1)]);
              reg2014 <= ($signed(reg1886) >= reg1878);
              reg2015 <= $unsigned({($signed(reg1829) != $unsigned((8'hba)))});
              reg2016 <= reg1838;
              reg2017 <= (($signed(((reg1897 - reg1991) >> (reg1928 >= reg1894))) ?
                      ((+(reg1860 ? reg1822 : reg1992)) ?
                          {$signed(reg1804),
                              (reg2000 ? reg1993 : reg1884),
                              reg1991[(1'h0):(1'h0)]} : $signed((reg1840 * (8'haa)))) : reg1803) ?
                  (reg1839 == (7'h4b)) : reg1804);
            end
          reg2018 <= $signed($unsigned(({reg2006, (~reg1967), {reg1782}} ?
              ({reg1814, reg1843, reg1883} ?
                  $unsigned(reg1891) : $unsigned((8'h9c))) : $unsigned(reg1855))));
        end
      else
        begin
          reg1995 <= ($unsigned((^~reg1987[(1'h0):(1'h0)])) + (7'h45));
          if ({$unsigned({(~^$unsigned(reg1914)),
                  $signed((reg1799 ? reg1768 : reg2017))}),
              $signed($unsigned((+{reg1981, reg1985, (7'h50)})))})
            begin
              reg1998 <= reg1877;
              reg2003 = $unsigned((((reg1808 * (reg1917 - wire1765)) & (&{reg1839,
                      reg1923})) ?
                  $signed((reg1928[(4'h9):(2'h3)] ?
                      $unsigned(reg1808) : reg1869)) : $unsigned({reg1839[(4'hd):(3'h7)],
                      $signed((8'hbc))})));
              reg2005 = $unsigned({$unsigned($signed((^~wire1763))),
                  ($signed((+reg1796)) != (~&$unsigned(reg1857))),
                  (+($signed(reg1846) ?
                      $unsigned((7'h44)) : $unsigned(reg1981)))});
              reg2008 = $unsigned(reg1998);
            end
          else
            begin
              reg1996 = $unsigned((!reg1891));
              reg1998 <= {reg2012};
              reg2003 = ({reg1857,
                  reg1777[(1'h1):(1'h1)],
                  wire1764[(4'hf):(4'ha)]} * (8'ha3));
              reg2004 <= reg1893[(3'h7):(1'h0)];
            end
          if ((({(-reg1962[(1'h0):(1'h0)]),
                  ($unsigned(wire1761) <= (reg1946 ? reg1839 : reg2000))} ?
              ($signed(reg1940) >> $unsigned({reg1962,
                  reg1915})) : (({reg2015} || (reg1928 ?
                  reg1836 : (8'h9d))) - (reg1846 ?
                  (reg1878 < reg1878) : reg1797))) < $signed(reg1897)))
            begin
              reg2009 <= (((~($signed((7'h50)) ?
                  {reg2011} : $signed(reg1923))) << (+(~(!reg1811)))) != reg1868[(1'h1):(1'h0)]);
            end
          else
            begin
              reg2009 <= ($unsigned(reg1915[(3'h6):(3'h4)]) ~^ reg1908[(1'h1):(1'h1)]);
              reg2010 <= {{($unsigned($signed(wire1765)) <<< ({reg1878} ?
                          (^~reg1897) : $unsigned(reg1892))),
                      (|(&reg1935))}};
            end
          reg2014 <= {(reg2011[(1'h0):(1'h0)] >= {((+reg1803) & $signed(reg1900)),
                  reg1858[(3'h6):(2'h3)]})};
          for (forvar2015 = (1'h0); (forvar2015 < (2'h3)); forvar2015 = (forvar2015 + (1'h1)))
            begin
              reg2016 <= reg2004;
              reg2019 = (+((^~(~^$unsigned(reg1933))) <<< $unsigned($signed((^forvar2015)))));
              reg2020 <= (($signed(($signed(reg1785) ?
                      {reg1956, reg1875} : (^~reg1993))) ?
                  $signed((-(reg1771 && reg1999))) : reg1777) & $signed((($signed(reg1883) ?
                  ((7'h56) || reg2004) : reg1864) || reg1788[(3'h7):(3'h7)])));
              reg2021 <= (!$unsigned(reg1811));
              reg2022 = $signed($unsigned((+reg1911)));
              reg2023 <= reg1840;
            end
          if ((^reg1777))
            begin
              reg2024 = {$unsigned((~|$unsigned($unsigned(reg1950)))),
                  $unsigned((reg1967[(4'hd):(3'h5)] > {$signed(reg2012),
                      (reg1803 + reg1905),
                      {(8'ha9), reg1884}})),
                  (~|reg2023[(4'he):(3'h4)])};
              reg2025 = (!($signed($signed($unsigned((7'h4f)))) ^ (forvar2005[(5'h10):(5'h10)] >= reg1880)));
              reg2026 = reg1836[(1'h0):(1'h0)];
            end
          else
            begin
              reg2024 = (~^(&(|$signed((8'hb1)))));
              reg2027 <= reg2017;
              reg2028 <= (~^reg2005[(3'h6):(3'h4)]);
              reg2029 <= ($unsigned($unsigned(reg2002[(1'h0):(1'h0)])) ?
                  (&((~&reg1928[(4'hd):(3'h4)]) ?
                      ($unsigned(reg1800) ?
                          (^~(8'ha9)) : (reg1875 ?
                              (7'h48) : reg1928)) : reg1804)) : (~&$signed($unsigned($unsigned((8'h9e))))));
              reg2030 <= ({reg2023} ?
                  (^~$signed({reg1824})) : $signed((^~$unsigned(((8'h9f) < reg1891)))));
            end
          reg2031 = $unsigned(reg2000[(4'ha):(4'ha)]);
        end
      for (forvar2032 = (1'h0); (forvar2032 < (1'h1)); forvar2032 = (forvar2032 + (1'h1)))
        begin
          if (reg2030)
            begin
              reg2033 = $unsigned($signed((($signed(reg1819) == (reg2004 ?
                      reg2019 : reg1997)) ?
                  $unsigned((reg1811 && forvar2010)) : (reg1999[(4'ha):(2'h3)] | reg1818[(3'h6):(3'h5)]))));
            end
          else
            begin
              reg2033 = $unsigned(($unsigned({$unsigned(reg1973),
                      ((8'ha0) ? reg1946 : reg1935),
                      (^reg1905)}) ?
                  {$unsigned((reg1886 ? reg1800 : reg1936))} : reg2028));
            end
          reg2034 = ($unsigned((~reg1993[(3'h4):(3'h4)])) ?
              ({(8'ha7)} >= reg2018[(4'h8):(1'h0)]) : ({reg1987} ?
                  ($unsigned((reg1997 ? (8'hb5) : (7'h40))) + {(reg1878 ?
                          reg1928 : reg1868)}) : ($unsigned(reg1791[(1'h1):(1'h1)]) >> $signed(reg2003[(1'h0):(1'h0)]))));
          for (forvar2035 = (1'h0); (forvar2035 < (2'h2)); forvar2035 = (forvar2035 + (1'h1)))
            begin
              reg2036 = (+$signed((reg1978[(3'h4):(2'h2)] - $signed($unsigned(reg1911)))));
              reg2037 <= forvar2015[(5'h18):(4'hf)];
              reg2038 <= reg2028;
              reg2039 <= reg1935[(2'h3):(1'h0)];
              reg2040 = (-reg2033[(3'h5):(1'h0)]);
              reg2041 = (reg1978 ? $unsigned((7'h55)) : reg1932[(3'h7):(1'h0)]);
            end
          reg2042 <= (|(~|(((~^reg1923) ~^ reg2011) ?
              (~&$unsigned(reg1855)) : reg1806)));
        end
    end
  assign wire2043 = ($signed({wire1760[(5'h10):(4'h9)],
                            ((reg1885 ? wire1761 : reg1797) ?
                                {reg1768, reg1933} : ((7'h4d) ^~ reg1855)),
                            reg1824[(4'h8):(3'h5)]}) ?
                        $signed((7'h46)) : reg2020);
  always
    @(posedge clk) begin
      for (forvar2044 = (1'h0); (forvar2044 < (1'h1)); forvar2044 = (forvar2044 + (1'h1)))
        begin
          if ((~&$signed($signed(reg1861[(4'h8):(1'h1)]))))
            begin
              reg2045 = $unsigned(reg1832);
              reg2046 <= ((~$signed((((8'h9e) >>> reg1788) >= $signed(reg1822)))) ?
                  {reg1777} : {$signed(((reg1993 ?
                          reg1940 : reg2028) == reg1933[(3'h4):(3'h4)]))});
              reg2047 <= $unsigned(reg1775[(3'h5):(1'h0)]);
              reg2048 <= $unsigned($signed($signed($unsigned((^reg1999)))));
            end
          else
            begin
              reg2045 = $signed(reg2014);
            end
        end
      reg2049 <= reg1794[(4'hc):(3'h4)];
      reg2050 = (wire1896 ?
          ($unsigned(((8'ha7) && (reg1768 ?
              reg1869 : reg1803))) << $unsigned(reg2028[(5'h10):(3'h7)])) : (((~^(7'h58)) > (reg1785[(2'h2):(2'h2)] ?
                  reg2048 : reg1904[(3'h5):(2'h2)])) ?
              ($signed((reg1846 != reg1799)) >>> $signed((-reg1935))) : $unsigned(reg1877[(1'h0):(1'h0)])));
      for (forvar2051 = (1'h0); (forvar2051 < (1'h0)); forvar2051 = (forvar2051 + (1'h1)))
        begin
          if ($unsigned((!((|{reg1855, reg1956, reg1855}) ?
              ((~^(7'h4a)) | (~|reg1799)) : (forvar2051[(4'h8):(2'h3)] ?
                  reg2015 : {reg1923, (7'h4b), reg1818})))))
            begin
              reg2052 <= $unsigned($signed((|reg1794[(2'h2):(1'h1)])));
              reg2053 <= ($signed(reg1769[(4'hc):(2'h2)]) <= (reg1999 <= reg1774));
              reg2054 <= reg1893;
              reg2055 = $unsigned(reg1962[(3'h6):(2'h2)]);
            end
          else
            begin
              reg2052 <= ((|($signed(reg2048[(3'h5):(3'h4)]) + $unsigned((~reg2006)))) ?
                  reg1774 : wire1762[(3'h5):(2'h3)]);
              reg2053 <= reg1777;
              reg2054 <= $unsigned(($signed(reg2007) | $signed(reg1875)));
              reg2056 <= (^reg1783[(3'h4):(3'h4)]);
            end
          reg2057 <= ({{$unsigned((+reg1900)), (7'h51)},
              (7'h46),
              (reg1966 <<< (reg2039[(3'h7):(2'h2)] < $unsigned(reg1838)))} <<< (+{$signed((reg1933 ?
                  (8'hb4) : reg1991))}));
          for (forvar2058 = (1'h0); (forvar2058 < (3'h5)); forvar2058 = (forvar2058 + (1'h1)))
            begin
              reg2059 = reg1880;
              reg2060 <= ($unsigned((7'h42)) ?
                  $signed(($unsigned((reg2020 << reg2016)) ?
                      (reg2037 >= (reg2030 ?
                          reg1940 : reg1923)) : $unsigned((reg1915 ?
                          reg1848 : (8'had))))) : $signed($signed(reg2010[(4'h9):(3'h5)])));
              reg2061 = $unsigned(reg2052);
              reg2062 <= reg2004[(4'hd):(1'h1)];
              reg2063 <= $unsigned((~|($signed($signed(reg1878)) ?
                  $signed(reg1877) : ((~&reg2015) ?
                      $unsigned(reg1904) : reg1880))));
            end
          reg2064 <= $signed($unsigned(wire1761));
          reg2065 <= (7'h46);
        end
      reg2066 <= (-(^~reg1961[(1'h1):(1'h1)]));
      reg2067 <= $unsigned($unsigned(reg1904[(3'h4):(2'h2)]));
    end
  always
    @(posedge clk) begin
      if (reg1775)
        begin
          reg2068 = $signed((($signed($unsigned(reg1796)) ?
              $unsigned(reg1891[(2'h2):(1'h1)]) : (^~$unsigned(reg1853))) > reg1981[(4'hf):(3'h5)]));
          reg2069 = ((-reg1869) ?
              reg2014[(4'hb):(3'h4)] : $unsigned($unsigned($unsigned((reg1869 ?
                  (7'h58) : reg1783)))));
        end
      else
        begin
          reg2068 = $unsigned({(8'haa)});
          reg2070 <= $unsigned(((reg1923 & $unsigned(((8'ha0) ?
              (8'hb3) : reg1883))) << reg1791[(2'h2):(1'h1)]));
          reg2071 <= reg1832[(1'h1):(1'h1)];
        end
      if ((reg2052 ?
          reg1768[(4'ha):(4'ha)] : ($unsigned($signed((reg2010 <<< reg1804))) ?
              (~$unsigned($signed(reg1956))) : reg2038[(4'h8):(2'h3)])))
        begin
          for (forvar2072 = (1'h0); (forvar2072 < (3'h6)); forvar2072 = (forvar2072 + (1'h1)))
            begin
              reg2073 <= $unsigned({$signed($signed((-reg1923)))});
              reg2074 = (^($signed((|$signed(reg1940))) ~^ $signed($signed(reg2015[(4'h9):(3'h7)]))));
            end
          for (forvar2075 = (1'h0); (forvar2075 < (3'h5)); forvar2075 = (forvar2075 + (1'h1)))
            begin
              reg2076 = ($signed(reg1902) ?
                  $unsigned($unsigned(reg1814[(3'h4):(2'h3)])) : {(!$unsigned({reg1985,
                          reg1808}))});
            end
          if ((((($signed(reg1923) ? (~wire1762) : $signed(wire1896)) ?
                      (!(7'h47)) : (-{reg1846})) ?
                  reg2015[(3'h7):(1'h1)] : (8'hb7)) ?
              ($signed((~&$signed(reg1956))) ?
                  (~&((^~reg2056) <<< reg1769)) : $signed(((~^reg1897) << reg1861[(1'h0):(1'h0)]))) : reg1875))
            begin
              reg2077 = $unsigned((((-(reg1942 >= reg2064)) ?
                  reg1804 : $signed((reg1847 ?
                      reg1829 : reg1840))) == reg1950[(5'h19):(4'h8)]));
              reg2078 <= $unsigned(reg2018[(1'h0):(1'h0)]);
              reg2079 = (reg2002[(2'h3):(1'h1)] ?
                  ($unsigned((^~(reg2030 <<< forvar2072))) ?
                      $unsigned(reg2066[(1'h1):(1'h1)]) : $signed((7'h53))) : (!reg1782[(2'h3):(2'h3)]));
              reg2080 = reg1936[(1'h0):(1'h0)];
              reg2081 = $unsigned($signed($signed($signed((reg2079 >= reg1932)))));
            end
          else
            begin
              reg2077 = $unsigned(((8'haa) ?
                  reg1777 : ($unsigned((reg1884 ? reg1878 : reg2010)) ?
                      (7'h54) : reg1904[(3'h5):(2'h3)])));
            end
        end
      else
        begin
          reg2072 = ($signed((7'h56)) ?
              (^~$unsigned({wire2043, (^reg1838)})) : ({{reg1768,
                      reg1832[(1'h1):(1'h1)]},
                  ($signed(reg2063) + (reg1883 || reg2010)),
                  {(~&reg2056), {reg1796}}} >= (~|$unsigned((7'h42)))));
          for (forvar2073 = (1'h0); (forvar2073 < (2'h2)); forvar2073 = (forvar2073 + (1'h1)))
            begin
              reg2075 <= reg1794[(5'h10):(3'h7)];
              reg2076 = (reg1768 ?
                  (reg2063[(2'h3):(2'h2)] <<< ($unsigned(reg1768) ?
                      $unsigned(reg1915) : $signed((forvar2073 >> (8'haf))))) : {$unsigned((~$signed(reg1825))),
                      (&$unsigned($signed((8'hba)))),
                      ((^~reg1933) ?
                          ({reg2075} ?
                              reg2009 : reg1806) : (reg2009[(3'h7):(2'h2)] ?
                              (|reg1914) : $unsigned(reg1769)))});
              reg2078 <= $unsigned((-(reg1829 ?
                  $unsigned($unsigned(reg1777)) : ((reg2049 ^ (8'hbd)) != (reg2015 & reg2062)))));
              reg2079 = (~|$signed((reg1903 ?
                  reg2002 : reg2081[(5'h13):(1'h0)])));
              reg2080 = reg1943;
              reg2082 <= (~&reg1940);
            end
        end
      reg2083 = $signed((reg1942 ?
          $signed(reg1814[(5'h11):(3'h5)]) : reg1825[(5'h13):(3'h5)]));
    end
  always
    @(posedge clk) begin
      for (forvar2084 = (1'h0); (forvar2084 < (3'h5)); forvar2084 = (forvar2084 + (1'h1)))
        begin
          for (forvar2085 = (1'h0); (forvar2085 < (1'h0)); forvar2085 = (forvar2085 + (1'h1)))
            begin
              reg2086 = (&(~($signed((reg1936 * (7'h4c))) ?
                  (reg2065[(4'h9):(3'h7)] ?
                      (reg2070 * (7'h44)) : $unsigned(reg2023)) : reg1811[(5'h11):(5'h10)])));
              reg2087 = $unsigned($signed((&(-$unsigned(reg1875)))));
              reg2088 <= (^~(~&reg1915));
              reg2089 = ((({$unsigned(reg1936)} ?
                      reg2006[(4'hd):(4'hd)] : reg1933[(4'hf):(3'h7)]) || (&reg1800)) ?
                  (8'ha8) : (reg1954 ?
                      $signed($signed($signed(reg2015))) : (reg1891 ^~ $signed(reg1857))));
              reg2090 = reg1818[(1'h0):(1'h0)];
              reg2091 <= reg1935;
              reg2092 = $signed($unsigned(($signed((|wire1761)) ?
                  reg2020[(5'h11):(5'h10)] : reg1822)));
            end
          reg2093 <= (-$signed((^~(reg1774[(4'hb):(4'hb)] ?
              (~reg2015) : $unsigned(reg1777)))));
          reg2094 <= (8'ha1);
          reg2095 <= $unsigned(((~($signed(reg1855) ?
                  (+reg1982) : $unsigned(reg1911))) ?
              {reg1860[(4'he):(4'h9)],
                  reg2091[(1'h1):(1'h1)],
                  {((8'hbd) >> reg1796)}} : (+(~|(reg2029 && reg1777)))));
          for (forvar2096 = (1'h0); (forvar2096 < (2'h2)); forvar2096 = (forvar2096 + (1'h1)))
            begin
              reg2097 <= $unsigned($unsigned(reg1846));
              reg2098 <= ((($signed(reg2042) ?
                          reg1771 : ((reg2091 >= reg1954) + (reg1893 || reg1818))) ?
                      $signed(((reg1995 >= (8'h9d)) || reg1796)) : $unsigned(reg1819[(1'h1):(1'h1)])) ?
                  $unsigned(reg1839) : ($signed(reg2092[(4'h9):(2'h3)]) ?
                      reg2090[(4'h8):(1'h0)] : $unsigned($signed($unsigned(reg1826)))));
            end
          for (forvar2099 = (1'h0); (forvar2099 < (3'h5)); forvar2099 = (forvar2099 + (1'h1)))
            begin
              reg2100 = $signed((~reg1869[(3'h5):(2'h3)]));
              reg2101 = $signed(({((reg2009 ? reg1768 : (8'h9e)) ?
                          (|reg1808) : {(8'hb5)}),
                      {$signed(reg1797),
                          {reg2053, reg1861},
                          (reg2070 ^~ (8'had))}} ?
                  $unsigned($unsigned(reg1900[(5'h17):(1'h1)])) : (~^$signed($signed((7'h56))))));
              reg2102 = reg1942;
            end
        end
      for (forvar2103 = (1'h0); (forvar2103 < (2'h2)); forvar2103 = (forvar2103 + (1'h1)))
        begin
          reg2104 <= reg1923;
          reg2105 = (~&$signed(((reg1877 ?
                  $signed(reg1783) : reg1832[(2'h2):(1'h0)]) ?
              $unsigned((&reg1979)) : (((7'h40) != reg2053) ^~ (!reg1875)))));
          if (reg2101)
            begin
              reg2106 = $signed($unsigned(($signed(reg2004[(1'h0):(1'h0)]) ?
                  $unsigned({reg2073}) : (reg1966 ^~ (reg1800 ?
                      reg2065 : reg1785)))));
              reg2107 <= (!reg2089[(2'h3):(1'h1)]);
              reg2108 <= {(reg1904 ?
                      (reg1935 ?
                          $unsigned((reg1868 ?
                              forvar2085 : reg1906)) : reg1993[(2'h3):(1'h0)]) : (!(^(reg2094 ?
                          (7'h55) : reg1903))))};
              reg2109 <= (~|reg1839[(4'h9):(3'h6)]);
              reg2110 <= $signed(reg1861);
              reg2111 <= {($unsigned(($unsigned(reg1993) << (&forvar2096))) ?
                      reg1923 : reg1940[(5'h10):(2'h2)])};
            end
          else
            begin
              reg2106 = reg2007[(5'h13):(4'hc)];
              reg2107 <= reg1990[(2'h2):(2'h2)];
              reg2112 = $unsigned($signed((7'h55)));
              reg2113 = reg1766[(1'h0):(1'h0)];
              reg2114 <= reg1966[(5'h12):(4'hb)];
            end
        end
      if (reg2071)
        begin
          if ((^reg2046[(4'hc):(4'h8)]))
            begin
              reg2115 <= ((reg2053[(5'h11):(4'hb)] ?
                  (reg1791[(2'h2):(1'h1)] + reg2017) : (reg1926[(3'h7):(1'h1)] ?
                      (reg1892 ?
                          (reg2107 == reg1904) : reg1978) : ($signed(reg1826) ?
                          reg1973[(5'h12):(4'h9)] : reg1926[(1'h0):(1'h0)]))) - $unsigned(reg1936));
              reg2116 <= ((&wire1896[(3'h5):(1'h0)]) ?
                  ({reg1822,
                      $signed((reg1915 < reg1893))} & (+(reg1998 << {(7'h45),
                      reg1885,
                      reg1892}))) : (~^reg1796));
              reg2117 <= $signed(reg2066);
              reg2118 <= $signed((~|{(+(reg2101 ? reg1791 : (8'h9e)))}));
              reg2119 = reg1999[(2'h2):(1'h1)];
            end
          else
            begin
              reg2115 <= $signed(reg1961);
            end
        end
      else
        begin
          if ($signed({reg1861[(2'h2):(1'h0)]}))
            begin
              reg2115 <= ({(7'h50),
                  reg2097,
                  (~|(reg1843 ?
                      reg2065[(4'he):(4'he)] : $signed(reg1950)))} | (~|{{reg2064,
                      reg2104[(1'h0):(1'h0)],
                      {reg1848}},
                  reg2004[(4'hc):(1'h0)],
                  (^~(8'ha6))}));
              reg2116 <= {reg2073};
              reg2119 = (reg2020 ?
                  {$unsigned((+wire1763[(2'h3):(1'h1)]))} : ($unsigned(((reg1943 ?
                          (8'ha1) : (7'h46)) ?
                      $signed(reg2023) : {reg2015,
                          (7'h53),
                          reg2010})) >> reg1962));
              reg2120 = ($unsigned(reg2102) > $unsigned(((reg1788 <<< reg1917[(4'hf):(3'h5)]) ?
                  reg1942[(3'h7):(2'h2)] : reg2082[(1'h0):(1'h0)])));
              reg2121 <= (^wire1765);
              reg2122 = ({{$signed((reg1943 ^~ wire1761)),
                      (reg1848[(1'h0):(1'h0)] ?
                          $signed(reg1819) : $signed((8'h9e))),
                      reg1806}} ^~ {reg2088[(4'ha):(4'h8)]});
              reg2123 = (reg1869[(1'h1):(1'h0)] + (reg1869 ?
                  (~$unsigned(forvar2096[(2'h2):(2'h2)])) : (reg1987[(4'h9):(3'h6)] ?
                      (&$unsigned((8'h9c))) : ({(8'hbe), (8'hbb), reg2116} ?
                          (|reg1981) : $signed(reg1940)))));
            end
          else
            begin
              reg2119 = reg1816[(5'h14):(4'h8)];
              reg2121 <= reg1977;
              reg2122 = $unsigned(reg2060);
              reg2124 <= (-((|$unsigned(reg1926[(3'h6):(3'h4)])) ?
                  $unsigned(reg1806) : {(reg1956[(4'h8):(1'h1)] - {reg1940}),
                      $unsigned((|reg1803))}));
              reg2125 = reg1912;
              reg2126 = (reg1940 <<< $signed((&reg1914[(5'h11):(4'hb)])));
            end
          reg2127 = $signed($signed(($unsigned({reg2071,
              reg1884}) <= (!$unsigned(reg2090)))));
          reg2128 = $signed(reg2052);
        end
      reg2129 = ($unsigned($unsigned((!$unsigned((7'h54))))) >>> (({reg1806} || ($unsigned(reg1768) + (~reg1797))) ?
          reg2001 : reg1788));
      if (((&$signed((~$signed(reg2028)))) ?
          (((+((8'h9c) ?
              (7'h51) : reg2067)) && (~&(reg1948 >= reg2002))) | (7'h52)) : (-(8'ha9))))
        begin
          reg2130 = {(!reg1769[(4'h8):(3'h7)]),
              $unsigned((reg1825 ?
                  (~&reg2004[(1'h0):(1'h0)]) : ($signed(reg1796) ?
                      ((8'ha6) <= reg1917) : $signed(reg1766)))),
              reg1838[(5'h12):(5'h12)]};
          for (forvar2131 = (1'h0); (forvar2131 < (1'h0)); forvar2131 = (forvar2131 + (1'h1)))
            begin
              reg2132 <= {$signed((($unsigned(reg1825) ?
                          $unsigned((8'hbe)) : (8'haf)) ?
                      reg2007[(5'h18):(5'h17)] : $unsigned((reg1806 ?
                          reg2105 : reg2071)))),
                  (&((reg1768[(4'hd):(2'h3)] && (reg2070 >>> forvar2099)) ^ reg2047)),
                  ((^~reg1990) ?
                      reg1956[(5'h11):(4'h8)] : ({(reg2110 ? reg1797 : reg2125),
                          reg2004[(1'h1):(1'h1)]} ^ reg1836[(1'h0):(1'h0)]))};
              reg2133 = ((!$signed(($signed(reg1962) ?
                  (reg1914 || forvar2103) : $unsigned((8'ha6))))) ^ (8'hbe));
              reg2134 = ((reg1803 && ((reg1843[(2'h2):(2'h2)] ?
                          (reg2018 ? reg1796 : reg2132) : $signed(reg2089)) ?
                      (!reg2065[(5'h14):(3'h7)]) : reg1818[(3'h4):(2'h2)])) ?
                  (reg2117[(4'h8):(1'h0)] + $signed(($unsigned((7'h40)) ?
                      reg1783 : reg1906))) : (~&reg1948[(2'h3):(1'h1)]));
            end
        end
      else
        begin
          reg2131 <= ($unsigned(reg1950[(4'hf):(4'hd)]) >> $signed({($signed((7'h48)) ?
                  wire1760[(4'hc):(3'h5)] : reg2039),
              $signed((reg2028 < reg1774)),
              $unsigned(reg2091)}));
          reg2133 = reg2128;
          reg2135 <= $unsigned($unsigned(reg2020[(5'h17):(1'h1)]));
          if (({(wire1896[(3'h4):(2'h2)] ?
                  reg2129 : $signed((reg2134 ? reg2095 : (8'hab)))),
              (8'hb3)} << {(&(^(-reg1833)))}))
            begin
              reg2136 <= $unsigned(((~&((reg2067 ?
                      (7'h48) : reg1926) << $unsigned(reg2082))) ?
                  reg2093[(1'h0):(1'h0)] : $unsigned((forvar2103[(5'h10):(4'h8)] ?
                      (reg2009 >= reg2046) : $unsigned(reg2030)))));
              reg2137 = ($signed((reg1826[(3'h4):(1'h1)] <<< reg2010[(1'h1):(1'h1)])) >>> (&((~&reg1982) ?
                  $signed($signed(forvar2131)) : (8'hb3))));
              reg2138 = ($unsigned((reg1794 ~^ ((reg1775 ?
                      reg1806 : reg1816) != reg2121[(3'h5):(2'h3)]))) ?
                  $unsigned(({(7'h53)} <= (reg1839[(3'h4):(2'h3)] ?
                      reg1855[(1'h1):(1'h1)] : (7'h41)))) : ($unsigned($unsigned($unsigned((8'haf)))) != ($signed(reg1884[(3'h6):(1'h1)]) ?
                      (((7'h41) == reg2115) <= reg2117) : $signed($signed(reg2114)))));
              reg2139 = (~&({$unsigned($signed(reg1806))} && (^(7'h53))));
              reg2140 = $unsigned($unsigned($signed((reg1804[(2'h2):(2'h2)] && (reg1839 ~^ reg1936)))));
              reg2141 = ({$unsigned(reg2107[(3'h4):(2'h3)]),
                  (8'hba),
                  {reg2086[(2'h2):(1'h1)],
                      ((&reg1954) ?
                          (reg2109 ?
                              (8'hb1) : reg1848) : $signed(reg2122))}} & reg2102[(1'h0):(1'h0)]);
            end
          else
            begin
              reg2137 = $signed($unsigned({(~^(|reg2098)),
                  {(reg1797 ? reg1982 : reg1956), $unsigned(wire1763)},
                  $unsigned(reg2130)}));
              reg2138 = $unsigned($signed(((-reg1914) || reg2111)));
              reg2142 <= {{(((|reg2113) ?
                              (reg2115 ^ (7'h53)) : ((8'hb8) >= reg2002)) ?
                          $signed($unsigned(reg1999)) : (8'ha3)),
                      (((reg2108 | wire1765) | reg1885) ?
                          {{reg1880}} : ($unsigned(reg1848) ?
                              {reg1967, reg2093} : wire1761))}};
              reg2143 <= (($unsigned($unsigned((reg1811 ?
                      (8'hb9) : reg2116))) + (($unsigned(reg1804) >> $unsigned((7'h46))) != ($signed(reg2073) && reg1926))) ?
                  ((^reg2121[(2'h2):(1'h0)]) ?
                      $signed((^reg2124[(4'hd):(4'hc)])) : ($signed(((7'h45) ?
                              reg1932 : reg2048)) ?
                          $unsigned(reg1948[(2'h2):(1'h0)]) : $signed({wire1765,
                              (8'had)}))) : (reg2000 < reg2117[(4'hd):(3'h4)]));
              reg2144 = (~^((-$unsigned(reg1818)) & (8'ha5)));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2145 = (1'h0); (forvar2145 < (1'h1)); forvar2145 = (forvar2145 + (1'h1)))
        begin
          reg2146 = $signed($signed(($unsigned({reg2131}) ^ ((wire1761 ?
              reg2014 : reg1819) ~^ {reg1880, (8'hb2)}))));
          for (forvar2147 = (1'h0); (forvar2147 < (1'h0)); forvar2147 = (forvar2147 + (1'h1)))
            begin
              reg2148 <= $unsigned(reg1857[(2'h2):(1'h1)]);
              reg2149 <= reg1875[(3'h5):(1'h1)];
              reg2150 <= (+reg1956);
              reg2151 <= (|$unsigned(reg2063));
            end
          if ($unsigned(reg1869[(2'h2):(1'h1)]))
            begin
              reg2152 <= $unsigned($signed($signed($unsigned(reg2009[(1'h1):(1'h1)]))));
              reg2153 <= $signed((+(7'h46)));
            end
          else
            begin
              reg2152 <= $signed(reg1790);
              reg2154 = reg2124[(4'he):(4'h9)];
              reg2155 = $signed($unsigned(reg1768));
              reg2156 = (|((+reg2023) - (($unsigned(reg1885) <= reg1905[(1'h0):(1'h0)]) >>> {{reg2016,
                      forvar2145},
                  $signed(reg1900)})));
              reg2157 = {$unsigned(reg1785),
                  (-(|$signed({reg2000, reg1775, reg1884}))),
                  {({(~|reg1917), reg1892, {reg1868, reg1819, reg1790}} ?
                          (reg2109[(4'h9):(4'h9)] || (reg2053 - reg1982)) : (wire1760[(2'h3):(2'h3)] <<< (reg2135 || reg1808))),
                      (($unsigned(reg2009) ?
                              reg2046[(4'h9):(3'h6)] : (|reg2015)) ?
                          $unsigned((-reg2046)) : ($unsigned((8'haa)) || (reg1967 ?
                              reg1836 : reg1948)))}};
            end
          for (forvar2158 = (1'h0); (forvar2158 < (1'h1)); forvar2158 = (forvar2158 + (1'h1)))
            begin
              reg2159 = (wire1765[(2'h3):(1'h1)] > (^$unsigned($unsigned(reg2155[(1'h0):(1'h0)]))));
              reg2160 <= ({$unsigned((|reg2062)),
                      $unsigned((-reg1800[(3'h6):(3'h5)]))} ?
                  $unsigned($unsigned(wire1896[(3'h5):(2'h2)])) : reg1775);
              reg2161 <= reg1962[(3'h4):(2'h2)];
              reg2162 = $unsigned(reg2054);
              reg2163 = reg2001[(3'h6):(2'h3)];
              reg2164 = reg1946;
              reg2165 <= reg1917;
            end
        end
      if ($signed((7'h47)))
        begin
          for (forvar2166 = (1'h0); (forvar2166 < (2'h2)); forvar2166 = (forvar2166 + (1'h1)))
            begin
              reg2167 = (&$unsigned((wire1765 ?
                  reg2004[(5'h10):(1'h0)] : ((reg1923 | reg1788) < $signed((7'h4a))))));
              reg2168 <= $signed($unsigned(reg1911));
              reg2169 <= reg2097;
              reg2170 = ((8'ha5) ? reg2135 : (reg1979 | reg1785));
            end
          reg2171 <= reg2121;
          if (reg1990)
            begin
              reg2172 = $unsigned(((((reg2156 == reg1892) ?
                      $unsigned(reg2014) : $unsigned(reg2160)) ?
                  $unsigned(reg2071) : {(&forvar2147)}) ^~ (reg2097[(5'h19):(4'hc)] ?
                  ({(7'h55), reg2163} ?
                      reg2065 : (reg1893 == reg1848)) : ($unsigned(reg2000) ?
                      $unsigned(wire1763) : $unsigned((7'h40))))));
              reg2173 = $signed((&reg1803[(2'h2):(1'h1)]));
            end
          else
            begin
              reg2172 = ({($unsigned((reg2066 >>> wire1762)) ^~ reg2017),
                      ((8'hbf) ^ reg1869),
                      (~&((reg2028 ? reg1791 : reg1829) <= $signed((8'ha2))))} ?
                  ((~&(~^(8'h9e))) ?
                      ({$unsigned(reg1869),
                              (^reg1982),
                              (reg1940 ? reg2104 : (8'ha6))} ?
                          reg1860 : {reg2028[(1'h1):(1'h1)]}) : ($signed((reg2148 ?
                          reg2009 : reg2070)) << reg2010)) : $signed((!reg1950[(5'h1c):(4'hb)])));
            end
          reg2174 = (!(&$signed(((reg1956 & (7'h58)) ?
              (reg1768 ? reg1993 : wire1765) : reg1884))));
          if ((reg1825 < reg2027))
            begin
              reg2175 <= ((reg2157 ?
                  $unsigned(($unsigned(reg2052) ?
                      $signed(reg2053) : $unsigned(reg2167))) : (reg2028 ?
                      $unsigned((reg2027 >>> reg2000)) : ($unsigned(reg1928) ^~ reg1923))) >= $unsigned(({((8'hbb) ?
                          reg2042 : reg1864),
                      $unsigned(reg2073)} ?
                  reg2159[(5'h10):(4'h8)] : $signed(((7'h46) + reg1977)))));
              reg2176 <= $signed((~^(~^reg2136[(2'h3):(1'h1)])));
              reg2177 <= reg2149[(5'h14):(5'h11)];
            end
          else
            begin
              reg2175 <= reg1902[(3'h4):(1'h1)];
              reg2176 <= $unsigned(((reg2114[(1'h1):(1'h1)] ?
                  reg2121[(3'h5):(1'h0)] : (reg1788 <<< (reg2132 ?
                      reg2037 : reg1991))) ~^ reg1940[(1'h1):(1'h0)]));
              reg2177 <= ((reg1978 <= $unsigned(reg1928[(2'h2):(1'h0)])) <<< (!$unsigned(((8'hac) ?
                  (reg1995 < reg2053) : reg1824[(1'h0):(1'h0)]))));
              reg2178 = $signed(reg2151);
              reg2179 = ((~^reg2028) ?
                  $signed(reg2154) : $signed((!(reg2067[(3'h7):(2'h2)] ?
                      reg2175[(4'ha):(3'h6)] : reg2110[(5'h11):(3'h5)]))));
            end
        end
      else
        begin
          for (forvar2166 = (1'h0); (forvar2166 < (3'h4)); forvar2166 = (forvar2166 + (1'h1)))
            begin
              reg2167 = reg2114;
            end
          if ((reg2098 ?
              $signed(($signed((reg2157 ?
                  (7'h48) : reg1928)) <= $unsigned((reg2037 ?
                  (7'h54) : reg2143)))) : reg1838[(4'he):(3'h4)]))
            begin
              reg2168 <= reg2027;
              reg2169 <= {{$unsigned(((reg2142 | (8'ha3)) ?
                          $signed(reg2148) : (~|reg1902))),
                      $signed($unsigned(reg1816[(3'h6):(1'h0)])),
                      (8'hb4)},
                  ((~|$unsigned(reg2017[(2'h2):(1'h0)])) >= reg2131)};
              reg2171 <= $unsigned(reg1777);
            end
          else
            begin
              reg2170 = ((~^(~|$signed((reg1886 > reg1777)))) ^ forvar2147[(5'h10):(4'hb)]);
              reg2172 = (-reg1860);
              reg2175 <= $unsigned($signed({(!$signed(reg1848)),
                  (~^reg1894),
                  $unsigned($unsigned((8'hac)))}));
              reg2178 = (reg2161[(1'h0):(1'h0)] >>> (($unsigned(reg1846[(3'h7):(2'h2)]) && reg1839) != reg1914[(4'hc):(2'h2)]));
              reg2180 <= ($unsigned(reg2065) <<< $unsigned((-$signed((reg2148 <<< (7'h56))))));
              reg2181 = reg2176[(5'h11):(3'h4)];
            end
          for (forvar2182 = (1'h0); (forvar2182 < (1'h1)); forvar2182 = (forvar2182 + (1'h1)))
            begin
              reg2183 = reg1861;
              reg2184 = $unsigned((reg2042[(2'h2):(1'h0)] ?
                  reg1900 : $signed(reg2073)));
              reg2185 = (reg1950 * reg2135[(4'h8):(3'h6)]);
              reg2186 = $unsigned((7'h40));
              reg2187 <= (((-($signed((8'hb9)) || reg1897[(3'h6):(1'h0)])) >= $unsigned(reg2071[(2'h3):(2'h2)])) != reg2170);
              reg2188 = ((reg2107 <= $unsigned(reg1869[(1'h0):(1'h0)])) ^ (~&{((reg2098 * reg2170) ?
                      reg1905[(2'h3):(2'h2)] : (reg2150 != forvar2145))}));
              reg2189 = reg1846;
            end
          for (forvar2190 = (1'h0); (forvar2190 < (3'h4)); forvar2190 = (forvar2190 + (1'h1)))
            begin
              reg2191 = (reg1783[(3'h7):(3'h5)] ?
                  (+(({reg1836} ?
                      $unsigned(reg1838) : $signed(reg1956)) != $signed((reg2151 ?
                      reg1961 : reg2107)))) : (^~(($signed(reg1860) ?
                      reg1840 : (reg2030 ?
                          reg1892 : reg1942)) + (reg2111 <<< (reg1799 == reg2037)))));
              reg2192 = $signed((~&$signed(((reg2179 ? (8'hab) : reg1804) ?
                  reg2169[(5'h13):(3'h4)] : (reg2116 ? reg1936 : reg1814)))));
              reg2193 = $signed({($unsigned(reg1785[(3'h5):(2'h2)]) ?
                      ((reg1950 == reg1946) ?
                          (reg1811 + reg1979) : {reg1775,
                              (8'hb0),
                              (7'h47)}) : (reg1902 == $signed(reg1894)))});
              reg2194 <= reg1995[(5'h10):(4'hc)];
              reg2195 <= forvar2145[(3'h4):(1'h0)];
            end
          reg2196 <= (($unsigned(reg2030[(4'hb):(3'h6)]) <= reg2131) - reg2023);
          for (forvar2197 = (1'h0); (forvar2197 < (3'h6)); forvar2197 = (forvar2197 + (1'h1)))
            begin
              reg2198 <= (^~$unsigned({({forvar2190,
                      reg1803,
                      reg2181} >> (wire1762 ? reg2157 : reg1891))}));
              reg2199 = reg2030[(5'h12):(5'h10)];
              reg2200 <= $signed(($unsigned(reg2136[(3'h5):(1'h0)]) ?
                  $signed((^((8'had) << reg2002))) : {((~&reg2062) ?
                          reg1956[(4'h9):(2'h3)] : $unsigned(reg2015)),
                      reg2198[(4'h8):(2'h3)],
                      (reg2030[(2'h2):(1'h1)] ?
                          $unsigned((7'h48)) : (^~(7'h4a)))}));
              reg2201 = reg2065[(4'h8):(3'h4)];
              reg2202 = $unsigned(reg2200);
              reg2203 = reg1886;
            end
        end
      for (forvar2204 = (1'h0); (forvar2204 < (2'h2)); forvar2204 = (forvar2204 + (1'h1)))
        begin
          for (forvar2205 = (1'h0); (forvar2205 < (2'h2)); forvar2205 = (forvar2205 + (1'h1)))
            begin
              reg2206 = (reg1935 ? reg1864 : reg1982[(3'h7):(3'h4)]);
            end
        end
    end
  assign wire2207 = reg1961;
  assign wire2208 = ($signed((^$signed($signed(reg1962)))) && (&(7'h4a)));
  always
    @(posedge clk) begin
      if (reg2017[(3'h6):(2'h3)])
        begin
          for (forvar2209 = (1'h0); (forvar2209 < (3'h6)); forvar2209 = (forvar2209 + (1'h1)))
            begin
              reg2210 <= (reg1829 < reg1915);
              reg2211 = reg2023[(4'hb):(4'h9)];
              reg2212 = {(($unsigned(reg1962) ?
                          (~|(7'h52)) : ($unsigned(reg1788) ^ reg2095)) ?
                      reg1946[(3'h4):(2'h2)] : reg2151),
                  $signed((|{$unsigned((8'hba)), reg1840}))};
              reg2213 = (8'had);
            end
          if ($unsigned(({(^~$unsigned(reg1892)),
              {reg1966},
              ((reg2007 ? reg1869 : reg2052) ?
                  (reg1905 ? reg1811 : (7'h4e)) : {(8'hbe),
                      reg2180})} & $unsigned($signed((~&reg1942))))))
            begin
              reg2214 <= (+$unsigned($signed($unsigned(reg2007[(5'h16):(5'h11)]))));
              reg2215 <= {($unsigned((reg2057 ?
                          $unsigned(reg2066) : $unsigned(reg2111))) ?
                      $unsigned((reg2165 ?
                          $signed(reg2030) : (wire2207 >> reg1966))) : reg2165)};
              reg2216 <= ($unsigned(((reg2020[(4'h9):(4'h9)] << (reg1804 ?
                      reg2017 : reg2075)) ?
                  ((wire1760 > (8'hb2)) - (~&reg2153)) : (wire1761 | (reg2071 ?
                      reg1875 : reg2009)))) >= $signed($signed($signed((8'haf)))));
              reg2217 <= reg1848;
              reg2218 <= {((+{$signed(reg1981),
                          (reg1868 ? reg2110 : reg2152),
                          (reg1973 != reg1942)}) ?
                      (($signed(reg2198) ?
                          reg1818 : $signed((8'hae))) - $signed({reg1923})) : (8'hb6))};
            end
          else
            begin
              reg2219 = $signed(($unsigned(reg1806) ?
                  (-{(^~wire1761),
                      reg1796}) : $unsigned($unsigned(reg1799[(5'h17):(5'h16)]))));
            end
          reg2220 <= reg2001[(1'h0):(1'h0)];
          if (($unsigned(((reg2118[(2'h3):(2'h2)] + (reg1908 << reg1892)) ?
                  (~^$unsigned(reg2121)) : reg2117[(3'h5):(3'h4)])) ?
              $signed((~|(+$signed(reg2169)))) : $signed((((reg2078 | reg2049) * $signed(reg1973)) ?
                  reg2131 : ((^~reg1985) ?
                      {reg1785, reg1803} : (reg1855 & (7'h51)))))))
            begin
              reg2221 <= $unsigned(reg1993[(4'hc):(2'h2)]);
            end
          else
            begin
              reg2221 <= $signed(reg1961);
              reg2222 = reg2213;
            end
          reg2223 <= ((({reg1985[(3'h6):(3'h5)]} ?
                  $unsigned(((7'h4e) ? reg1840 : reg1905)) : reg1766) ?
              $unsigned(reg1811) : $signed(($signed(reg1897) ?
                  reg1915[(2'h3):(1'h1)] : reg1885[(1'h1):(1'h0)]))) & (((~&$signed(reg2213)) ?
                  reg1981[(4'hc):(3'h4)] : reg2108) ?
              $signed($signed({reg2064, reg1766})) : {$unsigned((~^reg2037)),
                  $unsigned((reg2098 ? reg2161 : reg1791)),
                  reg2196[(3'h6):(1'h0)]}));
          if ($unsigned((!forvar2209[(4'hc):(4'ha)])))
            begin
              reg2224 <= $signed((|$signed((reg1905 ?
                  {reg2118, (7'h52), reg2221} : $signed(reg1808)))));
              reg2225 = ($unsigned($unsigned($unsigned($signed(reg2016)))) && ($signed(reg1906[(2'h2):(2'h2)]) ?
                  $unsigned($signed(reg1987)) : reg2002[(1'h1):(1'h0)]));
              reg2226 <= $unsigned({$signed(($unsigned(reg2187) ?
                      (reg1857 + reg1788) : $unsigned(reg2198)))});
              reg2227 = {$unsigned($signed((reg1824[(1'h1):(1'h1)] ^~ reg2116)))};
              reg2228 = $signed((&{((~&(8'ha9)) | {reg1855})}));
            end
          else
            begin
              reg2225 = (~{(reg2153 >>> ($signed(forvar2209) >> ((7'h50) <= (8'ha8)))),
                  $signed({$unsigned(reg2049)}),
                  {$unsigned(((7'h41) ? reg2088 : reg1891))}});
              reg2227 = ($signed($unsigned($signed({reg1833}))) ?
                  reg2222 : $unsigned(({$unsigned(reg2048),
                      $unsigned(reg2219)} >> reg2052[(4'hb):(2'h2)])));
              reg2229 <= $unsigned((((reg1956[(1'h1):(1'h0)] != reg2152[(3'h4):(1'h1)]) ^~ ((reg2131 >> reg2067) | reg2121[(3'h4):(1'h0)])) ?
                  ({$signed(reg1832)} ?
                      $unsigned($signed(reg2180)) : reg2002[(2'h2):(1'h1)]) : $unsigned($unsigned((reg2227 ?
                      reg1897 : reg1868)))));
              reg2230 = reg2224[(3'h6):(2'h2)];
              reg2231 <= $signed($signed(reg2117));
              reg2232 = (~^(~|reg2056[(3'h4):(3'h4)]));
              reg2233 = reg1791;
            end
        end
      else
        begin
          if ((+$unsigned(({(~reg1824),
              $unsigned(reg2029)} < reg2225[(5'h14):(5'h12)]))))
            begin
              reg2209 <= reg2180;
              reg2210 <= reg1768[(2'h3):(1'h0)];
              reg2214 <= reg2095;
            end
          else
            begin
              reg2209 <= ($signed(((!$signed(reg1908)) < $signed($unsigned((8'hb9))))) ?
                  (reg1897 || $unsigned((reg2229[(5'h13):(4'ha)] <= reg1954[(2'h2):(2'h2)]))) : $unsigned((~|reg1840)));
              reg2211 = ({(reg2115 ?
                      $unsigned($unsigned(reg2073)) : $signed(reg2224)),
                  (-$unsigned({reg1766, (7'h42)}))} >>> reg2073[(2'h2):(2'h2)]);
              reg2212 = ($unsigned($signed($unsigned((reg1800 ?
                  reg1878 : reg2082)))) ~^ {{($unsigned(reg1839) ?
                          {(7'h47)} : reg2056[(4'ha):(4'ha)]),
                      ({(7'h58), reg2115} >> $unsigned(reg1966))},
                  reg1993[(4'hf):(1'h0)]});
              reg2214 <= (reg2152 >= (reg2078[(5'h13):(5'h11)] ?
                  $unsigned(reg1886) : reg2057));
              reg2219 = reg2222;
            end
          reg2222 = (~|(^~(~|(~(reg2028 ? reg2230 : reg1811)))));
          for (forvar2223 = (1'h0); (forvar2223 < (2'h3)); forvar2223 = (forvar2223 + (1'h1)))
            begin
              reg2225 = reg2046;
              reg2227 = ((+((~|$signed(reg2161)) ?
                  (reg2148 ?
                      $unsigned((7'h48)) : (~|reg2109)) : (reg1943[(1'h0):(1'h0)] == reg1948[(1'h1):(1'h1)]))) >>> ($unsigned({(reg2098 ?
                          forvar2223 : reg1917),
                      (^reg2067)}) ?
                  ((reg1892 ?
                          $signed((8'hb0)) : ((8'haa) ? reg2049 : reg1885)) ?
                      (^(8'hb5)) : (~reg2071)) : $signed({$signed(reg1917),
                      (reg2018 ? wire1762 : reg2161),
                      $unsigned(reg1814)})));
              reg2228 = reg1961;
              reg2229 <= (^$signed($signed($unsigned((^reg2215)))));
              reg2231 <= (-(~|reg1797[(5'h11):(4'hd)]));
              reg2234 <= $signed(reg1828);
            end
        end
      reg2235 = ((~reg2220[(3'h5):(3'h5)]) * $unsigned($unsigned({$unsigned((8'h9f)),
          $signed(reg2071),
          (^~reg2088)})));
      if ((reg1857[(1'h0):(1'h0)] ^~ $signed(reg2067[(3'h5):(3'h4)])))
        begin
          reg2236 = {((($unsigned(reg1769) > (~|reg1819)) == $unsigned({reg1905,
                      reg1961})) ?
                  $signed(((~^(8'hb5)) <<< reg1883)) : $signed(($unsigned(reg1962) ^ (reg2073 ?
                      (7'h4a) : reg1774)))),
              (($signed((^reg2007)) ?
                  reg2219 : reg1878) + reg2230[(4'hb):(4'h8)])};
          reg2237 = (-reg2073[(2'h2):(1'h1)]);
          reg2238 <= reg1905[(2'h3):(2'h2)];
          if ((reg2046 ?
              {$signed(((reg2097 > reg1915) ? (~reg2107) : $unsigned(reg2211))),
                  (~|$signed(reg1906))} : ((~&$unsigned((reg2148 ?
                  reg1777 : reg2221))) <= (reg1982[(5'h14):(5'h11)] | $signed($unsigned(reg2211))))))
            begin
              reg2239 = ((reg1775[(3'h4):(1'h1)] ?
                  reg1979[(2'h3):(2'h3)] : $signed($signed({reg2160}))) <= reg1978);
              reg2240 <= {($unsigned((8'ha2)) ?
                      reg2136 : (+((7'h46) ?
                          {(7'h4f), (7'h4c), reg2198} : {(8'ha2)}))),
                  (&reg2064),
                  $unsigned($unsigned($unsigned((!reg2177))))};
              reg2241 <= {{reg1832[(2'h2):(1'h0)],
                      $signed(((|reg2108) >= $signed(reg2237))),
                      ((8'ha5) ?
                          reg2042[(4'h8):(2'h3)] : (reg2020 ?
                              (|reg2136) : (reg1777 << reg2038)))},
                  reg2023};
              reg2242 <= (!(~|{{reg1832,
                      (reg2020 ? reg2065 : (8'hb6)),
                      $unsigned(reg2073)},
                  {(reg2067 ? reg2212 : (7'h54))},
                  $signed(reg1967)}));
              reg2243 <= $signed((~|{(^$signed(reg2091)),
                  ($unsigned((7'h4b)) * {reg1833, (8'h9f), (7'h55)}),
                  reg1923[(1'h0):(1'h0)]}));
              reg2244 <= $signed(reg2243[(1'h0):(1'h0)]);
            end
          else
            begin
              reg2239 = $unsigned(reg1766[(3'h6):(1'h0)]);
              reg2245 = $signed((~&reg1987[(4'h8):(3'h7)]));
              reg2246 = {reg2065};
            end
          reg2247 = reg2054[(4'h9):(2'h3)];
        end
      else
        begin
          if ($unsigned(reg2018[(3'h6):(1'h0)]))
            begin
              reg2238 <= ((~|{reg2116[(2'h2):(1'h0)]}) | reg1853[(2'h3):(1'h0)]);
              reg2239 = reg2224;
              reg2240 <= (!($unsigned($signed((reg2148 != reg2238))) && (~|reg1843)));
              reg2245 = {{reg1788, (-(-(reg1818 >>> reg1977)))}, reg2121};
              reg2248 <= {(reg1926 ? (~&reg2195) : reg2245)};
              reg2249 <= $unsigned(($signed($unsigned($unsigned((8'had)))) ?
                  ({reg1816[(4'hf):(1'h1)],
                          $signed((7'h55)),
                          (reg1829 << wire2043)} ?
                      {reg2245} : $unsigned((~|reg2245))) : reg2196));
              reg2250 <= (|reg1825[(4'hf):(1'h1)]);
            end
          else
            begin
              reg2236 = {((8'hab) ^ $signed($signed((reg1990 ?
                      reg2247 : reg2176))))};
              reg2238 <= (&wire2207);
              reg2239 = reg2095;
              reg2245 = $unsigned(($unsigned((reg2042[(3'h5):(1'h1)] << (reg2171 ?
                      reg1981 : reg1915))) ?
                  $signed(reg2121[(4'hc):(3'h4)]) : $signed(({reg1886,
                      reg2020} >= reg1990[(1'h0):(1'h0)]))));
              reg2248 <= $unsigned($signed(reg1782[(5'h11):(5'h10)]));
              reg2251 = $unsigned((~^reg2010));
            end
          reg2252 <= {reg1833[(5'h10):(4'ha)],
              (^~$signed((~^reg2229))),
              reg2108};
          reg2253 = reg1906[(3'h4):(1'h0)];
          for (forvar2254 = (1'h0); (forvar2254 < (3'h4)); forvar2254 = (forvar2254 + (1'h1)))
            begin
              reg2255 <= ($unsigned(wire2207[(4'hb):(1'h0)]) | (((~|(forvar2223 ?
                  reg1804 : reg2021)) <= reg1928[(5'h10):(4'h8)]) && $signed(reg1811)));
              reg2256 = (~|$unsigned((reg1990 ?
                  ((^~reg1790) ?
                      reg1833[(5'h1a):(5'h15)] : $unsigned(reg2233)) : wire2207)));
              reg2257 = reg2242[(5'h19):(2'h3)];
              reg2258 <= ((~|$unsigned(reg2097[(5'h12):(4'hb)])) > $signed((($signed(reg1847) ?
                      $signed(reg2010) : {(7'h41)}) ?
                  reg1886[(1'h1):(1'h0)] : reg1905)));
              reg2259 = {($signed(reg1848[(1'h1):(1'h0)]) ?
                      (((reg2056 & (8'ha0)) >> reg1990[(2'h2):(1'h1)]) ?
                          ($unsigned(reg1861) <= reg1902) : (~&$unsigned(reg1840))) : reg2121),
                  reg2016,
                  ((((reg2240 * reg2149) ?
                          (reg1935 ?
                              wire1760 : (7'h4a)) : reg2210[(5'h18):(2'h2)]) >> {reg2075,
                          (~reg1788),
                          reg2094}) ?
                      ({(reg2228 ^ reg2065),
                              (reg2115 != reg2143),
                              (reg1880 ? reg2014 : reg1838)} ?
                          ({reg2149, (8'hab), reg1814} >>> (reg1935 ?
                              (7'h42) : reg1967)) : $signed($unsigned(reg1981))) : ($unsigned($unsigned(reg2018)) ?
                          ($signed(reg1948) != (reg2107 ?
                              reg2143 : reg2241)) : $unsigned({(7'h4e),
                              (8'ha7)})))};
            end
        end
      if ({(reg2116[(3'h4):(3'h4)] ?
              (~&(reg2136[(1'h1):(1'h1)] ?
                  ((8'ha9) == reg1769) : $unsigned(reg2256))) : (-($unsigned((8'ha5)) <= $unsigned(reg1886)))),
          $signed((~&(!((8'ha8) ? reg2016 : forvar2254)))),
          ({$unsigned((wire1760 * reg2000)),
                  ({reg2253} ? (reg2136 ? reg1894 : reg2017) : {reg2237}),
                  reg2004} ?
              $unsigned({{reg2194, reg1846, reg1923}}) : reg2042)})
        begin
          for (forvar2260 = (1'h0); (forvar2260 < (3'h6)); forvar2260 = (forvar2260 + (1'h1)))
            begin
              reg2261 = reg2111;
              reg2262 <= (~&{reg2180});
              reg2263 <= reg1840;
              reg2264 <= (-{reg2056,
                  (+$signed((reg2258 ? reg1840 : reg2230)))});
              reg2265 <= $unsigned(($unsigned($unsigned(reg1875)) ?
                  $unsigned((~|((7'h47) ?
                      reg2108 : (8'hba)))) : {(~&(reg2228 | reg1991)),
                      $unsigned($signed(reg2023)),
                      reg2094}));
              reg2266 = $signed((reg1977 ?
                  reg2009[(4'ha):(1'h1)] : $unsigned((wire2043 ?
                      $unsigned(reg1766) : reg2020))));
            end
          reg2267 = $signed($unsigned(reg2245[(4'hf):(4'h9)]));
          reg2268 <= reg1846[(5'h10):(4'h9)];
          reg2269 = $signed($signed(($signed({reg2211, (8'had), reg1998}) ?
              (reg2094[(3'h7):(3'h7)] ?
                  $unsigned(reg2231) : (reg2027 != reg2258)) : reg1928)));
          reg2270 <= $signed(reg1932);
          reg2271 <= reg2104[(1'h1):(1'h1)];
        end
      else
        begin
          if (reg1908)
            begin
              reg2260 <= (((((reg1797 ? reg2060 : reg1900) != {(8'h9f),
                  (7'h58),
                  reg2030}) | reg2121) >= $unsigned({(reg2171 - (8'hb1))})) - reg2108);
              reg2262 <= reg2194;
              reg2263 <= (reg1991 ^ reg1768);
              reg2266 = {reg2114};
              reg2268 <= $unsigned(((((reg1869 ?
                      reg1995 : (8'ha3)) != (wire1765 << reg2150)) ^ reg2253) ?
                  reg2023[(4'he):(2'h3)] : ((^reg1911[(4'hf):(1'h1)]) * ($unsigned(reg2222) ?
                      {(7'h4a), reg1885} : reg1839[(4'ha):(3'h6)]))));
              reg2269 = reg2241[(4'he):(3'h4)];
              reg2270 <= $unsigned(($unsigned({(reg1885 ^~ reg2006),
                      reg1840[(2'h2):(2'h2)]}) ?
                  (reg1933[(1'h0):(1'h0)] ?
                      (8'ha7) : (((8'hb2) ? reg2109 : reg2110) ?
                          $signed(reg2261) : (reg1839 ?
                              reg2132 : reg2153))) : (reg1904 ?
                      $signed($signed(reg1788)) : (8'hb6))));
            end
          else
            begin
              reg2261 = reg2030[(4'hf):(4'hb)];
              reg2262 <= $unsigned(reg2038);
              reg2266 = reg2269[(3'h6):(3'h5)];
              reg2267 = $signed(($signed(reg2212) ?
                  ((reg1766[(3'h5):(1'h0)] > $signed(reg2243)) ?
                      reg1954 : (|$unsigned((7'h56)))) : reg2194));
              reg2268 <= $unsigned(({$unsigned($unsigned(reg2211)),
                  $unsigned((&reg2252))} < (+$signed((reg1885 ?
                  reg2224 : wire1764)))));
              reg2269 = $signed(($signed({$signed(reg1991)}) ?
                  $unsigned(($unsigned(reg2224) ?
                      $unsigned(reg2261) : reg1962[(3'h5):(3'h4)])) : reg1904));
              reg2272 = reg1884[(4'h9):(3'h7)];
            end
          reg2273 = $signed($signed($signed(reg2171)));
          for (forvar2274 = (1'h0); (forvar2274 < (3'h6)); forvar2274 = (forvar2274 + (1'h1)))
            begin
              reg2275 <= (~&$unsigned({{{reg2253}, (8'hab), (&wire1760)}}));
              reg2276 = ((|{reg2017[(4'h9):(2'h2)]}) ?
                  $signed($signed({reg1897,
                      reg2220,
                      $signed(reg1848)})) : (&(($signed(reg2217) <<< $unsigned((8'hb0))) ?
                      (~reg2149[(4'hc):(4'hc)]) : reg2169[(4'h8):(2'h2)])));
              reg2277 = reg1833;
              reg2278 = ($signed($signed(reg2136[(3'h6):(2'h3)])) ?
                  reg2056 : $signed({$unsigned(reg1814)}));
              reg2279 <= $signed(((reg2250[(5'h1c):(5'h11)] ^~ ({reg1811,
                          reg1935,
                          wire1761} ?
                      {(8'hbe), reg2276} : $unsigned(reg2063))) ?
                  (+$unsigned($signed(reg2217))) : $unsigned((8'hab))));
              reg2280 = reg1908[(3'h6):(3'h6)];
              reg2281 = (|$signed(($unsigned(reg1999) ?
                  reg2030[(4'hc):(3'h4)] : $signed($unsigned(reg2236)))));
            end
          for (forvar2282 = (1'h0); (forvar2282 < (2'h2)); forvar2282 = (forvar2282 + (1'h1)))
            begin
              reg2283 = (^reg1999);
              reg2284 <= $unsigned(reg2198);
              reg2285 <= ((reg1861 >= reg2057[(3'h5):(2'h3)]) > (~^$unsigned(reg2135[(4'hc):(3'h7)])));
              reg2286 <= reg1915[(2'h3):(1'h0)];
              reg2287 <= reg2277;
              reg2288 = ($signed(($unsigned((~|reg2213)) ?
                  reg1794 : (~^(reg1843 ?
                      reg2264 : (8'hb3))))) && $signed({$unsigned((wire1765 - reg2233)),
                  ($unsigned(reg2234) ? $unsigned(wire2207) : $signed(reg2091)),
                  (-$signed(reg2016))}));
              reg2289 <= ((((&$signed((8'haa))) ?
                      reg2153[(1'h0):(1'h0)] : (reg2007 - (+(8'ha0)))) ?
                  {(~&$signed(wire1896)),
                      reg1853[(3'h4):(2'h3)],
                      reg2279} : {$signed({(7'h49),
                          reg2056})}) >> ((~|reg1912[(4'hb):(3'h6)]) != (reg1966[(5'h16):(4'hd)] ?
                  ((reg1860 >> (8'hbe)) && reg2111[(1'h0):(1'h0)]) : $unsigned((reg2275 ?
                      reg2245 : reg2124)))));
            end
          reg2290 = ((~^(($unsigned((8'hbf)) || ((7'h51) & reg1950)) + $signed({reg2065}))) ?
              reg1771[(3'h5):(3'h5)] : reg1885[(4'hd):(3'h6)]);
          if (($signed((($signed(reg2241) ?
              {reg1782} : (reg2054 - (8'hbb))) >> (^(~reg1999)))) | (reg2168[(3'h4):(3'h4)] ?
              reg1860 : {$unsigned($signed(reg1950)), reg2175})))
            begin
              reg2291 = (reg2219 ?
                  reg1769[(2'h2):(1'h1)] : ($signed($unsigned($signed(reg2258))) >>> reg1814[(4'hd):(4'h8)]));
              reg2292 = reg1966[(5'h13):(5'h11)];
              reg2293 <= (^~reg2117);
              reg2294 = (~&reg2000[(5'h12):(3'h7)]);
              reg2295 <= reg2117;
              reg2296 = ({$signed(reg2078),
                  $signed($unsigned((wire2207 & reg2171))),
                  ((reg1799[(5'h17):(4'hf)] ? (^reg1978) : (~|(8'ha0))) ?
                      reg2004[(1'h1):(1'h1)] : reg2248)} || reg2028[(5'h10):(4'hc)]);
            end
          else
            begin
              reg2291 = (reg1838 + reg1858);
              reg2293 <= (^~(($signed({(7'h42),
                      (7'h4c)}) == $unsigned(reg2247)) ?
                  reg2250[(5'h1b):(4'he)] : (~$signed({reg1824,
                      reg2109,
                      (8'ha9)}))));
              reg2294 = (~reg2238);
              reg2295 <= (!{((~|(reg2111 ? (8'ha7) : reg2114)) ?
                      (~&reg2247) : (reg2062 > $signed(reg2177))),
                  reg2001[(1'h1):(1'h1)]});
              reg2297 <= (~&$unsigned(((^~(!reg2251)) ?
                  $unsigned((~|forvar2254)) : ((^reg2236) ~^ {reg1774}))));
              reg2298 = {$signed(($unsigned((reg1858 ?
                      reg2242 : reg2276)) != $unsigned($signed(reg1818))))};
            end
        end
      reg2299 <= (^($unsigned(((reg2216 ? reg2177 : reg2149) ?
              (8'hb2) : reg2259[(3'h7):(1'h0)])) ?
          ($signed((8'hb5)) <<< reg2091) : $signed(reg2284[(4'he):(2'h2)])));
      for (forvar2300 = (1'h0); (forvar2300 < (3'h5)); forvar2300 = (forvar2300 + (1'h1)))
        begin
          reg2301 <= (($signed(reg1819[(4'hd):(3'h5)]) ^~ ($signed((reg2299 == (8'ha4))) <<< reg2115[(4'hb):(3'h4)])) + $signed($signed(reg2281[(5'h11):(3'h6)])));
          reg2302 <= reg2250;
          for (forvar2303 = (1'h0); (forvar2303 < (3'h5)); forvar2303 = (forvar2303 + (1'h1)))
            begin
              reg2304 <= $unsigned((~$unsigned($unsigned((forvar2223 && (8'h9c))))));
            end
        end
      if (reg1917)
        begin
          if (({(($unsigned(reg2047) < reg2287) ?
                  (reg2265[(2'h2):(2'h2)] ?
                      $unsigned(reg2098) : $unsigned((7'h41))) : reg2018),
              $unsigned(reg2014)} || ($unsigned(((reg2267 ?
                  reg1987 : (8'ha4)) > $unsigned(reg2021))) ?
              (reg2292 ?
                  $unsigned((^reg1847)) : ($signed(reg2302) ?
                      (reg2180 ? reg2224 : reg2267) : (reg2226 ?
                          reg2215 : reg2066))) : (reg2196 >>> (((7'h51) > reg1822) ?
                  $signed(reg2262) : reg2237)))))
            begin
              reg2305 <= {(^~$unsigned((^{reg2131, reg2018})))};
              reg2306 = (reg2049 <= reg2216[(2'h3):(2'h2)]);
            end
          else
            begin
              reg2306 = reg2060[(5'h11):(3'h7)];
              reg2307 <= (reg2048 ?
                  (($signed($signed(reg2078)) >>> reg2151[(1'h0):(1'h0)]) ?
                      $signed(((reg1936 ? reg1788 : (7'h4a)) >= (reg2242 ?
                          (7'h4b) : reg1967))) : ((~^$signed(reg2210)) ?
                          (8'ha8) : ((reg2027 | reg2217) < (~&reg2278)))) : $signed((7'h43)));
            end
          reg2308 <= (!$unsigned(reg1875[(3'h6):(2'h3)]));
          for (forvar2309 = (1'h0); (forvar2309 < (1'h0)); forvar2309 = (forvar2309 + (1'h1)))
            begin
              reg2310 = ((((+$signed(reg2229)) <= reg2217[(4'ha):(1'h0)]) ?
                  $signed($unsigned((reg2236 ?
                      reg2056 : reg1928))) : (((reg1956 ?
                          forvar2223 : (8'ha1)) ?
                      (reg2257 ?
                          reg2299 : wire1765) : $unsigned(reg2042)) <<< reg2109)) && reg2187);
              reg2311 <= reg2219[(3'h7):(3'h7)];
              reg2312 = $signed({(8'ha5),
                  (reg2053 ?
                      (~^{reg2066,
                          reg2064,
                          reg2269}) : ($unsigned(reg2021) && $signed((8'hab))))});
              reg2313 = {{$signed($signed(reg2078)), reg1803},
                  (~|{({wire2207, (7'h56), reg1788} ^ (reg2142 ?
                          reg2030 : reg2015)),
                      (7'h4e),
                      reg1775}),
                  ((&($signed(reg2242) ?
                      $unsigned((8'hba)) : {reg1942})) ^~ (($unsigned((7'h53)) ^ (|(8'ha1))) ?
                      ($signed(forvar2260) <= $signed(reg2222)) : ((reg2276 && reg2217) ?
                          $signed(reg2258) : reg2297)))};
              reg2314 = (!(reg2135 >= reg1912[(4'hb):(4'h8)]));
            end
          reg2315 = (reg2131 ?
              (({$signed(reg1799)} != ((reg2091 ?
                  reg1981 : reg2219) + (wire1762 <= reg1928))) - forvar2274) : $signed((reg2258[(4'h8):(3'h7)] ?
                  $signed($unsigned(reg2114)) : reg2028[(4'hb):(1'h1)])));
          reg2316 <= $unsigned(((~|reg1936[(4'he):(4'hc)]) >>> (~&((+(8'ha4)) ?
              reg2136 : ((8'ha2) ? reg2272 : reg2028)))));
          for (forvar2317 = (1'h0); (forvar2317 < (1'h1)); forvar2317 = (forvar2317 + (1'h1)))
            begin
              reg2318 <= ((reg2298[(4'h8):(3'h5)] ?
                  $signed({$unsigned(reg2088)}) : (^~reg2021[(1'h1):(1'h0)])) >= reg2066);
              reg2319 = $signed((reg1790[(3'h6):(3'h6)] ?
                  (reg1803[(1'h1):(1'h0)] != ($signed(reg1777) ?
                      {reg1808} : reg2225)) : $signed($signed((&reg2233)))));
            end
        end
      else
        begin
          if ((~^$signed($unsigned($unsigned((reg2116 * reg2002))))))
            begin
              reg2305 <= $unsigned($signed({$signed($signed(reg1848))}));
              reg2306 = reg1991[(5'h11):(4'h9)];
              reg2309 = (($unsigned(($signed(reg2259) ^ (~|reg2310))) ?
                      (((|(7'h4e)) ?
                          (reg2107 ~^ reg2265) : {reg1973,
                              reg2108}) && ($signed(reg2150) ?
                          reg2132[(2'h2):(2'h2)] : {reg2171,
                              reg1962})) : $signed(reg2233[(1'h0):(1'h0)])) ?
                  reg2210[(4'hb):(3'h6)] : reg1840[(3'h7):(3'h4)]);
              reg2311 <= ((($signed((reg1811 ?
                          reg1832 : reg2149)) >> wire2043) ?
                      $unsigned((reg1880 || {reg1978,
                          (7'h4e),
                          (8'hbc)})) : reg2067[(2'h2):(1'h0)]) ?
                  $unsigned((($unsigned(reg2258) == $unsigned(reg1814)) ?
                      ($signed(forvar2209) | (reg2093 ?
                          reg1838 : reg2049)) : (8'hab))) : (reg2307 != ($unsigned((8'h9d)) ?
                      {reg2310[(4'h8):(1'h1)],
                          reg1791,
                          reg1991} : {reg2219[(3'h6):(1'h1)],
                          (reg1791 ? reg1868 : reg1796)})));
              reg2312 = reg2028;
            end
          else
            begin
              reg2305 <= reg2198;
              reg2306 = ($signed((~&(|reg2054))) ?
                  ((-$unsigned({reg1967,
                      reg2028})) - ($signed((reg2116 && reg1775)) - $signed((8'hb1)))) : $signed(reg2270[(2'h2):(2'h2)]));
              reg2307 <= $signed({(((reg2114 ? (8'ha0) : reg2293) ?
                      {(7'h42), reg1804, forvar2254} : (reg1923 ?
                          (8'hba) : (7'h50))) + reg2213)});
              reg2309 = reg2292;
            end
          reg2316 <= (forvar2274 >>> $signed($unsigned(((reg1768 ?
              forvar2317 : reg1788) == (|reg1814)))));
          reg2317 = ($unsigned($unsigned($signed((reg2054 < forvar2260)))) ?
              (^~$signed(reg1857[(4'h8):(3'h6)])) : reg2175[(1'h1):(1'h1)]);
          if ({(reg2218 ?
                  ((-(^reg2001)) ?
                      {(reg2023 != reg1977)} : {(forvar2309 ?
                              reg2264 : reg2311)}) : (^~(reg2021[(3'h5):(2'h2)] ?
                      $signed((8'h9c)) : $unsigned(reg1936))))})
            begin
              reg2318 <= $signed((reg1932[(4'hb):(2'h3)] && (reg1782 ?
                  reg2264[(1'h1):(1'h0)] : ((reg2131 ~^ reg2294) ?
                      (reg2021 ? reg1911 : wire1764) : (reg2198 * reg2111)))));
              reg2319 = $unsigned((|$unsigned(((+reg2056) ?
                  reg2243 : (reg2293 < reg2151)))));
              reg2320 <= $unsigned($signed((((reg2097 ? reg1893 : wire2043) ?
                  $signed(reg1783) : (~reg1893)) * ((reg2248 ?
                      (7'h43) : reg2286) ?
                  $unsigned(reg2056) : (reg1973 ? (7'h4e) : reg1794)))));
              reg2321 <= (-(-(^~reg2063[(1'h1):(1'h0)])));
              reg2322 <= {wire1763[(2'h2):(2'h2)]};
              reg2323 = $signed($signed({reg2196[(3'h6):(2'h3)],
                  $signed(reg2258[(3'h5):(3'h4)])}));
              reg2324 <= reg2220;
            end
          else
            begin
              reg2319 = (-((($signed(reg1857) ? (~^reg2316) : {reg2243}) ?
                      (reg2224 >>> (^~reg2109)) : reg2053) ?
                  (~&reg1796) : {reg2187[(3'h5):(1'h1)]}));
              reg2320 <= reg1846;
            end
        end
    end
  always
    @(posedge clk) begin
      if (({(|{$signed(wire1760), reg1973, $signed(reg1853)})} * reg2071))
        begin
          reg2325 <= ($unsigned(reg2149) ?
              {reg2097,
                  (|$signed({reg2010})),
                  (+(~^(~&reg2048)))} : ({$signed({reg2311})} <= (~reg1902)));
          if ((reg2262[(3'h7):(3'h6)] > $signed(reg2000)))
            begin
              reg2326 = $signed({reg2131,
                  $signed({reg2175[(4'hb):(4'hb)],
                      (reg1926 && reg1950),
                      $unsigned(reg1861)})});
              reg2327 = ($signed(($signed(reg2029) ?
                      ((reg2289 ?
                          reg2047 : (8'hb9)) <= (-reg2238)) : ($unsigned(reg2321) ?
                          (reg1990 != wire1762) : reg2220))) ?
                  reg1782 : $unsigned(reg2067));
              reg2328 = (~(~&(-reg1998)));
              reg2329 <= (&$unsigned(reg2284[(5'h13):(4'h8)]));
            end
          else
            begin
              reg2326 = (!$unsigned(reg2194[(2'h3):(1'h1)]));
              reg2329 <= reg1967[(1'h1):(1'h0)];
            end
        end
      else
        begin
          if ($signed(((reg1995 ?
              (~^reg1923) : $signed(((7'h54) ^ reg1891))) - $signed(reg2264))))
            begin
              reg2326 = ((&(((|reg2187) ?
                      reg2326[(3'h6):(2'h3)] : reg1998[(4'he):(3'h7)]) ?
                  ((reg2067 && reg2027) ?
                      $signed(reg2165) : reg2263) : $signed(reg2214))) >= ((8'h9d) ^~ ($unsigned(wire1764) ?
                  (-(~^reg2143)) : reg1814)));
              reg2327 = reg2116;
              reg2328 = $unsigned((-(((|reg2149) || (reg2039 ~^ reg2143)) ?
                  ((~&reg2082) ?
                      reg1869 : $unsigned(reg1832)) : $signed((reg2065 ?
                      reg1987 : reg1774)))));
            end
          else
            begin
              reg2326 = $unsigned(((!{$signed(reg2262)}) || reg1788[(2'h3):(2'h2)]));
            end
          reg2330 = ((8'h9e) < ($signed(reg1855[(3'h4):(1'h1)]) * $signed(reg1917[(3'h5):(3'h5)])));
          for (forvar2331 = (1'h0); (forvar2331 < (1'h1)); forvar2331 = (forvar2331 + (1'h1)))
            begin
              reg2332 <= ((reg2271[(3'h5):(1'h0)] * ((&reg1829[(4'h8):(3'h7)]) > $signed((&reg2255)))) ?
                  reg1796[(1'h0):(1'h0)] : $unsigned($signed(reg1790[(3'h7):(2'h3)])));
              reg2333 <= reg2002[(2'h3):(2'h3)];
              reg2334 <= $unsigned($signed({$unsigned(((8'hbc) > (8'ha4)))}));
              reg2335 <= $signed(reg1940);
              reg2336 <= reg1893[(3'h7):(3'h5)];
            end
          for (forvar2337 = (1'h0); (forvar2337 < (3'h5)); forvar2337 = (forvar2337 + (1'h1)))
            begin
              reg2338 = (-reg2161);
              reg2339 = $unsigned((reg1993[(5'h11):(4'he)] << $signed($unsigned($signed(reg1860)))));
              reg2340 <= ((^~($unsigned((~&reg1768)) | $signed(reg1771))) + reg1991);
              reg2341 <= {(reg1891[(3'h4):(1'h0)] < $signed(((reg1990 ?
                      reg2318 : reg2221) ^ reg2244[(3'h5):(3'h4)])))};
              reg2342 <= (reg2136[(1'h0):(1'h0)] <= ($unsigned($unsigned((7'h50))) <<< (~$unsigned((reg2067 + (7'h48))))));
            end
          for (forvar2343 = (1'h0); (forvar2343 < (2'h2)); forvar2343 = (forvar2343 + (1'h1)))
            begin
              reg2344 <= $unsigned({$unsigned($signed((reg2054 & reg2053))),
                  $signed($signed((!reg2143)))});
              reg2345 = reg1861[(1'h1):(1'h1)];
              reg2346 = $signed((~(+($signed(reg2279) ?
                  forvar2337[(1'h0):(1'h0)] : $unsigned(reg1833)))));
              reg2347 = {(((+$signed(reg2017)) + ($unsigned(reg2071) ?
                          (reg2067 ? reg2265 : reg1978) : reg2054)) ?
                      $unsigned(((^~(8'ha1)) ^ (reg1932 ?
                          (7'h42) : reg1905))) : reg2029)};
              reg2348 = $signed((8'hbb));
            end
          for (forvar2349 = (1'h0); (forvar2349 < (3'h5)); forvar2349 = (forvar2349 + (1'h1)))
            begin
              reg2350 = ($signed($signed(reg1769[(1'h1):(1'h1)])) ?
                  $unsigned($signed(((reg1797 ?
                      reg2286 : (8'hba)) | reg2109[(3'h4):(1'h0)]))) : (wire1762 ?
                      $unsigned(reg1843) : (!(-(!reg2047)))));
            end
          if ((~|$unsigned(reg2333)))
            begin
              reg2351 <= reg1771;
            end
          else
            begin
              reg2352 = $unsigned(reg2268);
            end
        end
      reg2353 = $unsigned(((((reg1826 ^ reg1785) & (reg2063 ~^ reg1808)) <<< ($unsigned((7'h40)) ^~ (wire1761 & reg2215))) > reg2114[(3'h7):(3'h7)]));
      reg2354 = $unsigned(((^~$signed($signed(reg2104))) ?
          (+(8'hb5)) : (^reg2334)));
      if ((reg2078 | ($unsigned(((-reg2009) ?
          (&reg1794) : {reg2241})) >>> reg1885)))
        begin
          reg2355 <= reg2243[(1'h0):(1'h0)];
          if (reg2064)
            begin
              reg2356 <= $signed(reg1911);
              reg2357 = reg2243;
              reg2358 = {((+((|reg2006) ~^ (reg1990 ?
                      reg1908 : reg1897))) - ($unsigned(((8'hb0) < reg2110)) < (+$signed(reg1877)))),
                  reg2262[(2'h2):(1'h1)]};
              reg2359 <= $signed((reg2307[(3'h4):(2'h2)] ?
                  ((reg2037[(3'h6):(3'h4)] <<< (reg2064 && reg1838)) ?
                      reg1768[(2'h3):(2'h3)] : reg1932) : reg2094));
              reg2360 <= $signed(reg1936);
            end
          else
            begin
              reg2357 = reg1993[(3'h7):(1'h0)];
              reg2359 <= (reg2224[(2'h3):(2'h3)] ?
                  reg2116[(1'h0):(1'h0)] : (reg2048 ?
                      ({(~^reg2226)} ? reg2271 : wire1764) : (&(|(reg2346 ?
                          reg2299 : reg1808)))));
              reg2361 = $signed((&$signed(($signed(reg2131) ?
                  (reg2244 && (8'ha2)) : $signed(reg2062)))));
              reg2362 = (|$signed((~|$unsigned($unsigned(reg1769)))));
              reg2363 <= ($unsigned((^{reg1848,
                      (reg1768 ? reg2111 : (8'haf))})) ?
                  (-reg2143) : ((~((|reg2094) ?
                          {reg1880} : ((8'hbc) ? reg1900 : reg2241))) ?
                      ((~&$unsigned(reg2334)) != (|$signed(reg1847))) : reg2171[(4'hc):(3'h7)]));
              reg2364 = $signed((|(7'h48)));
            end
          for (forvar2365 = (1'h0); (forvar2365 < (1'h0)); forvar2365 = (forvar2365 + (1'h1)))
            begin
              reg2366 = {($unsigned(((~^reg2075) ?
                      (^reg2220) : (reg2004 >>> reg2305))) > reg1912)};
              reg2367 = reg2352[(4'h9):(3'h6)];
              reg2368 <= (~^(~|(!reg1853[(1'h0):(1'h0)])));
              reg2369 = $unsigned({$signed((7'h4c)),
                  $unsigned(reg1942[(2'h2):(2'h2)])});
            end
          for (forvar2370 = (1'h0); (forvar2370 < (3'h6)); forvar2370 = (forvar2370 + (1'h1)))
            begin
              reg2371 = reg2171;
              reg2372 = reg2351[(4'he):(4'ha)];
              reg2373 = (+((reg2095[(1'h0):(1'h0)] <= (7'h4c)) ?
                  reg1811[(1'h1):(1'h1)] : $unsigned(($signed(reg1956) | reg1962))));
              reg2374 = $unsigned(reg1884);
              reg2375 = (-(!$signed((+$signed(reg1991)))));
              reg2376 <= reg2057;
            end
          for (forvar2377 = (1'h0); (forvar2377 < (2'h2)); forvar2377 = (forvar2377 + (1'h1)))
            begin
              reg2378 = reg1843;
            end
          for (forvar2379 = (1'h0); (forvar2379 < (2'h2)); forvar2379 = (forvar2379 + (1'h1)))
            begin
              reg2380 <= ((&(^(^~reg1961[(5'h10):(1'h0)]))) * {reg1839[(4'hd):(2'h2)]});
            end
          reg2381 = {{($signed(reg2258) ?
                      $unsigned({reg1998, reg2060, reg1826}) : reg2344),
                  reg1915}};
        end
      else
        begin
          for (forvar2355 = (1'h0); (forvar2355 < (1'h1)); forvar2355 = (forvar2355 + (1'h1)))
            begin
              reg2356 <= $signed({reg2056});
              reg2359 <= reg1940;
              reg2360 <= $unsigned((($signed($unsigned(forvar2379)) | (reg1883[(5'h16):(4'h9)] >>> (^~reg1814))) * $signed(reg2353)));
              reg2361 = (^reg2108);
            end
          for (forvar2362 = (1'h0); (forvar2362 < (3'h6)); forvar2362 = (forvar2362 + (1'h1)))
            begin
              reg2364 = $signed(reg2244[(2'h3):(2'h3)]);
              reg2365 = (|reg1847);
              reg2368 <= reg2333[(2'h3):(2'h3)];
              reg2370 <= (($signed(reg1838) ?
                  {{reg2301},
                      (+$unsigned(reg1892))} : reg2234[(4'hd):(4'hb)]) & {$signed(reg2347[(4'h9):(3'h7)]),
                  ({(&reg2262), (reg1869 ? reg2218 : reg2093)} ?
                      {(reg2341 ? reg1893 : reg2067)} : ($signed(reg2243) ?
                          reg2038 : (~|reg2255)))});
            end
          reg2376 <= $unsigned((7'h43));
        end
      if (((reg2336 ?
              (reg2308 ?
                  (^wire1762) : ((reg2007 * reg2114) + (reg1883 <= (7'h40)))) : $signed((~|(reg2218 ?
                  reg1782 : reg1911)))) ?
          reg2234[(4'hb):(4'ha)] : ((^~reg2347[(4'hb):(3'h5)]) ?
              reg1892[(4'ha):(4'h9)] : reg1961)))
        begin
          reg2382 = reg2372[(4'ha):(1'h0)];
          for (forvar2383 = (1'h0); (forvar2383 < (3'h6)); forvar2383 = (forvar2383 + (1'h1)))
            begin
              reg2384 <= $signed((8'ha7));
              reg2385 <= $unsigned($unsigned(reg2143));
              reg2386 = $unsigned((reg2196 ?
                  $signed(((-forvar2331) + (&reg1911))) : reg1926));
              reg2387 = reg1906;
              reg2388 <= (7'h52);
              reg2389 = reg2372[(5'h12):(3'h7)];
              reg2390 <= {(~^(|reg2271[(3'h4):(1'h0)])), reg2160};
            end
          reg2391 <= (~&$signed(($signed(reg2389[(3'h5):(3'h5)]) ?
              $unsigned($unsigned(reg2255)) : $unsigned((reg1923 * reg2329)))));
          reg2392 = ($signed(((!(reg2380 ? reg2252 : reg2114)) ?
                  reg1902[(4'h8):(3'h4)] : (~^(reg2330 - reg1880)))) ?
              $signed(((reg1833 >> $signed((7'h41))) * $signed(reg1961))) : (($unsigned($signed(forvar2331)) && ((^reg2082) ?
                  $unsigned(reg1923) : reg1948)) && (~|((-(7'h4b)) ?
                  reg2088[(5'h14):(5'h12)] : $signed(reg1883)))));
          reg2393 <= ({($signed((reg2352 | reg2231)) ?
                  ((~^reg2250) ?
                      (reg2042 * (8'hb8)) : $signed((8'hb3))) : reg1806[(4'h9):(4'h8)]),
              $signed(((~reg2370) ?
                  (reg2333 - (8'hb2)) : (reg2357 ?
                      (7'h4a) : (8'hbf))))} ~^ reg1875[(3'h4):(1'h1)]);
          for (forvar2394 = (1'h0); (forvar2394 < (2'h2)); forvar2394 = (forvar2394 + (1'h1)))
            begin
              reg2395 <= (|(+(((|reg2116) + (reg1847 ^ (8'h9f))) ?
                  reg1843[(3'h7):(2'h3)] : $unsigned((reg2161 ?
                      (7'h56) : reg2029)))));
              reg2396 <= {$unsigned({((~reg2063) > {reg2149, reg1839, reg2176}),
                      $signed(reg1877),
                      reg2165})};
              reg2397 = reg2264[(5'h12):(4'he)];
            end
          if ({($signed(reg2358[(2'h2):(1'h1)]) ?
                  (7'h41) : ((~&(reg1912 ?
                      reg1966 : reg1861)) + (((7'h42) && (8'hb4)) != (&reg2046)))),
              $signed((($signed(reg1829) * $unsigned(reg2363)) && $unsigned((reg2229 ?
                  (8'hbd) : reg2075)))),
              (reg2210 ?
                  {reg2046,
                      (reg2042 >> (reg1948 ^ reg2093))} : reg2243[(1'h0):(1'h0)])})
            begin
              reg2398 = (reg2234 ? (~|reg2017) : reg2169[(1'h0):(1'h0)]);
              reg2399 = {$unsigned(($unsigned(reg2384[(2'h3):(2'h3)]) ^ ($signed(reg2385) <<< reg2308[(3'h5):(2'h3)]))),
                  $unsigned($unsigned(($signed((8'ha0)) ?
                      reg2287 : $unsigned((8'hac))))),
                  $signed($signed(reg2151))};
              reg2400 <= $signed(($signed({$signed(reg2223),
                  $signed(reg1843)}) ^~ $unsigned(((reg2396 * reg2018) >>> (reg2007 ~^ reg1803)))));
              reg2401 <= (+$unsigned((~&(&(!reg2396)))));
            end
          else
            begin
              reg2398 = (-{$unsigned(reg2388[(3'h5):(1'h1)])});
              reg2400 <= reg2301[(1'h1):(1'h0)];
              reg2402 = $signed((($signed({reg2224, reg2330, (8'hb3)}) ?
                  reg2176 : ((+forvar2383) <= $unsigned(reg1796))) >>> $signed($signed($unsigned(reg1840)))));
            end
        end
      else
        begin
          if ($signed($unsigned({((reg2115 ? reg2378 : reg2114) ?
                  (reg2057 >= reg1885) : $signed(reg1940))})))
            begin
              reg2383 <= (({$unsigned($signed((8'hba))),
                      $unsigned(reg1771),
                      $unsigned((reg1826 <<< reg2378))} ?
                  reg2098[(5'h11):(4'h8)] : reg2375) < (reg2000[(3'h6):(3'h5)] ?
                  (reg2071 ?
                      ($unsigned(reg2234) << {reg2265}) : (~&{reg2136})) : $signed((~((8'hb8) ?
                      reg2369 : reg1791)))));
              reg2384 <= reg2332;
              reg2385 <= (reg1906 ?
                  (8'had) : ((reg1833 ?
                      $unsigned(reg2371[(1'h0):(1'h0)]) : $unsigned($unsigned((7'h41)))) >> (~&(~^(reg2355 != reg2264)))));
              reg2386 = $unsigned((($signed((reg2121 ?
                      reg2165 : reg2321)) << (+{reg1836, reg1768, (8'ha3)})) ?
                  reg2382[(4'h9):(3'h6)] : (reg2356 >> ((reg2318 ?
                      reg2161 : reg2308) & {(7'h40), (8'hab), reg1846}))));
              reg2388 <= reg2110[(5'h15):(5'h15)];
              reg2390 <= reg2028[(5'h13):(4'hf)];
              reg2392 = {((reg2063[(2'h2):(2'h2)] ?
                          {((8'hbe) && reg2002),
                              {reg2302,
                                  reg1956,
                                  reg2142}} : $unsigned(reg1839)) ?
                      (reg1966 ?
                          reg1853 : ($unsigned((8'ha2)) ?
                              $unsigned(reg2365) : reg2115[(4'ha):(1'h0)])) : $unsigned((~|(|reg1861))))};
            end
          else
            begin
              reg2382 = reg2365;
              reg2386 = $unsigned(((reg2335[(4'hd):(2'h3)] - (~&reg1785)) >>> reg2047));
              reg2388 <= reg2380[(4'h8):(3'h6)];
              reg2389 = $signed({reg2078,
                  ((^(reg2214 - reg2104)) ?
                      $signed($unsigned(reg1839)) : reg2151)});
            end
          reg2394 = ($unsigned(reg2385[(4'h8):(3'h7)]) ?
              $unsigned(reg2355[(3'h6):(1'h0)]) : (($unsigned((reg2229 ^ reg2330)) ?
                  (-reg2116) : ($unsigned(reg1885) ?
                      (reg2255 ^~ reg1791) : $unsigned(reg2297))) <<< (7'h55)));
          reg2395 <= ($signed($signed((^{reg1828}))) ?
              $unsigned((&(reg2389 <= reg2117))) : reg2132[(1'h0):(1'h0)]);
          if (((^~$signed((!reg2271))) ?
              (+reg1803) : ((~|({(7'h56), (8'hb9)} ?
                      (reg2275 >> reg2195) : reg2165)) ?
                  $signed(reg2302[(2'h3):(1'h0)]) : ($unsigned($unsigned((8'hb9))) ?
                      $signed((7'h48)) : reg2275))))
            begin
              reg2397 = (reg2284[(4'hb):(4'hb)] || $signed($signed($unsigned($unsigned((8'haf))))));
              reg2398 = (|((reg2338[(1'h1):(1'h0)] ?
                      ((^reg1979) ?
                          $signed(reg2390) : reg1832) : $unsigned(reg1973)) ?
                  ($unsigned(reg1892) ?
                      (reg2252[(3'h4):(2'h3)] * reg2354[(3'h4):(2'h3)]) : (~reg1848)) : reg2327));
              reg2400 <= ((reg2260 | ($unsigned((|reg2021)) ^~ $unsigned((reg1978 ?
                      (8'ha9) : forvar2355)))) ?
                  $signed(reg2342[(3'h5):(1'h0)]) : (^~((^(8'hbd)) <= reg1981)));
            end
          else
            begin
              reg2396 <= ($unsigned((8'ha0)) ?
                  ((8'ha3) ?
                      reg2380 : $signed($signed((reg1915 ?
                          (7'h47) : reg2046)))) : $signed((({(7'h52)} ?
                      (&(7'h47)) : (forvar2370 > (8'ha6))) || (^~(reg2373 ^ reg2262)))));
            end
          if (($unsigned(reg1999) > (wire2207 == ($signed(reg2368[(4'ha):(2'h3)]) ?
              $signed($unsigned(reg2329)) : reg2344[(4'h9):(1'h1)]))))
            begin
              reg2401 <= reg2329[(2'h3):(1'h0)];
              reg2403 <= ((reg2307 ?
                  reg2390 : ($unsigned($signed(reg2395)) ?
                      $unsigned((reg2347 ?
                          reg2107 : (8'hab))) : $unsigned(reg2002))) - $signed((reg2322 ?
                  ($signed(reg1911) ^ (^(7'h4e))) : (-$signed(reg1904)))));
              reg2404 <= (forvar2394[(5'h13):(4'ha)] != (-((~&$signed(reg1973)) ?
                  (~$unsigned(reg2360)) : (!(reg1928 | reg2341)))));
              reg2405 = (forvar2377[(3'h6):(3'h5)] ?
                  $signed((~$unsigned(reg2260[(4'hb):(3'h6)]))) : reg1897[(5'h1b):(4'hf)]);
              reg2406 = (&$unsigned($unsigned($unsigned($unsigned(reg2388)))));
              reg2407 <= $unsigned($unsigned((~|$unsigned($signed(reg2152)))));
              reg2408 <= (({reg2217[(3'h6):(3'h6)],
                  (8'hb5),
                  reg2001} < $unsigned(($unsigned((8'h9e)) <<< reg2187))) <<< ({((reg2004 ?
                              (8'hba) : reg2395) ?
                          (reg1846 + (7'h4c)) : {reg2327})} ?
                  ((reg2244[(3'h6):(1'h1)] ?
                      $unsigned((8'ha5)) : ((8'hbf) ?
                          reg2374 : reg2006)) || $unsigned((reg1977 ?
                      reg2200 : reg2342))) : $signed(((|reg1788) <= reg1991))));
            end
          else
            begin
              reg2402 = (reg1824[(4'ha):(4'h9)] == reg2215[(4'he):(2'h2)]);
              reg2403 <= reg2198;
              reg2404 <= reg1891;
              reg2405 = ({((8'hae) ?
                          reg1982[(5'h11):(3'h4)] : ($unsigned(reg2097) & {reg1869,
                              (8'hb0)}))} ?
                  (|$signed(((reg1811 ~^ (8'ha5)) < reg2143[(3'h5):(1'h0)]))) : (~&(reg2387[(4'he):(3'h7)] == reg2260)));
              reg2406 = (reg1966[(4'hd):(2'h3)] >>> reg2094[(1'h0):(1'h0)]);
            end
        end
      reg2409 <= $signed((reg2114 != reg2369[(5'h10):(1'h0)]));
      reg2410 <= $signed((&{(-reg2062[(3'h5):(2'h2)])}));
    end
  always
    @(posedge clk) begin
      for (forvar2411 = (1'h0); (forvar2411 < (1'h1)); forvar2411 = (forvar2411 + (1'h1)))
        begin
          if (wire1761)
            begin
              reg2412 = $unsigned(($unsigned($unsigned((-reg1788))) + (((reg2271 ?
                          reg1905 : reg2095) ?
                      ((8'hb6) ^ reg2149) : (~reg2223)) ?
                  {(reg2297 ? reg1828 : reg2248)} : ($signed(reg1855) ?
                      reg2270 : reg2075))));
              reg2413 <= ($signed(reg2066[(2'h2):(2'h2)]) && (($unsigned(reg1853[(3'h4):(1'h1)]) <= reg2360[(5'h10):(4'hf)]) ?
                  reg2066 : ($unsigned($signed(reg2263)) * $signed($unsigned(reg1819)))));
              reg2414 <= $unsigned(($signed((~{reg2242,
                  (7'h55),
                  reg1800})) < ((|$unsigned(reg2329)) << $signed(reg2409))));
            end
          else
            begin
              reg2413 <= (7'h57);
              reg2414 <= (~^$unsigned(($signed((~&reg2388)) ?
                  ($unsigned(reg2078) ?
                      (!reg1880) : $unsigned(reg2168)) : (^reg2037))));
              reg2415 = ($signed({$signed($unsigned(reg2175))}) ?
                  reg2244[(3'h5):(1'h1)] : $unsigned(($unsigned($signed(reg2047)) ?
                      $unsigned(reg2108[(2'h3):(1'h0)]) : (~&(7'h4c)))));
            end
          reg2416 = ($signed((($signed(reg1962) ?
                  reg1904[(2'h2):(1'h0)] : reg1993) || {(reg2176 ?
                      reg2221 : reg1940),
                  (reg1885 <= reg2054)})) ?
              {(((reg1814 ? reg2287 : reg2098) - (^reg1987)) + (7'h57)),
                  {reg2002[(2'h2):(1'h1)], {((8'ha5) >> reg2388)}},
                  (reg1771 ?
                      ($signed(reg2214) ?
                          (reg2070 | reg1977) : ((7'h55) ?
                              (7'h52) : (7'h4c))) : {(reg1804 || reg2070)})} : reg1861);
          reg2417 <= (&reg1911[(4'hf):(4'ha)]);
          if ((({((reg1956 & reg2311) ? (~^reg1904) : $signed(reg1774)),
                  $unsigned(reg2260)} >> ((reg2318 >> (reg2226 && reg1788)) ?
                  (~|{(8'hb6), reg2160}) : ((reg2048 * (7'h4b)) ?
                      {reg2316, reg1858, reg1828} : {reg1774, reg2039}))) ?
              $signed((8'hab)) : $signed((^$signed($unsigned((8'hbe)))))))
            begin
              reg2418 <= reg1999[(5'h15):(3'h7)];
              reg2419 = ($signed({reg2415}) ?
                  (^$unsigned(forvar2411[(2'h3):(2'h2)])) : {{$unsigned((reg2223 - reg2217)),
                          (!$signed(reg1839)),
                          ($signed(reg2218) >= reg1869)}});
              reg2420 <= reg2029[(5'h15):(4'hb)];
            end
          else
            begin
              reg2419 = $signed(reg2108[(4'hf):(2'h2)]);
              reg2421 = $signed(reg2171[(4'h8):(3'h7)]);
              reg2422 <= ((7'h41) & reg2332);
            end
          reg2423 = reg1891[(4'hd):(4'h9)];
          for (forvar2424 = (1'h0); (forvar2424 < (3'h4)); forvar2424 = (forvar2424 + (1'h1)))
            begin
              reg2425 = $signed(reg2255);
              reg2426 = {(~$unsigned((reg2255[(2'h2):(1'h1)] <<< (reg2195 ^~ reg2097)))),
                  reg2423,
                  $signed((+$unsigned(reg2175)))};
            end
          reg2427 = ($unsigned($signed(((-reg1771) ?
                  (reg2098 <= reg1991) : reg2056))) ?
              $unsigned({$unsigned((~^reg2264)),
                  reg2351[(4'h8):(3'h7)]}) : $unsigned((((reg2107 >= reg2117) || $unsigned(reg1794)) & {$unsigned((8'haf)),
                  reg2001,
                  (reg2029 ? forvar2411 : reg1832)})));
        end
    end
  always
    @(posedge clk) begin
      if ((!{$signed(reg1940)}))
        begin
          reg2428 = {reg2196[(3'h4):(2'h2)],
              (reg1903 ^~ ($signed((reg2136 ? reg1928 : reg2135)) ?
                  reg2065[(5'h15):(4'hf)] : ((7'h51) ?
                      (reg2038 < reg2067) : $signed(reg1846))))};
          reg2429 = ($unsigned(reg1825[(5'h14):(4'hb)]) ?
              (((8'haa) ?
                  {$unsigned(reg2360),
                      (reg2002 ? wire1764 : reg2363)} : ((wire1760 ?
                      (8'hbd) : reg1806) < reg1811[(2'h3):(1'h0)])) ^ (((reg2152 + reg2187) ?
                      reg2057[(3'h4):(2'h2)] : (reg1771 ? reg1783 : (8'hbd))) ?
                  $signed($unsigned(reg2221)) : ({(8'h9e)} < $unsigned(reg1857)))) : (-($signed({reg2218}) != $signed($unsigned(reg1885)))));
          reg2430 = ($signed({({reg2142, reg1897, reg2021} ?
                      (&(8'hbe)) : ((8'hac) ? (8'hb9) : reg1923)),
                  ($unsigned((8'hb1)) < $unsigned(reg1791))}) ?
              $unsigned({(^~(reg2169 ? reg2248 : reg2116)),
                  ($signed(reg2286) != (reg2305 & reg2062))}) : ($unsigned((~&reg1777[(4'h8):(1'h0)])) - reg2015[(4'h8):(3'h4)]));
          reg2431 = ({reg1987[(4'h9):(1'h0)],
                  $unsigned($signed(reg2038)),
                  (8'hb0)} ?
              reg2383[(4'hf):(1'h1)] : $signed((~(~^(reg1966 < reg1885)))));
          reg2432 = $signed((($signed($unsigned(reg2390)) ^~ ({reg2220} ?
              reg2223 : reg1977)) - (8'hbd)));
        end
      else
        begin
          reg2433 <= $unsigned($unsigned((^{(reg2243 <= reg1816)})));
          reg2434 = ((reg2082 - (((8'hb7) >> (reg1855 ^~ reg2169)) * reg1829)) ?
              (!$signed($signed((reg1825 | reg1782)))) : ($unsigned((&{(7'h4e),
                      (7'h43),
                      reg2082})) ?
                  ($unsigned(reg1877) < ($unsigned(reg2403) ?
                      $signed(reg2226) : (reg2088 << (8'hae)))) : (&reg2165)));
          for (forvar2435 = (1'h0); (forvar2435 < (3'h5)); forvar2435 = (forvar2435 + (1'h1)))
            begin
              reg2436 <= (((({reg1991} || (!reg1950)) ~^ reg2335) ?
                  reg2417 : reg2028[(5'h11):(3'h4)]) << (~{$unsigned(reg1803[(2'h2):(1'h0)])}));
              reg2437 <= (7'h55);
              reg2438 = {({(((8'ha7) < (8'hae)) ?
                              $unsigned(reg2422) : (^~(7'h54))),
                          ($unsigned(wire1765) * (~&reg1819))} ?
                      ($signed((reg2037 ? reg1880 : reg1948)) ?
                          (&(~reg2153)) : (^(reg2351 <<< reg2114))) : ({$unsigned(reg2048),
                          reg2388[(5'h1a):(5'h11)]} ^~ {(reg2356 ?
                              reg2422 : reg2324),
                          wire2208[(1'h0):(1'h0)],
                          reg2262[(3'h6):(1'h0)]})),
                  reg2118};
              reg2439 = reg1832;
            end
          reg2440 <= ((+$signed(reg1926[(4'ha):(3'h6)])) >> reg2161[(4'h8):(1'h1)]);
          if ($signed($unsigned((7'h53))))
            begin
              reg2441 = $unsigned(reg2268);
              reg2442 = (((-{reg2198,
                          $unsigned(reg2428),
                          reg2039[(3'h4):(2'h3)]}) ?
                      ($signed((~^reg2414)) < reg2248[(1'h0):(1'h0)]) : $signed((~^reg2078[(5'h11):(4'he)]))) ?
                  ((reg1985 > ((reg2216 <= reg1791) ?
                          reg2428[(3'h7):(1'h1)] : {reg1978, reg1766})) ?
                      $unsigned(reg2115) : $unsigned(((reg2318 >>> (7'h47)) ?
                          (&reg2279) : (reg1782 ?
                              reg1935 : reg2121)))) : $unsigned(($unsigned(reg1985) ?
                      ({reg1825,
                          reg1936,
                          reg1993} > (~|(7'h4d))) : $signed(reg1915[(3'h4):(3'h4)]))));
              reg2443 = reg1977;
              reg2444 <= $signed((-$signed($signed($unsigned(reg2368)))));
              reg2445 = $signed(((-(((8'haa) != reg2311) ?
                  $signed(reg1788) : (reg2376 > reg1993))) - (^wire1765[(3'h4):(1'h1)])));
            end
          else
            begin
              reg2441 = reg2429;
              reg2444 <= (8'hbb);
              reg2446 <= {reg1796,
                  $unsigned($signed(((wire1763 & (8'had)) && $signed(reg2320))))};
              reg2447 <= (!($unsigned((reg2334 ?
                      $signed((7'h54)) : $signed(reg1903))) ?
                  $unsigned(reg2075[(2'h3):(2'h3)]) : $signed(reg1954[(2'h2):(1'h1)])));
              reg2448 = reg2431[(2'h2):(1'h0)];
              reg2449 <= reg2048;
            end
          reg2450 <= $signed($signed($signed({$unsigned(reg1885),
              $unsigned(reg1869)})));
        end
      reg2451 = ({$unsigned($signed((reg1785 >>> reg1883)))} ?
          (^~({(reg1869 ? reg2443 : reg2393),
                  (~^wire1896),
                  reg1982[(3'h6):(1'h1)]} ?
              reg2414[(3'h5):(2'h3)] : reg1905[(3'h4):(1'h0)])) : reg2248);
      reg2452 = $signed({$signed((~|(reg2016 ? reg1906 : wire1763)))});
    end
  assign wire2453 = reg1782;
  always
    @(posedge clk) begin
      reg2454 <= ((7'h49) & ((8'hb9) * $signed($signed((reg2009 ?
          (7'h57) : reg1816)))));
      reg2455 = (reg1954 ?
          reg2341 : (reg1836 ?
              reg2149[(1'h1):(1'h1)] : ($unsigned((8'h9f)) <= (+(reg2038 > reg1775)))));
      for (forvar2456 = (1'h0); (forvar2456 < (2'h3)); forvar2456 = (forvar2456 + (1'h1)))
        begin
          for (forvar2457 = (1'h0); (forvar2457 < (1'h0)); forvar2457 = (forvar2457 + (1'h1)))
            begin
              reg2458 = (~&($signed((~&reg2265)) ?
                  $unsigned(((~^reg2231) & (reg1928 ~^ reg2287))) : $signed({(reg2384 < (7'h57))})));
              reg2459 = (({reg2260[(4'ha):(3'h5)],
                  reg2252[(1'h1):(1'h1)]} & $signed(((reg2057 ?
                      (7'h44) : reg2359) ?
                  reg2039[(3'h6):(3'h6)] : $signed(reg2047)))) ~^ $signed((~^reg2422)));
              reg2460 = ($signed(((|$unsigned(reg2401)) ?
                      ((8'hb6) <<< (|reg1782)) : $unsigned($unsigned(reg1769)))) ?
                  ({(~&{(7'h43)})} ?
                      reg2320[(4'h8):(3'h6)] : reg2009[(4'h9):(1'h1)]) : $signed(reg2160));
              reg2461 <= $signed($unsigned((7'h58)));
            end
          reg2462 = $signed((+(~&$unsigned((wire1765 == reg2241)))));
          for (forvar2463 = (1'h0); (forvar2463 < (3'h5)); forvar2463 = (forvar2463 + (1'h1)))
            begin
              reg2464 <= ($unsigned(wire2207) & $unsigned((reg2150[(3'h4):(2'h3)] ?
                  {reg1808, reg2250} : ({reg1884} ?
                      $unsigned(reg2223) : (~^reg2150)))));
            end
          for (forvar2465 = (1'h0); (forvar2465 < (3'h6)); forvar2465 = (forvar2465 + (1'h1)))
            begin
              reg2466 <= $unsigned(($unsigned(((8'hbd) & reg1814[(1'h1):(1'h0)])) ?
                  {{reg2383,
                          ((7'h4b) ? reg1950 : reg2029),
                          (reg2252 > reg1942)},
                      $unsigned((reg2396 ^ reg1967)),
                      (^~$unsigned(reg2115))} : $signed($unsigned(((7'h4b) ?
                      reg1966 : (7'h4f))))));
              reg2467 = (7'h4c);
              reg2468 = ((reg2016[(3'h4):(3'h4)] ?
                  ($signed(reg2413[(2'h3):(2'h2)]) >> reg1803[(1'h0):(1'h0)]) : reg2015[(2'h3):(2'h2)]) >= (reg2002[(2'h2):(1'h0)] ^ (((reg1824 ?
                          reg2454 : reg2116) ?
                      reg1814[(2'h2):(2'h2)] : (~&reg2038)) ?
                  ((reg2038 ?
                      reg2023 : reg1956) >>> (~|reg1950)) : {$unsigned(reg2265),
                      (reg2450 ? reg2433 : (8'had))})));
              reg2469 = $signed(reg1790[(3'h7):(2'h2)]);
              reg2470 <= $unsigned(reg1962);
              reg2471 <= $signed(((((~reg2336) && (reg2258 <<< reg2324)) ?
                      ((reg2360 ?
                          (8'hac) : (8'hb0)) | $unsigned((7'h44))) : ($signed(reg1855) ?
                          (reg2160 ? reg2455 : reg2115) : reg2248)) ?
                  reg2107[(4'ha):(3'h4)] : reg2057));
            end
          reg2472 = reg2054;
          reg2473 = reg1932[(4'h9):(2'h3)];
        end
      for (forvar2474 = (1'h0); (forvar2474 < (2'h2)); forvar2474 = (forvar2474 + (1'h1)))
        begin
          reg2475 = $signed($signed((|reg2088[(1'h0):(1'h0)])));
          reg2476 <= $signed(reg1894);
          if ($unsigned((wire1763 ?
              $signed(((reg2437 ^~ (8'hb2)) >> reg1902[(4'ha):(3'h7)])) : (($signed(reg1935) ^~ $signed(reg1948)) - $unsigned(reg1861[(3'h6):(2'h3)])))))
            begin
              reg2477 <= $signed(reg2136[(3'h5):(3'h4)]);
              reg2478 <= (8'hbd);
              reg2479 <= reg2131[(1'h1):(1'h1)];
              reg2480 <= $unsigned($signed(((~&(reg2226 | reg2390)) ?
                  (~|(^~reg2355)) : ({reg1766} ?
                      (reg2422 >> reg2304) : $signed(reg2091)))));
              reg2481 = (reg2422[(3'h5):(3'h4)] ?
                  (-((reg1982 == reg2307[(2'h2):(1'h1)]) ^~ $signed({reg2344,
                      wire1765}))) : ((~{(reg2234 & reg1774)}) ?
                      (7'h4b) : $unsigned(reg2194[(2'h3):(2'h3)])));
              reg2482 <= ($unsigned(reg2401) ?
                  ((~$signed($unsigned(reg2320))) <<< (^$unsigned($unsigned(reg1791)))) : $unsigned((^~$signed((reg2149 - (7'h55))))));
              reg2483 = reg2153[(4'ha):(4'ha)];
            end
          else
            begin
              reg2477 <= {reg2242, $signed((!reg1803))};
              reg2481 = reg2383;
              reg2483 = (reg1826 ?
                  (+reg1932[(3'h6):(3'h6)]) : (reg2481 ?
                      (reg2078 ?
                          $signed((reg2153 || reg2231)) : ($unsigned(reg1962) ?
                              {reg2329,
                                  reg2007} : (~(7'h4f)))) : reg2226[(3'h7):(2'h3)]));
              reg2484 <= (^~$unsigned($unsigned((~&$signed(reg1894)))));
              reg2485 = $signed(reg2091);
            end
          reg2486 = (({reg1993[(3'h5):(1'h0)],
                      $signed(reg2410[(3'h5):(2'h2)])} ?
                  (reg1912 ?
                      reg2037 : {(~^reg2214),
                          (-reg1977)}) : (&$signed((reg2449 ?
                      reg2263 : reg1999)))) ?
              (($unsigned((-reg2380)) ?
                  ($unsigned(reg2275) ?
                      $unsigned(reg2057) : (reg2002 ?
                          reg1936 : reg2209)) : $unsigned((-reg2380))) + $unsigned((~|(^reg1790)))) : (+(8'hb5)));
          if (reg2368[(1'h1):(1'h0)])
            begin
              reg2487 <= (~|({(~^reg2484[(3'h6):(3'h5)])} >>> (reg2095 ~^ $unsigned(reg2152[(3'h4):(1'h1)]))));
              reg2488 = reg2094;
              reg2489 = reg2115[(4'ha):(2'h2)];
              reg2490 = $unsigned($signed(reg1987));
            end
          else
            begin
              reg2488 = $signed({(reg1905 ?
                      reg2124 : (^~((7'h53) ? reg1954 : reg2262))),
                  $signed($signed((^~reg2124)))});
            end
        end
    end
  always
    @(posedge clk) begin
      reg2491 = reg2335;
      if ({$signed((-reg2243)),
          reg1908,
          (reg1783[(3'h5):(3'h5)] ^ ((~|$unsigned(reg1905)) ?
              $signed((reg1981 ? reg2124 : reg2143)) : $unsigned({reg1911,
                  reg2018,
                  reg2070})))})
        begin
          for (forvar2492 = (1'h0); (forvar2492 < (1'h0)); forvar2492 = (forvar2492 + (1'h1)))
            begin
              reg2493 <= ($signed((|(reg1961[(3'h5):(2'h3)] && (reg2396 ?
                      reg2109 : (7'h50))))) ?
                  reg1864 : (~|$signed(reg1903)));
              reg2494 = ((+$unsigned($signed(reg2214))) <= ($unsigned(($unsigned(reg2023) > (8'hb0))) && {reg1800,
                  (reg1782 ? $signed(reg2301) : (reg2110 ? reg2002 : reg2066)),
                  ((reg1829 ? reg2243 : reg2414) ~^ $unsigned(reg2376))}));
              reg2495 = (reg2229[(5'h11):(4'hf)] >> ($signed((reg2320 ?
                      (reg2114 ? reg1900 : reg2218) : (wire1760 > reg2009))) ?
                  (((~|reg1768) ? reg2471[(1'h1):(1'h0)] : reg2238) ?
                      {((8'ha1) ? reg2444 : reg1826),
                          reg1979[(1'h1):(1'h0)],
                          $signed(reg1967)} : ((reg2380 >= reg2150) ?
                          (7'h4c) : (reg1981 ^ reg2410))) : reg2115[(5'h10):(3'h4)]));
            end
          if ((~&$unsigned(reg2333[(3'h5):(1'h0)])))
            begin
              reg2496 <= $unsigned(reg2214[(3'h7):(2'h3)]);
              reg2497 = (((+(!{(8'ha0), reg1942})) ?
                  $signed((reg1993[(3'h7):(3'h7)] ?
                      {reg1883, reg2333, reg2165} : (reg2046 ?
                          reg2220 : reg2054))) : $unsigned(((~|reg1847) ?
                      reg2115 : reg1906[(3'h5):(3'h5)]))) < reg2495);
              reg2498 <= (~^$unsigned((~&$unsigned(reg1848))));
              reg2499 <= reg2479[(4'hc):(2'h2)];
              reg2500 <= $unsigned(reg1998[(3'h7):(2'h2)]);
              reg2501 <= reg2284[(3'h5):(2'h3)];
              reg2502 <= {(|$signed(reg2440[(2'h3):(1'h1)])),
                  (~|reg1774),
                  (((((8'had) ? reg1768 : reg2073) ?
                          $signed((7'h4f)) : $signed(reg1790)) ?
                      (reg2214 ? reg2368 : {reg2136}) : {reg2135[(4'hc):(2'h2)],
                          reg1857,
                          reg2142[(2'h3):(1'h1)]}) << reg2027[(2'h3):(2'h2)])};
            end
          else
            begin
              reg2497 = ((~&{(!$unsigned(reg2198)),
                      ((reg2385 ? reg2477 : reg2115) <<< (~^reg1912))}) ?
                  reg1796 : {{((~^reg1956) ? reg1904 : reg2499)},
                      {($unsigned(reg2285) > reg2500[(4'hb):(4'h9)]),
                          {((8'h9d) >= reg2198)}},
                      reg2149});
              reg2498 <= (^reg1804);
              reg2503 = (~|(reg1858[(2'h2):(2'h2)] ?
                  reg1838[(4'h9):(2'h2)] : $signed(($unsigned(reg1771) > $signed(reg1806)))));
            end
          reg2504 = reg2056;
        end
      else
        begin
          reg2492 = $unsigned(reg2194[(2'h2):(1'h1)]);
          reg2494 = $signed($unsigned((7'h41)));
          reg2495 = (&$signed($unsigned(((reg1932 == (8'ha0)) - $unsigned((7'h42))))));
          for (forvar2496 = (1'h0); (forvar2496 < (3'h5)); forvar2496 = (forvar2496 + (1'h1)))
            begin
              reg2497 = (reg2324[(4'hc):(3'h6)] ?
                  $signed(reg1940[(4'hc):(3'h7)]) : $signed(reg2168[(2'h2):(2'h2)]));
              reg2498 <= (|(&{(!$signed(reg1832)),
                  ((&reg2440) || $unsigned(reg2417))}));
              reg2499 <= $signed(reg1785[(2'h3):(1'h1)]);
              reg2503 = ($signed(reg1891) || ($unsigned($unsigned($signed((7'h57)))) ?
                  wire1763[(2'h2):(1'h0)] : $unsigned(((reg2078 & reg2111) || (reg2334 ?
                      reg1794 : reg2384)))));
              reg2504 = $unsigned(((+$unsigned($signed(reg1908))) ?
                  reg2023[(3'h4):(3'h4)] : reg2180));
              reg2505 <= (((^~reg1900) || (reg2242[(4'ha):(3'h7)] ?
                  reg1857[(4'h8):(1'h1)] : (+reg2027))) & reg2418);
              reg2506 = ((((reg1991 ? $unsigned(reg2056) : $unsigned(reg1868)) ?
                  $signed($unsigned(reg1950)) : $signed((reg1808 >= reg1904))) != $signed(reg2094[(3'h6):(1'h1)])) + (^~((+{(7'h4e)}) ?
                  reg2356 : ($unsigned(reg1880) ?
                      ((8'hb6) ? reg1840 : reg2153) : reg2334))));
            end
          if ($signed((~&$signed(({reg2471,
              reg2215} != reg2248[(4'h8):(4'h8)])))))
            begin
              reg2507 = $signed(reg1857);
              reg2508 <= ((~^((~&(reg2470 || reg1917)) >>> reg2444)) && {(8'haf)});
              reg2509 = $signed($signed($signed(reg1861)));
              reg2510 <= (-$unsigned(reg2503));
              reg2511 = (reg2200 ?
                  reg1875 : (reg1981 ? reg2505[(3'h4):(2'h3)] : reg2299));
            end
          else
            begin
              reg2508 <= (reg2214 || $unsigned(reg2064));
              reg2509 = $unsigned(reg1853[(2'h2):(1'h1)]);
              reg2511 = {(reg1785[(3'h5):(2'h3)] ^ ((!reg2180) ?
                      $signed(reg1962) : $unsigned(((7'h50) ^ reg2242)))),
                  {((reg2017 ^ (reg2010 > reg2243)) ?
                          reg1956 : ({(8'ha4),
                              (8'hba),
                              reg2299} >= $unsigned((8'h9c))))},
                  reg2307};
            end
        end
      for (forvar2512 = (1'h0); (forvar2512 < (2'h2)); forvar2512 = (forvar2512 + (1'h1)))
        begin
          for (forvar2513 = (1'h0); (forvar2513 < (3'h5)); forvar2513 = (forvar2513 + (1'h1)))
            begin
              reg2514 <= reg2466;
              reg2515 = {reg2241[(4'ha):(3'h4)]};
              reg2516 <= reg2078[(4'hf):(4'hc)];
              reg2517 = (-(~&reg2229));
              reg2518 <= ((~&$unsigned($unsigned((8'ha9)))) ?
                  (8'hb8) : $unsigned(((^~reg1915[(4'ha):(2'h2)]) >= ((reg1869 ?
                      reg2215 : reg1833) << reg2407))));
              reg2519 = $unsigned(reg2258);
            end
          for (forvar2520 = (1'h0); (forvar2520 < (2'h3)); forvar2520 = (forvar2520 + (1'h1)))
            begin
              reg2521 = $unsigned($signed(reg1804));
              reg2522 = reg1824;
              reg2523 <= $signed({(reg2047[(1'h1):(1'h0)] | $signed(reg1855)),
                  (~reg1979),
                  $signed($unsigned(reg1775[(2'h2):(1'h1)]))});
            end
          if (reg1775)
            begin
              reg2524 = $unsigned($unsigned($unsigned((8'ha0))));
              reg2525 <= ({$unsigned(((reg2091 + reg2384) ?
                          $unsigned(reg2150) : reg1800)),
                      {$unsigned((reg2054 ? reg2518 : reg2450)),
                          (reg1936[(4'he):(4'h8)] != (reg2494 && reg2409)),
                          ((+reg1978) ?
                              (reg2243 ? reg2148 : reg2115) : {reg2021})}} ?
                  $unsigned($unsigned($signed(reg1811))) : (((~$unsigned(reg1985)) ?
                      reg1811[(5'h13):(4'hb)] : $signed((reg2502 > reg2066))) > reg1914[(5'h11):(4'h8)]));
              reg2526 = reg2344[(3'h4):(1'h1)];
            end
          else
            begin
              reg2524 = reg2334[(3'h4):(1'h0)];
              reg2525 <= reg1826[(5'h10):(1'h0)];
              reg2527 <= ((~&reg2466[(5'h16):(5'h16)]) ?
                  ({reg2295[(4'hc):(2'h3)],
                      ($unsigned(reg1791) ?
                          (reg2047 ? reg2052 : reg1769) : {reg1833}),
                      reg1860} != $signed(reg2341)) : reg1893);
              reg2528 <= (-(!(reg2370 ^ ((reg2503 != reg1962) ?
                  ((7'h54) != reg2344) : (|reg2284)))));
              reg2529 = $signed(wire2208);
              reg2530 = $unsigned(((7'h4c) << reg2342[(2'h3):(2'h3)]));
            end
        end
    end
  always
    @(posedge clk) begin
      if ((reg2446[(4'ha):(2'h2)] ?
          reg2065[(3'h5):(3'h4)] : $signed((((reg2136 != reg2071) ?
              (|reg1782) : $unsigned(reg1774)) <<< (^$signed(reg2454))))))
        begin
          reg2531 <= reg2015[(4'h8):(2'h2)];
          reg2532 = $unsigned($signed({(!$signed(reg2302)),
              reg2238[(3'h5):(2'h2)]}));
          if (reg2000[(4'hf):(4'he)])
            begin
              reg2533 = $unsigned((^reg2098[(5'h18):(4'he)]));
            end
          else
            begin
              reg2534 <= $signed(($signed(reg1777[(5'h12):(3'h5)]) ?
                  (((reg1942 ~^ reg2454) ?
                      (reg2007 ?
                          reg2304 : reg2095) : $unsigned(reg2286)) + ($signed(reg2039) & reg2340[(4'hf):(3'h5)])) : (~reg2143[(4'h8):(2'h2)])));
              reg2535 <= reg2088[(4'h9):(3'h7)];
              reg2536 <= (reg2177[(3'h4):(1'h0)] < ($unsigned(reg2446[(2'h3):(1'h1)]) << {(7'h43),
                  reg2226[(5'h11):(4'hf)]}));
            end
          for (forvar2537 = (1'h0); (forvar2537 < (1'h0)); forvar2537 = (forvar2537 + (1'h1)))
            begin
              reg2538 <= $unsigned($signed(reg2010[(4'ha):(4'ha)]));
              reg2539 = $signed((-$unsigned(((reg1843 | reg2393) < (~reg1891)))));
            end
          if ($signed(reg1932))
            begin
              reg2540 = $signed(reg2078[(3'h4):(2'h3)]);
              reg2541 = $unsigned((($signed((8'hae)) << (|(^~reg1878))) <<< {((reg2408 * reg2176) >> (~^reg2169)),
                  $unsigned(((8'hbf) ~^ reg2336))}));
              reg2542 = $signed(reg1962[(4'h8):(3'h5)]);
              reg2543 = $unsigned($unsigned({$unsigned(reg1962)}));
            end
          else
            begin
              reg2540 = reg2217[(5'h10):(4'h9)];
              reg2541 = (reg2270[(1'h0):(1'h0)] ~^ ((~&((reg1766 ?
                          reg2131 : (8'hb1)) ?
                      reg2073[(3'h5):(3'h5)] : wire2453[(2'h2):(1'h1)])) ?
                  $unsigned(reg1933[(3'h7):(3'h5)]) : (+reg2073[(3'h5):(3'h4)])));
              reg2544 <= (~&$signed((reg1966 < $unsigned((reg1902 ?
                  reg1977 : reg1818)))));
              reg2545 = reg2057[(4'hb):(3'h4)];
              reg2546 <= (reg1936[(1'h1):(1'h1)] == {(((^reg2010) - $unsigned(reg2066)) & ($signed((8'hbd)) > reg2271[(4'he):(3'h6)])),
                  (&$unsigned($signed(reg1771)))});
            end
        end
      else
        begin
          for (forvar2531 = (1'h0); (forvar2531 < (2'h3)); forvar2531 = (forvar2531 + (1'h1)))
            begin
              reg2532 = $signed(reg1884[(5'h10):(4'hc)]);
            end
          reg2534 <= (((($signed((8'ha5)) ?
                  reg1822 : $signed(reg2198)) != {((8'had) ?
                      reg1912 : reg1857)}) || reg2110) ?
              {$unsigned(reg1775),
                  $unsigned((7'h50))} : ((~{$unsigned(reg2418)}) ?
                  ($unsigned(((8'hbf) | reg2249)) || ($unsigned(reg1946) << $signed(reg2493))) : {{(8'hb2)},
                      $unsigned(reg1814)}));
          if ((+$signed($unsigned({(-reg2015),
              {reg2260},
              ((8'hb1) - (7'h40))}))))
            begin
              reg2537 = $unsigned($signed($signed(reg2152[(2'h2):(1'h0)])));
              reg2539 = (^((^$unsigned((reg2333 >> reg1981))) + (reg2437[(3'h5):(1'h0)] ?
                  $signed(reg2268) : {$unsigned(reg2344),
                      $signed((8'hb7)),
                      (reg2368 ? reg2046 : reg2401)})));
            end
          else
            begin
              reg2535 <= (~&(~^((~|$unsigned(reg2390)) != wire1896)));
              reg2537 = reg2322;
              reg2539 = $signed(($unsigned({$unsigned((7'h4b))}) | reg1954[(1'h1):(1'h0)]));
              reg2544 <= reg2243;
            end
          if ((reg2248[(4'ha):(3'h6)] ?
              ((&$unsigned((wire2208 ?
                  reg2318 : reg1878))) ~^ reg2286[(3'h6):(3'h5)]) : $signed({$signed($signed(reg2407))})))
            begin
              reg2546 <= reg2440[(2'h2):(1'h0)];
              reg2547 <= $unsigned($signed(($unsigned(reg1843) == reg2285[(1'h0):(1'h0)])));
              reg2548 <= $unsigned($unsigned((reg2248 ?
                  (((7'h43) ^ reg1998) ?
                      reg2396 : $unsigned(reg1811)) : $signed(reg2523))));
            end
          else
            begin
              reg2545 = {(~|$unsigned(reg1800[(3'h7):(2'h2)]))};
              reg2549 = (-$unsigned($unsigned((-(reg1981 ?
                  reg2333 : reg2160)))));
              reg2550 = $unsigned($signed($signed(reg2109[(4'hf):(4'he)])));
              reg2551 <= reg2152[(2'h3):(2'h3)];
              reg2552 <= $signed(((!($signed(reg1987) < $unsigned(reg1836))) << (~|($unsigned(reg1897) >> reg2376))));
              reg2553 <= (+$unsigned(reg2391));
              reg2554 = reg2229;
            end
          reg2555 = $unsigned(reg1785);
          reg2556 <= $unsigned($signed({reg1926,
              ($signed(reg1908) == $unsigned(reg2404)),
              $unsigned(reg1788[(4'he):(4'ha)])}));
        end
      reg2557 = (8'hb2);
      reg2558 <= (8'hab);
      for (forvar2559 = (1'h0); (forvar2559 < (1'h0)); forvar2559 = (forvar2559 + (1'h1)))
        begin
          if ({{reg1950[(4'hc):(4'ha)],
                  ((&reg2135) ? reg2548 : reg1993[(4'ha):(3'h4)]),
                  $signed((^~(!reg1869)))}})
            begin
              reg2560 <= ($signed((reg2053 * $signed((7'h55)))) ?
                  (~|wire2208[(5'h19):(5'h16)]) : (reg2440[(5'h17):(5'h11)] > $signed(reg1782[(3'h4):(2'h2)])));
              reg2561 = (({reg2094} ?
                      {(|(reg2299 ? reg2549 : reg2523)),
                          $signed((reg1903 ? reg1768 : reg1932)),
                          reg2318} : $signed(reg1961)) ?
                  {reg1848[(1'h1):(1'h1)], reg2325[(1'h0):(1'h0)]} : reg2243);
              reg2562 <= $unsigned(({(~&(reg2017 ? reg2370 : reg2240)),
                  {$signed(reg2476),
                      {reg2297, reg2042, reg2359},
                      (reg2433 ? reg2482 : reg1933)},
                  reg2408[(4'hc):(2'h2)]} ^~ $signed(reg2023[(4'hb):(4'ha)])));
            end
          else
            begin
              reg2560 <= reg2150;
              reg2561 = reg2150;
              reg2562 <= $signed((&(((~reg2447) ?
                  $signed(reg2160) : reg2385[(5'h11):(2'h3)]) ^ (&$signed(reg2464)))));
              reg2563 = {(~^(reg2264[(3'h6):(3'h5)] + reg2054[(4'hb):(4'hb)])),
                  ((-($unsigned(reg1838) ? $signed(reg1900) : reg2401)) ?
                      (^{(reg2052 != reg2527),
                          (reg2093 ?
                              reg2409 : reg1838)}) : (-(reg2214[(3'h6):(1'h1)] << $signed((8'h9e)))))};
              reg2564 <= reg2195;
            end
          reg2565 = reg2380[(5'h10):(5'h10)];
          reg2566 = reg2562;
          reg2567 <= $signed(reg2160[(2'h2):(2'h2)]);
        end
    end
  assign wire2568 = $unsigned((^~($unsigned(reg2065[(3'h4):(3'h4)]) ?
                        reg2409[(1'h1):(1'h0)] : {$unsigned(reg1800),
                            reg2218[(1'h0):(1'h0)],
                            (reg2221 | reg2200)})));
  always
    @(posedge clk) begin
      reg2569 <= reg2518;
      reg2570 <= {(reg2385[(5'h12):(4'h9)] ?
              reg1846[(1'h0):(1'h0)] : {$unsigned(((7'h40) <= reg2546))}),
          {($signed({reg1826, reg2501, reg2171}) ?
                  (^~reg2042) : reg1998[(3'h5):(1'h0)]),
              (({reg1985} ?
                  (reg1897 >= (7'h58)) : $unsigned(reg1811)) << $signed({reg2499,
                  reg2496}))},
          $unsigned($signed(reg2391))};
      reg2571 = $signed($signed(((reg1999 ? reg1811 : (|reg2066)) << reg1766)));
      for (forvar2572 = (1'h0); (forvar2572 < (2'h2)); forvar2572 = (forvar2572 + (1'h1)))
        begin
          reg2573 <= reg1943;
          reg2574 = {((+$unsigned($unsigned(reg2238))) | $unsigned(reg2132[(5'h13):(4'hb)])),
              {reg2263,
                  (-($unsigned(reg1818) * {reg2258})),
                  {($unsigned(reg2564) ? reg2004 : (~&reg2018)),
                      ($signed(reg1894) > reg1928),
                      reg2271}},
              {(+{reg2168}),
                  ({(~reg1911), reg1961, $signed(reg1914)} >= (~{reg2057})),
                  ((reg2121[(4'h8):(3'h6)] >= (reg2477 * reg2000)) ?
                      (reg2436 ^ $signed(reg1799)) : (&$unsigned((7'h48))))}};
          reg2575 = $unsigned($unsigned({{{reg2015}, reg1894}}));
          if ($signed($signed($signed($signed($signed((8'hac)))))))
            begin
              reg2576 = ($signed((~{$unsigned((7'h45)),
                  reg1819[(4'ha):(3'h6)]})) == reg1838);
              reg2577 = $unsigned(($unsigned((|reg2142)) ~^ ($unsigned(reg2226[(4'ha):(3'h6)]) ?
                  (reg2320[(1'h1):(1'h0)] ~^ (~|reg2318)) : reg2187[(5'h1c):(2'h3)])));
              reg2578 <= reg2556[(5'h15):(1'h1)];
              reg2579 = (|(~&reg2115[(5'h10):(3'h7)]));
              reg2580 = $unsigned({((~&(~|reg2028)) ?
                      $unsigned((~|reg2514)) : ({reg1995} ?
                          (reg2009 ?
                              reg2198 : (7'h56)) : (reg2057 - (8'hb5))))});
              reg2581 = ((-reg1860[(5'h16):(4'hd)]) ?
                  $unsigned((8'hb9)) : (!((-$signed(reg2420)) ?
                      $unsigned((~&reg2437)) : reg2578[(3'h7):(3'h5)])));
            end
          else
            begin
              reg2578 <= reg2318;
              reg2582 <= ((((+$signed((8'hb0))) >= reg1905) ?
                      ($unsigned((reg2066 == (7'h40))) ?
                          reg2479 : reg1782[(3'h6):(3'h6)]) : ((^(reg1977 ?
                              (8'hab) : reg1824)) ?
                          reg2418[(5'h1e):(5'h17)] : reg2342)) ?
                  reg2014[(3'h4):(1'h1)] : $signed($unsigned($signed(reg1993[(3'h7):(3'h5)]))));
              reg2583 = $unsigned(reg2355[(3'h5):(3'h4)]);
              reg2584 = (~|$unsigned($signed({(+(7'h4a))})));
            end
          reg2585 = reg1966[(2'h3):(1'h0)];
        end
      if (($unsigned($signed(($unsigned(reg2324) ?
          reg2238[(3'h4):(1'h1)] : reg2355))) ~^ (reg2351 >>> (~|(8'haf)))))
        begin
          for (forvar2586 = (1'h0); (forvar2586 < (1'h0)); forvar2586 = (forvar2586 + (1'h1)))
            begin
              reg2587 = reg2109;
              reg2588 = {({(~&(reg2587 ? reg2056 : (7'h52))),
                          $signed(((8'ha4) && reg1829)),
                          reg2136[(3'h4):(1'h1)]} ?
                      reg1966 : $unsigned($unsigned({reg2054}))),
                  $signed((((reg2400 ? reg2238 : wire1761) ^ (reg2322 ?
                          reg2466 : reg2039)) ?
                      reg2111 : reg1818[(3'h7):(3'h6)])),
                  reg1774};
              reg2589 <= (($signed(((+reg1804) ?
                  {reg2229} : $signed(reg2449))) + (8'hbb)) >> reg2305);
            end
          reg2590 = reg1774[(2'h2):(2'h2)];
          reg2591 <= $signed((~|$signed(reg2017)));
        end
      else
        begin
          reg2586 = $signed((-(reg2305 ?
              ($unsigned(reg2116) ?
                  {reg2057, reg2200, reg2341} : (-(7'h49))) : {reg2420,
                  $unsigned(reg1880),
                  reg2009[(3'h7):(3'h5)]})));
          if ((-($signed(reg2518[(3'h7):(1'h1)]) << ({(|reg1788),
              (^~reg2525),
              {(8'h9e), reg2569, reg2287}} & ($signed(reg2447) ?
              $unsigned(reg2413) : (reg1771 ? reg1914 : reg2523))))))
            begin
              reg2587 = {$signed((((reg2299 ?
                          (7'h4b) : reg1819) ~^ $unsigned((7'h4c))) ?
                      (+reg1794) : ($unsigned(reg2148) >> (~&(7'h55))))),
                  {(reg1768[(4'h8):(1'h0)] ^ reg2215[(1'h0):(1'h0)])},
                  reg2356[(4'he):(4'ha)]};
              reg2588 = {reg2558[(4'hd):(3'h7)],
                  (^{$unsigned((&reg2020))}),
                  $signed(reg2355)};
              reg2589 <= ((($unsigned(reg2171[(1'h0):(1'h0)]) ?
                      ((+reg1832) ?
                          (^~reg2010) : $signed(reg2028)) : (~^(reg2578 >= (7'h46)))) ?
                  reg2393 : {$signed((reg2004 ? reg2117 : reg2311)),
                      reg2053[(5'h1a):(5'h10)],
                      $signed($signed(reg2478))}) <= (~^$signed($signed(reg2548))));
              reg2591 <= $unsigned(((reg2575[(4'he):(4'he)] ?
                  (~^(reg2114 ?
                      reg2305 : reg1891)) : reg1822) < $signed(reg2265[(4'h9):(1'h1)])));
              reg2592 <= (reg2564 ? reg1788 : (-reg2215));
              reg2593 = (+(($signed(reg1905) ?
                      $unsigned(reg2316[(3'h4):(1'h0)]) : $signed({reg2376})) ?
                  reg1869[(1'h0):(1'h0)] : $signed(((8'hb9) >= (reg2220 ?
                      reg2115 : reg2535)))));
              reg2594 = {reg2293[(3'h4):(3'h4)]};
            end
          else
            begin
              reg2589 <= reg1926;
              reg2591 <= {(~&(+$signed((~^reg2308)))), reg2248};
              reg2593 = (~^(reg2243[(1'h0):(1'h0)] ?
                  (^~reg2118[(1'h1):(1'h1)]) : (reg2065 ?
                      {reg1966[(4'hb):(2'h3)],
                          reg2414[(4'hb):(4'hb)]} : reg2268)));
              reg2594 = reg1995[(2'h2):(2'h2)];
              reg2595 <= (&(~^reg1822));
              reg2596 = reg2308[(4'hd):(3'h7)];
            end
          if ((~$unsigned(reg1911)))
            begin
              reg2597 = ((-({(reg2516 >> reg2470), reg1880} ?
                  ((reg2289 ? reg2307 : reg2552) >> (reg2002 ?
                      reg2436 : reg1903)) : {reg2218,
                      $unsigned((8'ha3))})) ~^ (~&(+$unsigned((reg2047 ^ wire1764)))));
              reg2598 = $signed(({wire1762[(3'h6):(2'h3)],
                  ((reg1935 ?
                      reg2270 : (8'h9d)) ^~ reg2422)} < $unsigned(reg1791[(2'h2):(1'h1)])));
              reg2599 = reg2534;
              reg2600 = (~|(((8'hbe) >= $unsigned((^~reg2476))) * $unsigned((7'h4a))));
              reg2601 <= (8'ha6);
              reg2602 = reg2384;
            end
          else
            begin
              reg2597 = (reg2220[(3'h4):(1'h1)] ?
                  $signed(reg2407[(2'h3):(2'h3)]) : $signed(reg2249));
              reg2601 <= $unsigned(((7'h52) != (~|(-reg2307))));
              reg2603 <= {(+reg2073[(2'h3):(2'h3)])};
              reg2604 <= $unsigned(reg2599);
            end
          for (forvar2605 = (1'h0); (forvar2605 < (1'h0)); forvar2605 = (forvar2605 + (1'h1)))
            begin
              reg2606 <= (8'had);
              reg2607 <= (^reg2516[(2'h2):(1'h1)]);
              reg2608 = ($signed(reg2088) ?
                  reg2493[(5'h12):(3'h7)] : (($unsigned(reg1948) ?
                          reg2383 : (|{reg2047, (7'h40)})) ?
                      $signed((+reg2078)) : {reg1861[(2'h2):(1'h1)],
                          $unsigned($unsigned(reg1774)),
                          $unsigned((|reg2567))}));
              reg2609 = reg1950;
              reg2610 <= $unsigned(((-$signed((reg1892 > reg2409))) - $signed(($unsigned((8'ha5)) <<< ((8'haa) != (8'ha3))))));
              reg2611 = ($signed(((~|(reg2023 - reg2385)) ?
                      reg2336[(3'h4):(2'h3)] : (^(^~reg2470)))) ?
                  $signed((((reg1928 ^~ reg2376) ?
                      reg1936 : (8'hbf)) & {reg2131,
                      (~reg2238),
                      $signed(reg2588)})) : reg2482[(3'h7):(2'h3)]);
              reg2612 <= reg2408;
            end
          if ((-(8'hb1)))
            begin
              reg2613 <= ((-reg2585[(3'h6):(3'h4)]) ?
                  ($signed((~^$unsigned((8'ha1)))) & (^reg1869)) : ((~&reg1902) >> ((-$signed(reg2067)) ?
                      (|{reg1839}) : $unsigned(reg1816))));
              reg2614 = $unsigned(reg2243);
              reg2615 = $unsigned((-((forvar2586 ?
                  (^~reg2383) : $signed(reg2196)) >= (reg2114 ^ reg2505[(1'h1):(1'h0)]))));
            end
          else
            begin
              reg2613 <= reg1981;
              reg2616 <= $signed(reg2289);
              reg2617 = reg2240;
            end
        end
      if ($signed(((reg2168[(4'h8):(3'h7)] != ((reg2006 ?
          reg1906 : reg2477) + (~^reg1806))) >> (reg2581[(1'h0):(1'h0)] ?
          reg2220[(4'h9):(2'h2)] : (8'ha4)))))
        begin
          reg2618 <= (((~^(^reg2093)) ^~ (-(~$signed(reg1804)))) > {$signed(($signed((8'hb6)) ~^ (reg2596 ^~ reg1979))),
              $signed($signed($unsigned((7'h45))))});
          reg2619 = $signed(reg1833);
          if (reg1982[(2'h2):(1'h1)])
            begin
              reg2620 <= reg1861[(2'h3):(2'h2)];
              reg2621 = $signed($unsigned({((reg2418 ? wire2043 : reg1979) ?
                      {reg2593, reg1833, reg1912} : {reg2508}),
                  (reg2360 ^~ ((8'hbd) == reg1923))}));
              reg2622 <= $signed(reg2142[(2'h3):(2'h3)]);
            end
          else
            begin
              reg2621 = $signed(((~&$unsigned($signed((7'h58)))) ?
                  ($signed({reg2336}) + (8'hab)) : reg2585[(4'h9):(4'h8)]));
              reg2622 <= (reg2500[(2'h2):(2'h2)] ?
                  reg2066[(1'h1):(1'h0)] : $unsigned(reg2595));
              reg2623 <= (~&{reg2214, (+reg1869[(1'h0):(1'h0)])});
              reg2624 <= $unsigned((($signed((~&reg2356)) ?
                      ($signed(reg2470) <= {reg1875}) : reg2108) ?
                  (((-reg2589) ? $signed(reg2576) : (~^reg2250)) ?
                      $signed(reg2305) : ((reg1880 ? reg2596 : reg2621) ?
                          reg1990[(2'h3):(2'h3)] : $signed(reg2305))) : $signed($unsigned(reg2608[(4'he):(4'h9)]))));
              reg2625 <= reg2108[(3'h7):(3'h5)];
            end
          reg2626 <= $signed(reg2020);
        end
      else
        begin
          reg2619 = $unsigned((reg2335 - ($unsigned(reg1933[(4'hf):(3'h7)]) & reg2263[(2'h3):(2'h2)])));
          if (((($signed(reg2436[(1'h1):(1'h0)]) != $signed((^reg2297))) > ({{(8'ha9)},
              {reg2030}} && reg2594[(3'h4):(3'h4)])) || ($unsigned($signed((reg1977 ?
                  reg2570 : reg2322))) ?
              (($unsigned(reg2148) < {reg2594}) || (~^$unsigned(reg2287))) : (^reg1877[(2'h3):(1'h0)]))))
            begin
              reg2620 <= (7'h4b);
              reg2621 = (($unsigned(((reg1791 <<< reg2471) ?
                          (!reg2356) : reg2321)) ?
                      $signed($unsigned((reg2535 && reg1999))) : $unsigned(($unsigned((7'h49)) ?
                          $unsigned(reg1891) : (reg2553 ^ reg2150)))) ?
                  (({((8'hae) | reg2168), reg2293, reg2224[(2'h2):(1'h0)]} ?
                      reg2318 : reg2165) <<< $unsigned(((reg2271 ?
                      reg2570 : (7'h40)) <<< (reg1800 ?
                      reg2252 : (7'h46))))) : {reg2332,
                      ($signed(reg1825[(4'h8):(3'h4)]) << (7'h51))});
              reg2627 = ({reg2216[(2'h2):(1'h0)],
                  (reg2581[(1'h0):(1'h0)] ? reg2544 : reg2446),
                  reg2241} << (reg2446[(3'h7):(2'h2)] ^~ {($signed(reg1981) >= (~^reg2573)),
                  reg2547[(4'hf):(1'h0)]}));
              reg2628 <= {(reg1904[(3'h7):(1'h0)] ?
                      (reg2000 ?
                          $signed(reg2209[(2'h3):(2'h2)]) : (!(+reg2311))) : (~|((~|reg2413) && (~reg1833))))};
              reg2629 = (~|($unsigned(reg2258[(2'h2):(2'h2)]) <<< (+$unsigned(((8'ha3) ?
                  reg2477 : reg2604)))));
              reg2630 = (($unsigned((-reg1777[(4'hb):(4'h8)])) + reg2271[(1'h0):(1'h0)]) * ({($unsigned(reg1806) ?
                          $signed(reg2249) : reg2143[(2'h2):(1'h0)]),
                      reg2514[(1'h1):(1'h0)],
                      {reg2564[(3'h7):(1'h1)], $unsigned(reg2344), reg2518}} ?
                  reg1771 : reg1796[(1'h1):(1'h0)]));
            end
          else
            begin
              reg2621 = reg2258;
              reg2622 <= (reg1995[(5'h14):(5'h13)] ?
                  reg2336[(3'h4):(3'h4)] : {(reg1885 ^ (reg1912[(4'ha):(3'h4)] ~^ (reg2538 ?
                          reg1790 : (8'ha5))))});
              reg2627 = (7'h44);
              reg2628 <= $signed($signed($signed((reg2132 ?
                  (|reg2308) : reg2591[(1'h1):(1'h0)]))));
              reg2631 <= reg2301;
              reg2632 = (+reg1814);
              reg2633 <= $signed(reg2479);
            end
        end
    end
  always
    @(posedge clk) begin
      reg2634 <= {(reg2325[(1'h0):(1'h0)] < $signed(((~reg1987) >= reg1978))),
          reg2527};
    end
endmodule