
(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param1156 = {({(((8'h9d) <= (8'ha6)) ~^ (^~(8'h9c))), (~{(7'h41), (8'had)})} >> {({(8'h9f)} | ((8'haa) * (8'hbc))), (+((8'ha0) ? (7'h48) : (8'ha1)))})})
(y, clk, wire200, wire199, wire198, wire197, wire196);
  output wire [(32'hd58):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire200;
  input wire [(5'h13):(1'h0)] wire199;
  input wire signed [(5'h12):(1'h0)] wire198;
  input wire [(5'h10):(1'h0)] wire197;
  input wire [(3'h6):(1'h0)] wire196;
  wire [(4'h8):(1'h0)] wire1154;
  wire [(4'he):(1'h0)] wire1094;
  wire [(5'h16):(1'h0)] wire436;
  wire signed [(4'he):(1'h0)] wire389;
  wire signed [(2'h2):(1'h0)] wire336;
  wire signed [(3'h7):(1'h0)] wire291;
  wire [(5'h15):(1'h0)] wire287;
  wire signed [(4'ha):(1'h0)] wire286;
  wire [(5'h15):(1'h0)] wire284;
  wire signed [(5'h12):(1'h0)] wire204;
  wire [(5'h18):(1'h0)] wire203;
  reg [(3'h6):(1'h0)] reg477 = (1'h0);
  reg [(3'h4):(1'h0)] reg474 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg473 = (1'h0);
  reg [(5'h16):(1'h0)] reg470 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg469 = (1'h0);
  reg [(3'h6):(1'h0)] reg466 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg462 = (1'h0);
  reg [(2'h2):(1'h0)] reg460 = (1'h0);
  reg [(3'h6):(1'h0)] reg457 = (1'h0);
  reg [(4'he):(1'h0)] reg452 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg450 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg445 = (1'h0);
  reg [(4'h8):(1'h0)] reg444 = (1'h0);
  reg [(2'h2):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg440 = (1'h0);
  reg [(3'h7):(1'h0)] reg439 = (1'h0);
  reg [(5'h10):(1'h0)] reg435 = (1'h0);
  reg [(4'hd):(1'h0)] reg433 = (1'h0);
  reg [(4'hd):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg431 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg429 = (1'h0);
  reg [(5'h11):(1'h0)] reg428 = (1'h0);
  reg [(4'ha):(1'h0)] reg425 = (1'h0);
  reg [(3'h5):(1'h0)] reg419 = (1'h0);
  reg [(4'h9):(1'h0)] reg418 = (1'h0);
  reg [(4'hd):(1'h0)] reg415 = (1'h0);
  reg [(3'h4):(1'h0)] reg413 = (1'h0);
  reg [(5'h15):(1'h0)] reg412 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg410 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg409 = (1'h0);
  reg [(5'h13):(1'h0)] reg407 = (1'h0);
  reg [(2'h3):(1'h0)] reg403 = (1'h0);
  reg [(5'h10):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg398 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg394 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg391 = (1'h0);
  reg [(3'h5):(1'h0)] reg390 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg377 = (1'h0);
  reg [(4'hb):(1'h0)] reg385 = (1'h0);
  reg [(5'h16):(1'h0)] reg381 = (1'h0);
  reg [(5'h10):(1'h0)] reg380 = (1'h0);
  reg [(4'hd):(1'h0)] reg379 = (1'h0);
  reg [(4'hd):(1'h0)] reg375 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg374 = (1'h0);
  reg [(5'h16):(1'h0)] reg368 = (1'h0);
  reg [(5'h14):(1'h0)] reg367 = (1'h0);
  reg [(5'h14):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg365 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg362 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg361 = (1'h0);
  reg [(4'ha):(1'h0)] reg352 = (1'h0);
  reg [(5'h17):(1'h0)] reg347 = (1'h0);
  reg [(5'h11):(1'h0)] reg346 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg345 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg333 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg328 = (1'h0);
  reg [(5'h10):(1'h0)] reg327 = (1'h0);
  reg [(5'h12):(1'h0)] reg326 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg325 = (1'h0);
  reg [(4'hd):(1'h0)] reg322 = (1'h0);
  reg [(4'hf):(1'h0)] reg319 = (1'h0);
  reg [(5'h18):(1'h0)] reg317 = (1'h0);
  reg [(4'h9):(1'h0)] reg315 = (1'h0);
  reg [(5'h11):(1'h0)] reg310 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg306 = (1'h0);
  reg [(5'h11):(1'h0)] reg304 = (1'h0);
  reg [(4'h8):(1'h0)] reg303 = (1'h0);
  reg [(5'h17):(1'h0)] reg301 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg298 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg295 = (1'h0);
  reg [(4'hd):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg290 = (1'h0);
  reg [(5'h15):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1097 = (1'h0);
  reg [(4'h9):(1'h0)] reg1099 = (1'h0);
  reg [(4'he):(1'h0)] reg1102 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1104 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1101 = (1'h0);
  reg [(2'h2):(1'h0)] reg1108 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1109 = (1'h0);
  reg [(4'he):(1'h0)] reg1114 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1117 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1118 = (1'h0);
  reg [(3'h7):(1'h0)] reg1121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1124 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1126 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1127 = (1'h0);
  reg [(4'h9):(1'h0)] reg1130 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1132 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1135 = (1'h0);
  reg [(4'hd):(1'h0)] reg1136 = (1'h0);
  reg [(3'h4):(1'h0)] reg1138 = (1'h0);
  reg [(3'h6):(1'h0)] reg1139 = (1'h0);
  reg [(5'h16):(1'h0)] reg1141 = (1'h0);
  reg [(4'h8):(1'h0)] reg1142 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1146 = (1'h0);
  reg [(3'h7):(1'h0)] reg1148 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1149 = (1'h0);
  reg [(5'h15):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1151 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1152 = (1'h0);
  reg [(4'ha):(1'h0)] reg1153 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1137 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1147 = (1'h0);
  reg [(4'he):(1'h0)] reg1145 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1144 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1143 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1137 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1134 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1133 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1131 = (1'h0);
  reg [(4'ha):(1'h0)] reg1129 = (1'h0);
  reg [(4'h9):(1'h0)] reg1128 = (1'h0);
  reg [(5'h14):(1'h0)] reg1125 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1123 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1122 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1120 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1119 = (1'h0);
  reg [(2'h2):(1'h0)] reg1116 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1115 = (1'h0);
  reg [(3'h7):(1'h0)] reg1113 = (1'h0);
  reg [(4'hc):(1'h0)] reg1112 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1111 = (1'h0);
  reg [(2'h2):(1'h0)] reg1110 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1107 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1106 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1103 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1102 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1099 = (1'h0);
  reg [(4'hf):(1'h0)] reg1105 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1103 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1101 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1100 = (1'h0);
  reg [(3'h7):(1'h0)] reg1098 = (1'h0);
  reg [(4'hd):(1'h0)] reg476 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg475 = (1'h0);
  reg [(4'hb):(1'h0)] reg472 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg471 = (1'h0);
  reg [(4'hd):(1'h0)] reg468 = (1'h0);
  reg [(5'h10):(1'h0)] reg467 = (1'h0);
  reg [(5'h11):(1'h0)] reg465 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg464 = (1'h0);
  reg [(5'h10):(1'h0)] forvar463 = (1'h0);
  reg [(5'h14):(1'h0)] reg461 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar459 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg458 = (1'h0);
  reg [(3'h7):(1'h0)] reg456 = (1'h0);
  reg [(5'h15):(1'h0)] reg455 = (1'h0);
  reg [(5'h12):(1'h0)] forvar454 = (1'h0);
  reg [(5'h16):(1'h0)] reg453 = (1'h0);
  reg [(4'h8):(1'h0)] forvar451 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar443 = (1'h0);
  reg [(5'h13):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg448 = (1'h0);
  reg [(5'h12):(1'h0)] reg447 = (1'h0);
  reg [(3'h6):(1'h0)] reg446 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg443 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg442 = (1'h0);
  reg [(4'he):(1'h0)] reg438 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar437 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar434 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg430 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar427 = (1'h0);
  reg [(3'h5):(1'h0)] reg426 = (1'h0);
  reg [(3'h6):(1'h0)] reg424 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg423 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg422 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg421 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg420 = (1'h0);
  reg [(4'he):(1'h0)] reg417 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar416 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg414 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg411 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg408 = (1'h0);
  reg [(5'h12):(1'h0)] reg406 = (1'h0);
  reg [(5'h11):(1'h0)] reg405 = (1'h0);
  reg [(4'h8):(1'h0)] reg404 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg402 = (1'h0);
  reg [(5'h13):(1'h0)] reg401 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg399 = (1'h0);
  reg [(4'he):(1'h0)] reg397 = (1'h0);
  reg [(5'h15):(1'h0)] reg395 = (1'h0);
  reg [(2'h2):(1'h0)] forvar392 = (1'h0);
  reg [(5'h12):(1'h0)] reg382 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg388 = (1'h0);
  reg [(4'hf):(1'h0)] forvar387 = (1'h0);
  reg [(5'h14):(1'h0)] reg386 = (1'h0);
  reg [(5'h14):(1'h0)] reg384 = (1'h0);
  reg [(3'h7):(1'h0)] reg383 = (1'h0);
  reg [(4'hb):(1'h0)] forvar382 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg378 = (1'h0);
  reg [(4'he):(1'h0)] forvar377 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg376 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg370 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar364 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg373 = (1'h0);
  reg [(5'h13):(1'h0)] reg372 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg371 = (1'h0);
  reg [(4'h9):(1'h0)] forvar370 = (1'h0);
  reg [(5'h13):(1'h0)] reg369 = (1'h0);
  reg [(5'h15):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg363 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar360 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg359 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg358 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar357 = (1'h0);
  reg [(4'hb):(1'h0)] reg356 = (1'h0);
  reg [(3'h5):(1'h0)] forvar355 = (1'h0);
  reg [(5'h10):(1'h0)] reg354 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg353 = (1'h0);
  reg [(3'h7):(1'h0)] reg351 = (1'h0);
  reg [(5'h14):(1'h0)] reg350 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar348 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar344 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg342 = (1'h0);
  reg [(2'h3):(1'h0)] reg341 = (1'h0);
  reg [(5'h14):(1'h0)] reg340 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg339 = (1'h0);
  reg [(4'hd):(1'h0)] forvar338 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar337 = (1'h0);
  reg [(4'h8):(1'h0)] reg335 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg332 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg331 = (1'h0);
  reg [(4'h9):(1'h0)] reg330 = (1'h0);
  reg [(4'hc):(1'h0)] reg329 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg324 = (1'h0);
  reg [(5'h12):(1'h0)] reg323 = (1'h0);
  reg [(2'h2):(1'h0)] reg321 = (1'h0);
  reg [(5'h15):(1'h0)] reg320 = (1'h0);
  reg [(3'h7):(1'h0)] reg318 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar316 = (1'h0);
  reg signed [(4'he):(1'h0)] reg314 = (1'h0);
  reg [(4'hc):(1'h0)] reg313 = (1'h0);
  reg [(4'hd):(1'h0)] reg312 = (1'h0);
  reg [(5'h10):(1'h0)] reg311 = (1'h0);
  reg [(3'h5):(1'h0)] forvar310 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar304 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg309 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg302 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg299 = (1'h0);
  reg [(3'h5):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg293 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg292 = (1'h0);
  reg [(5'h15):(1'h0)] reg289 = (1'h0);
  reg [(4'hb):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg201 = (1'h0);
  assign y = {wire1154,
                 wire1094,
                 wire436,
                 wire389,
                 wire336,
                 wire291,
                 wire287,
                 wire286,
                 wire284,
                 wire204,
                 wire203,
                 reg477,
                 reg474,
                 reg473,
                 reg470,
                 reg469,
                 reg466,
                 reg462,
                 reg460,
                 reg457,
                 reg452,
                 reg450,
                 reg449,
                 reg445,
                 reg444,
                 reg441,
                 reg440,
                 reg439,
                 reg435,
                 reg433,
                 reg432,
                 reg431,
                 reg429,
                 reg428,
                 reg425,
                 reg419,
                 reg418,
                 reg415,
                 reg413,
                 reg412,
                 reg410,
                 reg409,
                 reg407,
                 reg403,
                 reg400,
                 reg398,
                 reg396,
                 reg394,
                 reg393,
                 reg391,
                 reg390,
                 reg377,
                 reg385,
                 reg381,
                 reg380,
                 reg379,
                 reg375,
                 reg374,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg362,
                 reg361,
                 reg352,
                 reg347,
                 reg346,
                 reg345,
                 reg334,
                 reg333,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg322,
                 reg319,
                 reg317,
                 reg315,
                 reg310,
                 reg308,
                 reg307,
                 reg306,
                 reg304,
                 reg303,
                 reg301,
                 reg298,
                 reg295,
                 reg294,
                 reg290,
                 reg1096,
                 reg1097,
                 reg1099,
                 reg1102,
                 reg1104,
                 reg1101,
                 reg1108,
                 reg1109,
                 reg1114,
                 reg1117,
                 reg1118,
                 reg1121,
                 reg1124,
                 reg1126,
                 reg1127,
                 reg1130,
                 reg1132,
                 reg1135,
                 reg1136,
                 reg1138,
                 reg1139,
                 reg1141,
                 reg1142,
                 reg1146,
                 reg1148,
                 reg1149,
                 reg1150,
                 reg1151,
                 reg1152,
                 reg1153,
                 reg1137,
                 reg1147,
                 reg1145,
                 reg1144,
                 forvar1143,
                 reg1140,
                 forvar1137,
                 forvar1134,
                 reg1133,
                 forvar1131,
                 reg1129,
                 reg1128,
                 reg1125,
                 forvar1123,
                 forvar1122,
                 reg1120,
                 reg1119,
                 reg1116,
                 reg1115,
                 reg1113,
                 reg1112,
                 reg1111,
                 reg1110,
                 reg1107,
                 reg1106,
                 reg1103,
                 forvar1102,
                 forvar1099,
                 reg1105,
                 forvar1103,
                 forvar1101,
                 reg1100,
                 reg1098,
                 reg476,
                 reg475,
                 reg472,
                 reg471,
                 reg468,
                 reg467,
                 reg465,
                 reg464,
                 forvar463,
                 reg461,
                 forvar459,
                 reg458,
                 reg456,
                 reg455,
                 forvar454,
                 reg453,
                 forvar451,
                 forvar443,
                 reg437,
                 reg448,
                 reg447,
                 reg446,
                 reg443,
                 reg442,
                 reg438,
                 forvar437,
                 forvar434,
                 reg430,
                 forvar427,
                 reg426,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg417,
                 forvar416,
                 reg414,
                 reg411,
                 reg408,
                 reg406,
                 reg405,
                 reg404,
                 reg402,
                 reg401,
                 reg399,
                 reg397,
                 reg395,
                 forvar392,
                 reg382,
                 reg388,
                 forvar387,
                 reg386,
                 reg384,
                 reg383,
                 forvar382,
                 reg378,
                 forvar377,
                 reg376,
                 reg370,
                 forvar364,
                 reg373,
                 reg372,
                 reg371,
                 forvar370,
                 reg369,
                 reg364,
                 reg363,
                 forvar360,
                 reg359,
                 reg358,
                 forvar357,
                 reg356,
                 forvar355,
                 reg354,
                 reg353,
                 reg351,
                 reg350,
                 reg349,
                 forvar348,
                 forvar344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 forvar338,
                 forvar337,
                 reg335,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg324,
                 reg323,
                 reg321,
                 reg320,
                 reg318,
                 forvar316,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 forvar310,
                 forvar304,
                 reg309,
                 reg305,
                 reg302,
                 reg300,
                 reg299,
                 reg297,
                 reg296,
                 reg293,
                 reg292,
                 reg289,
                 reg288,
                 reg202,
                 reg201,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg201 = (($unsigned($unsigned($unsigned(wire197))) ?
              $unsigned($signed(wire198[(1'h1):(1'h1)])) : (wire198[(2'h2):(2'h2)] >> ((8'ha2) ?
                  (wire197 - wire198) : {wire200, (7'h40)}))) ?
          (7'h47) : (~&(^~$unsigned($unsigned(wire200)))));
      reg202 = (~{(~&{(wire199 ? (8'haf) : reg201), {reg201, reg201}}),
          (($unsigned(wire198) ?
              ((8'ha7) ?
                  wire199 : reg201) : $signed(wire200)) <<< wire199[(4'he):(4'hc)])});
    end
  assign wire203 = ((~$unsigned(wire199[(4'ha):(3'h5)])) << $unsigned(($unsigned(wire199[(4'he):(4'ha)]) == $signed((8'hb3)))));
  assign wire204 = wire198;
  assign wire286 = ({wire196,
                           (wire197 ?
                               (7'h49) : ({wire196} ?
                                   wire198[(2'h2):(1'h1)] : $signed(wire197)))} ?
                       $signed(($unsigned(wire284[(1'h1):(1'h1)]) == (~^$signed(wire198)))) : (~(($signed((8'hae)) <<< (wire196 << wire284)) ?
                           {(wire200 ? (8'h9f) : wire199)} : (8'h9d))));
  assign wire287 = $signed(wire197[(2'h2):(2'h2)]);
  always
    @(posedge clk) begin
      reg288 = $signed(wire284);
      reg289 = (^$unsigned($unsigned((wire286 ?
          wire196[(2'h2):(1'h1)] : $signed(wire284)))));
      reg290 <= reg288[(4'h9):(1'h1)];
    end
  assign wire291 = {(~^({(wire199 ? wire200 : wire196),
                           $unsigned(wire284)} ^ (^wire203[(5'h17):(2'h2)]))),
                       (wire198[(4'h9):(1'h0)] ?
                           (((wire203 ?
                                   wire203 : wire284) || $unsigned(wire196)) ?
                               $unsigned(wire287) : ((wire284 ?
                                   wire197 : wire199) & $signed(wire204))) : wire200)};
  always
    @(posedge clk) begin
      if ($signed(($signed(($signed((7'h42)) ^~ $signed(reg290))) ?
          $unsigned($signed(wire204[(4'h8):(1'h1)])) : $signed(wire197))))
        begin
          reg292 = (~&(({(wire204 ? (7'h44) : wire204)} ?
              ((reg290 ~^ wire196) >>> (wire197 ?
                  wire287 : wire197)) : ((&wire287) ?
                  ((8'hae) ?
                      wire197 : wire203) : $unsigned(wire284))) >>> {((wire196 ?
                      wire197 : wire291) ?
                  $signed(wire291) : wire200)}));
          reg293 = {wire196[(2'h3):(1'h0)]};
          if ((+$signed((7'h42))))
            begin
              reg294 <= wire204[(4'hc):(2'h3)];
              reg295 <= ($signed($signed(wire291[(3'h5):(3'h5)])) ?
                  (reg293 ?
                      {{wire203},
                          $signed(((8'hb0) > wire200))} : $signed($unsigned((-wire291)))) : wire197[(4'hf):(3'h5)]);
              reg296 = wire198;
            end
          else
            begin
              reg296 = wire204[(4'hf):(4'hb)];
              reg297 = (|reg294[(1'h1):(1'h1)]);
              reg298 <= ({reg293[(4'hc):(4'h9)],
                      {wire284[(5'h15):(4'hb)], wire284}} ?
                  ((reg293[(5'h13):(3'h6)] << $unsigned(reg294[(1'h0):(1'h0)])) | $unsigned(($signed(reg292) << {wire197,
                      reg293}))) : wire284);
              reg299 = wire197[(2'h2):(1'h1)];
              reg300 = wire200[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg294 <= (($unsigned(($unsigned((8'h9e)) ~^ ((8'ha0) ?
                  reg298 : wire197))) > $signed(((wire199 ? wire291 : reg296) ?
                  {wire203, wire198} : (8'hb1)))) ?
              (8'hae) : ((+({reg293} ? wire284 : reg295[(2'h3):(1'h1)])) ?
                  $signed((&(reg292 != wire286))) : wire199));
        end
      reg301 <= {$signed($signed(wire291)), reg295[(3'h4):(1'h0)]};
      reg302 = (($unsigned(wire196[(3'h6):(3'h5)]) ?
              $signed(wire291) : wire204) ?
          $unsigned($signed(((wire200 == reg296) ?
              (~^wire196) : wire199[(4'h9):(3'h6)]))) : ($signed(((^wire203) ^~ (wire196 ?
                  wire287 : wire199))) ?
              wire286 : (~|reg290)));
    end
  always
    @(posedge clk) begin
      if ((&($unsigned(wire196) * (!{wire198, $unsigned(wire286)}))))
        begin
          if ((|(8'hb7)))
            begin
              reg303 <= ((^~(~&$signed(wire196))) < ($unsigned(($signed((8'hb8)) ?
                      $unsigned(reg301) : reg290)) ?
                  ({(wire197 - wire196), (&wire203)} - ($unsigned(wire196) ?
                      $signed((8'hbc)) : reg301)) : ({(~^wire286)} * ({wire204} ?
                      (reg295 & wire198) : (reg294 ? reg290 : reg290)))));
              reg304 <= $unsigned(wire198);
            end
          else
            begin
              reg305 = wire196;
              reg306 <= reg303[(2'h2):(1'h1)];
            end
          reg307 <= {reg304[(5'h11):(2'h3)]};
          reg308 <= wire204;
          reg309 = $unsigned((reg304 != ($unsigned(reg304) ~^ (!(~&(8'hb1))))));
          reg310 <= ((~&($signed({wire198, reg305}) ?
              (^(&wire197)) : $signed($signed(reg295)))) - ($unsigned((~^$unsigned(wire291))) < {reg290[(2'h3):(2'h3)]}));
        end
      else
        begin
          reg303 <= $unsigned(wire284);
          for (forvar304 = (1'h0); (forvar304 < (2'h3)); forvar304 = (forvar304 + (1'h1)))
            begin
              reg306 <= $signed(reg308);
              reg309 = (reg307[(3'h5):(3'h4)] || $unsigned($unsigned(reg305[(3'h5):(3'h4)])));
            end
          for (forvar310 = (1'h0); (forvar310 < (3'h4)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 = ((7'h49) ?
                  ((((~wire196) ^~ (reg306 - (8'hb3))) >>> ($signed(forvar310) ?
                          reg294 : forvar310[(1'h0):(1'h0)])) ?
                      reg304 : (^((8'hbc) >= ((8'ha6) <= forvar310)))) : (~&reg306));
              reg312 = (8'hbc);
              reg313 = ((reg301[(4'ha):(3'h7)] ?
                      wire287[(4'h8):(3'h5)] : $unsigned(forvar310[(1'h0):(1'h0)])) ?
                  wire204[(3'h4):(2'h3)] : (&(|(((8'ha7) ?
                      (8'hb3) : forvar310) && $signed(forvar304)))));
              reg314 = $signed((reg304 ?
                  $unsigned((8'h9c)) : ({$signed(reg313)} && (forvar310 ?
                      wire199 : reg305[(1'h0):(1'h0)]))));
              reg315 <= ($unsigned(((wire198[(4'ha):(3'h4)] < $signed(reg301)) & wire203)) >>> $unsigned(reg295));
            end
        end
      for (forvar316 = (1'h0); (forvar316 < (2'h2)); forvar316 = (forvar316 + (1'h1)))
        begin
          if ((8'hb4))
            begin
              reg317 <= (+wire199);
              reg318 = wire204;
              reg319 <= reg303;
            end
          else
            begin
              reg318 = (-(&(($signed(wire200) ?
                      $unsigned(reg301) : forvar310[(1'h0):(1'h0)]) ?
                  $unsigned({(8'hbc)}) : {(-reg298),
                      forvar304[(1'h0):(1'h0)]})));
              reg319 <= reg307;
              reg320 = forvar304[(2'h3):(2'h3)];
            end
          if (reg303)
            begin
              reg321 = reg317[(5'h17):(5'h11)];
              reg322 <= (~|reg290[(3'h5):(3'h5)]);
            end
          else
            begin
              reg322 <= $unsigned($signed(reg322[(4'hd):(3'h7)]));
              reg323 = $signed((^$unsigned(((wire204 != forvar310) ~^ (wire197 >= reg321)))));
              reg324 = (wire198 ?
                  ({reg317,
                          ((reg320 ? reg298 : wire284) != $unsigned(wire196))} ?
                      reg320 : reg319[(4'hc):(4'hb)]) : (8'hb4));
              reg325 <= $unsigned((reg301[(1'h0):(1'h0)] >>> $signed(wire198)));
            end
          if ($unsigned(reg322[(1'h0):(1'h0)]))
            begin
              reg326 <= wire284;
              reg327 <= $signed($signed($unsigned($unsigned((&reg303)))));
              reg328 <= (~^(wire287[(4'h8):(3'h5)] ?
                  {({wire198, reg323} ?
                          reg306[(3'h5):(3'h4)] : wire197[(4'ha):(3'h7)]),
                      wire287[(3'h6):(3'h6)]} : (8'h9d)));
              reg329 = ($unsigned((^~(8'haa))) ~^ {reg326[(1'h0):(1'h0)]});
            end
          else
            begin
              reg329 = reg290;
              reg330 = (reg307 <<< $unsigned($unsigned(reg305)));
              reg331 = {$signed($unsigned($signed((~&wire200))))};
            end
        end
    end
  always
    @(posedge clk) begin
      reg332 = reg303[(3'h4):(2'h2)];
      reg333 <= $unsigned($signed((-wire199)));
      reg334 <= reg326[(3'h5):(1'h1)];
      reg335 = reg319[(1'h1):(1'h0)];
    end
  assign wire336 = $signed({($signed((wire204 ~^ reg328)) ?
                           reg306 : {$unsigned(reg298)})});
  always
    @(posedge clk) begin
      for (forvar337 = (1'h0); (forvar337 < (1'h0)); forvar337 = (forvar337 + (1'h1)))
        begin
          for (forvar338 = (1'h0); (forvar338 < (3'h4)); forvar338 = (forvar338 + (1'h1)))
            begin
              reg339 = (&($signed(((^~reg306) >= $signed(reg301))) << (~&{(!(8'hba)),
                  (^wire336)})));
              reg340 = $signed({reg294});
              reg341 = reg317[(4'ha):(2'h2)];
              reg342 = reg341[(1'h0):(1'h0)];
              reg343 = wire198;
            end
          for (forvar344 = (1'h0); (forvar344 < (3'h4)); forvar344 = (forvar344 + (1'h1)))
            begin
              reg345 <= $unsigned(((!(!$signed((8'ha4)))) > wire284[(3'h7):(2'h3)]));
              reg346 <= reg345;
            end
          reg347 <= {(^$unsigned({wire284, $signed((8'haf))})),
              $signed({((~^reg339) + (wire287 ? wire286 : reg310)), reg315})};
        end
      for (forvar348 = (1'h0); (forvar348 < (2'h3)); forvar348 = (forvar348 + (1'h1)))
        begin
          reg349 = (+$unsigned(wire203));
          if ({reg307[(2'h3):(1'h1)], reg304[(1'h0):(1'h0)]})
            begin
              reg350 = reg326;
              reg351 = reg304[(5'h11):(3'h5)];
              reg352 <= reg306;
              reg353 = (&$unsigned(reg322));
              reg354 = ($signed((~|$signed((reg328 ? reg325 : reg325)))) ?
                  $signed(((^~reg349) <= (8'ha8))) : ((reg304 ?
                      reg298 : (~|reg351[(3'h4):(1'h1)])) & $unsigned($unsigned(reg315))));
            end
          else
            begin
              reg350 = (&{((-reg346[(1'h0):(1'h0)]) >> $unsigned((reg328 ?
                      forvar348 : reg345)))});
            end
        end
      for (forvar355 = (1'h0); (forvar355 < (1'h0)); forvar355 = (forvar355 + (1'h1)))
        begin
          reg356 = forvar338;
        end
    end
  always
    @(posedge clk) begin
      for (forvar357 = (1'h0); (forvar357 < (2'h3)); forvar357 = (forvar357 + (1'h1)))
        begin
          reg358 = {(wire200[(4'ha):(1'h1)] & ((reg317[(5'h17):(1'h1)] || $unsigned(reg310)) & (|(wire286 ?
                  wire286 : wire203)))),
              (wire196 ? reg333 : reg295[(3'h4):(1'h0)])};
        end
      reg359 = reg358[(4'h9):(3'h7)];
      for (forvar360 = (1'h0); (forvar360 < (1'h1)); forvar360 = (forvar360 + (1'h1)))
        begin
          reg361 <= ({wire336} ?
              (&(($unsigned(reg328) ?
                  (reg315 ?
                      (8'ha9) : wire198) : (|wire284)) && wire291[(3'h5):(2'h2)])) : reg326);
          reg362 <= (reg345 ?
              {reg345,
                  (~|$unsigned((wire204 ?
                      reg295 : reg352)))} : (&$signed((8'haf))));
          reg363 = $signed($unsigned(reg362));
        end
      if (reg346[(4'ha):(2'h2)])
        begin
          if ($signed($unsigned(forvar360)))
            begin
              reg364 = ({$unsigned($signed(reg303[(3'h4):(3'h4)]))} ?
                  ({wire286[(3'h5):(2'h2)], (|(reg345 ? (7'h45) : (7'h40)))} ?
                      $signed((-reg301)) : (8'ha5)) : $unsigned(reg362));
              reg365 <= {reg298[(1'h0):(1'h0)]};
              reg366 <= (~|(+reg301[(3'h4):(1'h1)]));
              reg367 <= ({wire286[(4'h9):(3'h6)]} >> ((&(reg328[(1'h1):(1'h0)] ?
                      (8'ha4) : (reg315 ? reg359 : reg326))) ?
                  (~&reg359) : wire336[(1'h0):(1'h0)]));
              reg368 <= reg303;
            end
          else
            begin
              reg364 = $signed($unsigned({(reg352 ? (reg364 < reg317) : reg308),
                  ((&reg307) ^ (~&reg290))}));
              reg365 <= reg333[(4'hc):(4'h8)];
              reg369 = $signed((&(($unsigned(wire203) && ((8'hb0) & wire284)) ?
                  $unsigned($signed(reg298)) : $signed({reg326, reg301}))));
            end
          for (forvar370 = (1'h0); (forvar370 < (1'h0)); forvar370 = (forvar370 + (1'h1)))
            begin
              reg371 = {reg327[(1'h0):(1'h0)], wire196[(2'h2):(2'h2)]};
              reg372 = wire336[(1'h0):(1'h0)];
              reg373 = $unsigned(reg319);
              reg374 <= (($signed(reg345[(3'h7):(3'h6)]) >= $signed((reg371 ?
                  (reg301 >>> reg347) : reg361[(3'h5):(2'h2)]))) * $unsigned(reg319));
              reg375 <= (+(wire196[(2'h2):(2'h2)] == reg317));
            end
        end
      else
        begin
          for (forvar364 = (1'h0); (forvar364 < (1'h1)); forvar364 = (forvar364 + (1'h1)))
            begin
              reg369 = ($signed((~$signed($signed((7'h45))))) | reg345[(1'h0):(1'h0)]);
              reg370 = reg306;
              reg371 = forvar370;
              reg372 = $unsigned((7'h46));
              reg374 <= $signed($signed(reg365[(4'ha):(2'h2)]));
            end
          reg376 = $unsigned(((^((-reg358) ?
                  wire196[(1'h0):(1'h0)] : $signed(wire287))) ?
              ((~&wire199) <<< {wire204[(1'h0):(1'h0)],
                  wire200}) : ((reg347[(3'h7):(3'h5)] ?
                      forvar360[(1'h0):(1'h0)] : (^reg352)) ?
                  $unsigned((reg346 <<< reg308)) : reg301[(5'h15):(5'h15)])));
        end
      if ($signed(($unsigned(reg303) ?
          {(^~(wire286 ? (8'h9d) : wire197)),
              ($signed(reg307) ?
                  $signed((8'ha1)) : (~&reg345))} : $unsigned((^~(wire336 << forvar357))))))
        begin
          for (forvar377 = (1'h0); (forvar377 < (2'h2)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg378 = forvar370[(2'h2):(1'h0)];
              reg379 <= ((reg306 ? $unsigned((!$unsigned(reg376))) : (8'h9c)) ?
                  {((reg370 ? {reg294} : $signed((8'hae))) ?
                          ($unsigned(reg290) != forvar377[(2'h3):(2'h3)]) : $unsigned((~&reg307)))} : $signed($signed($signed($signed(reg358)))));
              reg380 <= ((~&wire197) ?
                  wire291[(1'h1):(1'h0)] : $unsigned({($unsigned(wire291) << (^~reg346))}));
              reg381 <= ((($unsigned($unsigned(reg325)) | reg376[(4'ha):(2'h2)]) <<< $unsigned($signed((forvar357 ?
                      reg308 : forvar370)))) ?
                  reg308[(3'h4):(3'h4)] : ($signed(forvar370) >> $unsigned(reg379[(1'h1):(1'h1)])));
            end
          for (forvar382 = (1'h0); (forvar382 < (1'h1)); forvar382 = (forvar382 + (1'h1)))
            begin
              reg383 = (~^reg301[(5'h16):(5'h10)]);
              reg384 = {{wire197[(3'h4):(3'h4)]},
                  $unsigned(forvar377[(3'h4):(3'h4)])};
            end
          reg385 <= reg298[(1'h0):(1'h0)];
          reg386 = reg295;
          for (forvar387 = (1'h0); (forvar387 < (1'h0)); forvar387 = (forvar387 + (1'h1)))
            begin
              reg388 = ($signed((($unsigned(reg381) ?
                      (~reg383) : wire203[(1'h1):(1'h1)]) * $signed((reg345 ?
                      reg358 : wire336)))) ?
                  (8'h9c) : (($signed($unsigned(reg358)) << ($unsigned(reg364) == (wire286 ?
                      (8'hbd) : reg327))) ^ (($signed(reg303) ?
                      reg372 : (forvar364 ?
                          reg306 : reg298)) < $unsigned($signed(reg303)))));
            end
        end
      else
        begin
          reg377 <= reg298;
          if (((&{((wire291 || reg371) ?
                      (^reg365) : (reg290 ? reg306 : wire203)),
                  ((forvar377 * wire291) ? {reg333} : (~&reg334))}) ?
              ($signed((forvar360 ? (&reg322) : (wire284 ? wire287 : reg363))) ?
                  {reg372[(4'ha):(1'h1)], (^(wire336 << reg290))} : (((reg362 ?
                      reg374 : reg334) && {reg315,
                      reg352}) == forvar387[(4'hc):(1'h0)])) : ($unsigned(wire197) != reg376[(5'h10):(2'h3)])))
            begin
              reg378 = (~^reg328[(2'h2):(2'h2)]);
              reg382 = $unsigned($signed($signed((~&$signed(reg359)))));
              reg383 = (((((~&reg295) | ((7'h49) ?
                      reg345 : reg303)) - ((+reg304) ?
                      (~forvar387) : (wire199 ? (8'hab) : reg365))) ?
                  $unsigned(reg373[(4'h8):(3'h5)]) : $signed((((8'hbb) ?
                      reg385 : (7'h49)) & ((7'h46) ?
                      wire197 : wire196)))) && (($signed(((8'ha2) || reg378)) ?
                      reg382[(4'h9):(1'h0)] : ($signed(wire196) ?
                          (|(8'hb9)) : $unsigned((8'h9c)))) ?
                  ($signed(forvar370[(2'h2):(1'h0)]) + $signed(reg352[(4'h8):(4'h8)])) : forvar357[(2'h3):(2'h2)]));
            end
          else
            begin
              reg379 <= {(8'ha3),
                  (forvar377 && {$signed((!reg310)),
                      {wire204, (forvar370 <= reg317)}})};
            end
          reg384 = (($unsigned(reg301) - wire198) ?
              forvar364 : ((forvar364 ?
                      (reg363[(4'hf):(4'hf)] * (reg359 ?
                          wire197 : (8'hb1))) : $unsigned(forvar360[(1'h1):(1'h1)])) ?
                  ((8'h9f) >>> (~^(^reg295))) : (!$unsigned($unsigned(forvar370)))));
          reg386 = {($unsigned((8'hab)) ?
                  (-wire287) : (({reg352, forvar387} ?
                          (&wire199) : $signed(reg301)) ?
                      $unsigned($unsigned(wire199)) : (^~((8'ha4) ?
                          forvar377 : forvar370)))),
              $unsigned(reg374[(1'h1):(1'h0)])};
        end
    end
  assign wire389 = $signed(reg310[(3'h4):(2'h2)]);
  always
    @(posedge clk) begin
      reg390 <= reg377;
    end
  always
    @(posedge clk) begin
      reg391 <= {$signed($signed(reg317[(1'h1):(1'h1)]))};
      for (forvar392 = (1'h0); (forvar392 < (2'h3)); forvar392 = (forvar392 + (1'h1)))
        begin
          reg393 <= {{$signed($signed({reg368, reg365}))}};
          reg394 <= reg377;
          reg395 = (-((($unsigned(reg379) ?
                      (reg325 ? reg315 : wire286) : wire197[(2'h2):(2'h2)]) ?
                  ($signed((8'hb7)) ^~ (~&reg390)) : reg365[(3'h4):(1'h1)]) ?
              ($unsigned($unsigned(reg317)) ?
                  ((reg379 ?
                      wire286 : reg326) < $signed(reg380)) : (-wire284)) : $unsigned((8'haf))));
          reg396 <= reg379;
        end
      if ((8'hb6))
        begin
          reg397 = (|(!reg326[(4'h9):(4'h9)]));
        end
      else
        begin
          if ((&wire203[(5'h16):(5'h13)]))
            begin
              reg398 <= reg395;
              reg399 = ($signed($signed(reg368)) <<< (($signed(reg391[(5'h15):(4'h9)]) || {$unsigned(reg362)}) ~^ {$signed(reg362[(4'hd):(1'h1)]),
                  reg390[(1'h1):(1'h1)]}));
              reg400 <= $unsigned((&reg294));
              reg401 = (!{reg390[(3'h5):(1'h1)],
                  (wire284 ?
                      ($unsigned(reg295) ?
                          (reg315 >>> reg294) : reg319) : reg327)});
            end
          else
            begin
              reg397 = reg374[(3'h6):(3'h5)];
              reg399 = reg322[(3'h6):(1'h0)];
              reg401 = (reg398 ^ $signed(reg400[(5'h10):(4'h8)]));
              reg402 = (^reg399[(3'h4):(1'h0)]);
            end
          if (reg304)
            begin
              reg403 <= (~^(~^((reg345 ? (reg401 == forvar392) : reg325) ?
                  $unsigned(wire204[(5'h10):(3'h7)]) : ((reg366 < reg294) ?
                      (reg317 ? wire286 : reg375) : reg326))));
            end
          else
            begin
              reg404 = forvar392;
              reg405 = (reg390 && $unsigned((8'h9c)));
              reg406 = (reg347 ?
                  reg379[(1'h1):(1'h1)] : {((&reg294) ?
                          ({reg352, reg326} ?
                              (|(8'ha4)) : $unsigned(reg403)) : (((8'hb6) == reg317) & $unsigned((8'ha1))))});
              reg407 <= {($signed(($unsigned(reg385) ?
                          (wire284 ? reg307 : reg294) : $signed(reg406))) ?
                      $unsigned(($unsigned(reg400) ?
                          (reg385 != (8'hba)) : $unsigned((8'hbb)))) : reg290),
                  $unsigned(reg362[(4'hd):(3'h6)])};
            end
          reg408 = reg362;
        end
    end
  always
    @(posedge clk) begin
      if ((~|($unsigned(($signed(reg334) ?
              reg310 : (reg377 ? reg301 : reg381))) ?
          {((~|reg379) ~^ reg400[(4'h8):(3'h5)])} : reg345[(2'h3):(2'h3)])))
        begin
          reg409 <= wire287;
          reg410 <= reg294[(1'h0):(1'h0)];
        end
      else
        begin
          reg409 <= wire197;
          reg411 = ({reg294, (+$signed(reg381))} - $unsigned({{reg379},
              (((8'h9f) ? reg303 : reg409) ?
                  (wire286 << reg303) : $signed(wire199))}));
          if ($signed(((reg308 ? wire286 : reg381) <= wire198)))
            begin
              reg412 <= wire197[(1'h1):(1'h1)];
              reg413 <= $signed($signed((+$unsigned($signed(reg374)))));
            end
          else
            begin
              reg412 <= ((^~$unsigned((7'h43))) ?
                  (((&$unsigned((8'hbd))) ?
                      $unsigned(reg315[(2'h3):(2'h3)]) : $signed($unsigned(reg409))) < reg301) : reg381[(4'hc):(4'hb)]);
              reg414 = $unsigned(reg367);
              reg415 <= wire389;
            end
          for (forvar416 = (1'h0); (forvar416 < (2'h3)); forvar416 = (forvar416 + (1'h1)))
            begin
              reg417 = (~(reg303 >>> (^~(|$unsigned(wire198)))));
              reg418 <= (&{$unsigned($signed($signed((8'hb2)))),
                  reg398[(4'h9):(3'h7)]});
              reg419 <= wire198;
            end
          if (((reg367[(3'h6):(3'h5)] & reg304) ?
              $unsigned($unsigned({$signed(reg381)})) : $signed((wire389 >> reg306))))
            begin
              reg420 = (reg346 ?
                  wire204 : ((+reg380[(2'h2):(2'h2)]) ?
                      $signed((((8'hb6) ?
                          wire199 : reg328) ~^ $signed(reg306))) : reg310[(4'hb):(2'h2)]));
              reg421 = reg394[(1'h1):(1'h1)];
              reg422 = (reg413[(1'h0):(1'h0)] ?
                  wire197[(3'h5):(3'h4)] : (~|wire389[(2'h2):(1'h0)]));
            end
          else
            begin
              reg420 = ((~|reg394) ?
                  $signed((&$unsigned($unsigned(forvar416)))) : $unsigned(reg400));
            end
        end
      reg423 = $unsigned((^{(8'ha8), reg333[(4'hc):(4'hb)]}));
      reg424 = (reg391 != (~^$signed($signed(reg391[(4'hb):(4'h9)]))));
      reg425 <= (((^reg418[(3'h7):(3'h5)]) ?
          $signed((^$unsigned(reg415))) : (($signed(reg352) ^~ (8'ha4)) ~^ $unsigned((reg368 == (8'hb8))))) != ($unsigned(wire287[(4'hc):(1'h0)]) ?
          reg419[(1'h0):(1'h0)] : reg421));
    end
  always
    @(posedge clk) begin
      reg426 = (-wire197[(4'hf):(4'he)]);
      for (forvar427 = (1'h0); (forvar427 < (1'h1)); forvar427 = (forvar427 + (1'h1)))
        begin
          if (((8'hb9) ?
              {(reg380 ?
                      (~(reg385 && reg400)) : $unsigned((wire198 ?
                          reg317 : reg400)))} : reg413[(3'h4):(2'h2)]))
            begin
              reg428 <= (((!reg365) ~^ (reg418 & (reg347 < (~|reg400)))) - (!reg333[(4'hb):(2'h3)]));
              reg429 <= reg412[(5'h14):(4'hd)];
              reg430 = (($signed($signed($signed(wire286))) ?
                  (reg365[(1'h1):(1'h1)] >>> reg393) : ({reg308[(3'h5):(3'h4)],
                          wire336[(1'h1):(1'h0)]} ?
                      reg374 : $unsigned(reg385[(4'ha):(3'h5)]))) >>> reg400);
            end
          else
            begin
              reg428 <= $signed(reg298[(3'h5):(3'h4)]);
              reg430 = $signed(reg415);
            end
          reg431 <= $unsigned($signed(wire286[(2'h2):(2'h2)]));
          reg432 <= reg394;
          reg433 <= ({(($signed(reg326) <= (wire203 >> wire198)) ?
                      ($unsigned(reg394) ?
                          (!reg415) : (reg385 ? reg365 : wire197)) : reg322)} ?
              $signed((reg319[(3'h5):(1'h1)] ?
                  (reg306[(1'h1):(1'h1)] ?
                      $signed(reg377) : reg407) : $unsigned((^~wire200)))) : ({(~(wire196 >= wire389))} != $signed(($unsigned(wire198) + (wire197 <<< reg334)))));
        end
      for (forvar434 = (1'h0); (forvar434 < (3'h4)); forvar434 = (forvar434 + (1'h1)))
        begin
          reg435 <= (7'h43);
        end
    end
  assign wire436 = ((reg410[(2'h3):(1'h0)] ?
                           $signed((!{reg325, (8'haf)})) : reg308) ?
                       $signed(reg415) : reg394);
  always
    @(posedge clk) begin
      if (reg290)
        begin
          for (forvar437 = (1'h0); (forvar437 < (2'h3)); forvar437 = (forvar437 + (1'h1)))
            begin
              reg438 = $signed(reg290);
              reg439 <= ({(~&reg379),
                  $signed(($unsigned(reg394) ?
                      (&wire204) : (!reg375)))} != wire284);
              reg440 <= (|(+reg315));
            end
          if ((reg413 ?
              $signed(reg306) : $signed(($signed((~^reg428)) - (reg304 ?
                  (wire203 ? reg432 : wire284) : (+reg366))))))
            begin
              reg441 <= reg325[(3'h4):(2'h2)];
              reg442 = (|(^~(($signed(reg319) | (&reg381)) ?
                  (!(reg412 ?
                      reg438 : reg290)) : ($signed(reg295) ^ reg439[(2'h3):(1'h0)]))));
              reg443 = ((reg347 ~^ (((~|reg433) | $signed((8'hae))) >= (wire436 < (^~reg438)))) >= reg362[(5'h13):(3'h7)]);
              reg444 <= (~^{($unsigned($signed(reg328)) <<< reg325)});
            end
          else
            begin
              reg441 <= $unsigned(((^~reg433[(3'h7):(3'h4)]) <= {$signed(reg440[(2'h2):(1'h1)])}));
              reg444 <= (8'ha2);
              reg445 <= ($unsigned({($unsigned(reg381) <= {wire203,
                          (7'h44)})}) ?
                  (|(~&$signed(reg435[(4'hc):(2'h2)]))) : reg367);
              reg446 = reg439;
              reg447 = ({$signed($signed((wire291 - wire336)))} ?
                  ((((&wire336) >>> $unsigned(wire287)) ^ $unsigned($signed(reg304))) ?
                      (^~((~^reg290) ~^ wire291[(1'h0):(1'h0)])) : $signed(((~&(8'hbc)) != (~^reg410)))) : {reg362[(4'he):(3'h5)],
                      reg375[(1'h1):(1'h0)]});
            end
          reg448 = reg403;
        end
      else
        begin
          if (wire389)
            begin
              reg437 = $signed((-$unsigned(reg407[(4'hf):(3'h6)])));
              reg438 = {reg412};
              reg442 = $unsigned((((|(reg352 >>> reg310)) ?
                  $unsigned(reg396) : $signed($signed(reg442))) - $signed($signed($unsigned(reg410)))));
            end
          else
            begin
              reg439 <= (~$signed($signed(((8'hb5) >= $unsigned((8'h9e))))));
            end
          for (forvar443 = (1'h0); (forvar443 < (1'h0)); forvar443 = (forvar443 + (1'h1)))
            begin
              reg446 = (&reg308[(3'h5):(1'h1)]);
              reg447 = $unsigned($signed(((7'h42) ?
                  {(reg375 * reg352), $unsigned(reg375)} : reg308)));
              reg449 <= $signed((~^($signed(reg391) | ((reg368 ?
                  reg425 : reg390) && $signed(reg437)))));
              reg450 <= (8'hb9);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar451 = (1'h0); (forvar451 < (2'h2)); forvar451 = (forvar451 + (1'h1)))
        begin
          reg452 <= ((~|reg304) ?
              (reg306 != $signed($signed(((7'h48) ?
                  reg345 : reg375)))) : wire291);
          reg453 = (|{(~|reg328[(1'h1):(1'h1)]),
              $signed($unsigned($unsigned(reg301)))});
          for (forvar454 = (1'h0); (forvar454 < (1'h1)); forvar454 = (forvar454 + (1'h1)))
            begin
              reg455 = (-{$unsigned(reg407)});
              reg456 = (!(reg418[(3'h6):(1'h0)] >> {(wire336[(1'h0):(1'h0)] ?
                      $signed(reg391) : (|reg352))}));
              reg457 <= $signed($signed($signed($unsigned(wire203[(4'hb):(2'h2)]))));
              reg458 = ((8'ha8) != ((($signed(reg306) || {reg440, reg298}) ?
                  $unsigned((reg412 ~^ reg326)) : reg390[(1'h0):(1'h0)]) | ((^$signed(reg328)) ?
                  reg325 : reg428)));
            end
          for (forvar459 = (1'h0); (forvar459 < (2'h2)); forvar459 = (forvar459 + (1'h1)))
            begin
              reg460 <= {(~^$signed($unsigned(reg433))),
                  $signed(($signed($unsigned(reg306)) < (reg432 ?
                      (-reg429) : ((8'haa) | reg361))))};
              reg461 = reg450[(3'h7):(2'h3)];
            end
          reg462 <= reg326[(1'h0):(1'h0)];
        end
      if (($signed(({(reg385 ^ wire203)} ?
              $unsigned((reg432 + reg290)) : ($unsigned(wire203) ?
                  $unsigned(wire291) : {reg450}))) ?
          (wire287[(5'h15):(4'he)] != (reg319[(4'hb):(4'h9)] ?
              (+$unsigned(reg365)) : $unsigned($unsigned((8'ha3))))) : (($unsigned($signed(reg304)) && (8'hb1)) + (!$unsigned((8'h9e))))))
        begin
          for (forvar463 = (1'h0); (forvar463 < (1'h0)); forvar463 = (forvar463 + (1'h1)))
            begin
              reg464 = (((8'hb3) ^~ $signed((+{wire197}))) ?
                  $signed($unsigned($signed(((8'hbd) > reg400)))) : (~{reg306}));
              reg465 = reg326[(4'hf):(4'hb)];
              reg466 <= {(($signed(((7'h46) == reg458)) && {((8'h9c) ?
                              reg403 : reg346)}) ?
                      (8'hbd) : forvar463[(1'h0):(1'h0)]),
                  $signed(((7'h47) ?
                      reg306[(1'h0):(1'h0)] : $unsigned({reg366, wire436})))};
              reg467 = (|(8'ha9));
            end
          if ($unsigned($signed($signed(reg385[(3'h4):(1'h1)]))))
            begin
              reg468 = (+reg466[(3'h5):(1'h1)]);
              reg469 <= reg441;
              reg470 <= (reg345[(3'h4):(3'h4)] ?
                  reg462[(5'h13):(4'h9)] : reg457);
              reg471 = (!reg400[(4'he):(1'h0)]);
            end
          else
            begin
              reg469 <= ((((((8'haa) ? (8'hb0) : wire291) ?
                          (~&reg361) : reg445) > $unsigned((wire200 ^ reg415))) ?
                      $unsigned($unsigned($signed(reg418))) : $unsigned($unsigned((reg457 ?
                          (8'had) : reg381)))) ?
                  {(~^$signed($signed(reg308)))} : reg433[(4'hc):(2'h3)]);
              reg470 <= reg303[(1'h0):(1'h0)];
              reg471 = reg428[(5'h11):(4'ha)];
              reg472 = reg435[(1'h1):(1'h1)];
              reg473 <= ((~(($signed(reg452) ?
                      reg315[(1'h0):(1'h0)] : (reg400 * reg322)) || (8'hb5))) ?
                  $unsigned($signed((~^((7'h46) && reg322)))) : {(reg440 ?
                          (~(~^reg452)) : reg439)});
            end
        end
      else
        begin
          for (forvar463 = (1'h0); (forvar463 < (1'h0)); forvar463 = (forvar463 + (1'h1)))
            begin
              reg466 <= $signed((~|(((reg419 != reg375) ?
                  $signed(reg418) : $signed(reg464)) * reg433)));
            end
          if (forvar459)
            begin
              reg467 = $signed($signed(($unsigned({wire286,
                  reg325}) >= (!(+reg390)))));
              reg469 <= $signed(reg439[(3'h7):(2'h3)]);
              reg470 <= ((((((7'h41) && reg381) ?
                          (wire204 ? reg469 : reg413) : (^reg465)) ?
                      $signed($unsigned(reg295)) : ((reg432 <<< reg390) - $unsigned(forvar459))) ?
                  reg441 : ((reg445[(4'hb):(1'h0)] != (reg471 ?
                          reg407 : reg407)) ?
                      reg467[(4'he):(3'h4)] : (|{reg298,
                          reg393}))) || {({(reg464 ^~ reg306),
                          $unsigned(reg415)} ?
                      $signed((reg352 >>> forvar451)) : $unsigned((reg465 + (8'hb5)))),
                  ((-wire336) ? (^~$signed(reg325)) : (|(reg456 < wire389)))});
              reg473 <= {((reg322 != (reg362[(4'ha):(3'h5)] ?
                      (!wire200) : reg361[(3'h4):(3'h4)])) & (reg308[(4'h8):(1'h1)] || $signed($signed(reg431))))};
              reg474 <= $unsigned($unsigned(($unsigned((~^reg464)) > ((reg306 ?
                      (7'h48) : reg403) ?
                  (reg301 ? (8'hb7) : wire203) : {reg465, reg453}))));
            end
          else
            begin
              reg469 <= $signed({(^~(!(reg310 & (8'ha3))))});
            end
          reg475 = {(reg362[(3'h5):(2'h2)] ?
                  (!reg474[(1'h0):(1'h0)]) : (|(~^$signed(reg307)))),
              (8'hb1)};
          reg476 = ({$signed(($signed(reg315) && $signed(reg464))),
                  reg413[(2'h3):(2'h3)]} ?
              reg307 : $unsigned((8'h9f)));
        end
      reg477 <= (~^$signed((^wire196)));
    end
  always
    @(posedge clk) begin
      reg1096 <= reg295[(1'h0):(1'h0)];
      reg1097 <= $signed((reg301[(4'hb):(3'h6)] ?
          wire203[(4'ha):(2'h2)] : {(+wire286[(4'h9):(4'h8)]),
              (wire284 ? $signed(reg361) : reg466)}));
      reg1098 = ((|(&({reg415, (8'ha5)} ~^ {wire436}))) ?
          reg457[(1'h0):(1'h0)] : {($unsigned((+(7'h48))) <= reg445),
              $unsigned((reg379[(1'h1):(1'h0)] <= (reg441 ?
                  reg346 : reg403)))});
      if ($unsigned({((!reg1097[(3'h7):(1'h0)]) ?
              ({(8'ha6), reg410} ?
                  (&wire203) : {reg307}) : reg394[(2'h2):(1'h1)]),
          ((^~reg470) ? reg450 : ($signed((8'h9f)) < wire199[(4'he):(4'hd)]))}))
        begin
          reg1099 <= (($unsigned(($signed(reg362) ?
                  reg393[(4'hd):(4'h9)] : ((7'h40) ? wire1094 : reg469))) ?
              $unsigned(((^~(8'hb1)) ?
                  (reg413 ?
                      reg367 : (8'h9e)) : (reg441 | reg466))) : ($signed((wire284 > reg412)) ?
                  (wire199 ^ reg429) : (~^{wire1094, reg433}))) || (8'hbe));
          reg1100 = $unsigned((-reg412));
          for (forvar1101 = (1'h0); (forvar1101 < (2'h3)); forvar1101 = (forvar1101 + (1'h1)))
            begin
              reg1102 <= $signed(((!(wire287[(4'h8):(4'h8)] | $signed(reg1099))) != reg449[(3'h6):(2'h3)]));
            end
          for (forvar1103 = (1'h0); (forvar1103 < (3'h4)); forvar1103 = (forvar1103 + (1'h1)))
            begin
              reg1104 <= ($signed(wire389) ?
                  reg412[(5'h15):(1'h0)] : $signed(((reg418[(3'h4):(2'h3)] ?
                      reg327[(4'ha):(4'ha)] : $signed(reg345)) || wire198[(2'h3):(1'h0)])));
            end
          reg1105 = ((&(^~$unsigned((wire204 << reg474)))) >>> $unsigned($signed($signed(reg470[(2'h3):(2'h3)]))));
        end
      else
        begin
          for (forvar1099 = (1'h0); (forvar1099 < (1'h1)); forvar1099 = (forvar1099 + (1'h1)))
            begin
              reg1101 <= $unsigned(reg326);
            end
          for (forvar1102 = (1'h0); (forvar1102 < (1'h1)); forvar1102 = (forvar1102 + (1'h1)))
            begin
              reg1103 = wire198;
              reg1104 <= {wire199[(5'h13):(4'h8)]};
              reg1105 = ((8'hb7) + {$signed($signed($signed(reg413)))});
              reg1106 = reg419;
            end
          if ({((reg1097 && $signed($unsigned((8'hb6)))) ^ (|$unsigned(reg385))),
              reg333[(1'h1):(1'h0)]})
            begin
              reg1107 = $unsigned((-reg380[(4'ha):(4'h8)]));
              reg1108 <= reg428;
              reg1109 <= $signed(($signed(((wire198 ? reg334 : (8'h9d)) ?
                      $signed(reg452) : $unsigned(reg327))) ?
                  reg413 : reg1097[(4'h8):(1'h1)]));
            end
          else
            begin
              reg1107 = $unsigned(reg385);
              reg1110 = ((~$signed(reg1109[(4'hc):(3'h5)])) ?
                  $unsigned((~$unsigned(((8'ha8) - reg394)))) : reg374[(4'hb):(3'h7)]);
              reg1111 = (+(((+$unsigned(wire199)) >>> (~&(reg431 ?
                  (7'h49) : reg441))) + $unsigned(reg409[(1'h0):(1'h0)])));
              reg1112 = reg396[(4'hd):(2'h3)];
              reg1113 = (7'h42);
            end
        end
    end
  always
    @(posedge clk) begin
      if (wire389[(1'h0):(1'h0)])
        begin
          if ($unsigned((~^({(reg398 ? wire1094 : wire284)} ?
              (((8'hb2) ? reg435 : reg290) ?
                  $unsigned(reg394) : (^wire336)) : {(~|(8'h9e)), reg390}))))
            begin
              reg1114 <= $unsigned($unsigned($unsigned((reg407 ?
                  wire287[(2'h2):(2'h2)] : (-reg377)))));
            end
          else
            begin
              reg1115 = $unsigned({$unsigned($signed((reg328 - reg1099)))});
            end
          reg1116 = (~|(8'hb7));
          reg1117 <= wire287[(4'ha):(2'h3)];
          reg1118 <= (reg435 >> (~&$signed((+(reg374 >> reg445)))));
        end
      else
        begin
          if (((reg413[(1'h0):(1'h0)] ?
              wire198 : $signed(($unsigned(reg375) << (reg429 != (8'hac))))) << reg333))
            begin
              reg1114 <= (~|$unsigned(reg449));
            end
          else
            begin
              reg1114 <= (+reg1102);
              reg1117 <= reg380;
            end
          reg1119 = (wire287[(2'h3):(2'h3)] | {($signed({reg466}) * $signed(((8'hbf) & reg380)))});
          reg1120 = {($signed(((-(8'h9f)) ?
                      $signed(reg367) : $unsigned(reg452))) ?
                  (($signed(reg460) >= (~reg412)) ?
                      (^(reg412 ?
                          reg368 : wire291)) : (-wire286[(3'h7):(3'h5)])) : (7'h42))};
        end
      reg1121 <= (reg327[(4'hf):(3'h6)] ? ((!reg457) >= reg418) : reg470);
      for (forvar1122 = (1'h0); (forvar1122 < (2'h3)); forvar1122 = (forvar1122 + (1'h1)))
        begin
          for (forvar1123 = (1'h0); (forvar1123 < (2'h3)); forvar1123 = (forvar1123 + (1'h1)))
            begin
              reg1124 <= $signed(($unsigned((~|(reg439 && reg1120))) <<< (reg352 ?
                  $signed(reg396) : (~|(~&(8'hb7))))));
              reg1125 = $unsigned({{(&(reg315 ? (8'hae) : reg477))},
                  $signed($signed($signed((8'hbe))))});
              reg1126 <= wire389[(3'h5):(2'h2)];
            end
          if ({$signed($unsigned($signed((!(7'h42)))))})
            begin
              reg1127 <= (^reg334);
              reg1128 = $signed((reg1120[(4'hf):(4'hd)] ?
                  {(~&{wire287, reg1102}),
                      reg307[(2'h3):(1'h1)]} : $unsigned((+(-reg298)))));
            end
          else
            begin
              reg1127 <= {(8'hac)};
              reg1128 = (~&reg1128);
              reg1129 = reg1116[(1'h0):(1'h0)];
            end
          reg1130 <= $unsigned(wire286);
          for (forvar1131 = (1'h0); (forvar1131 < (1'h0)); forvar1131 = (forvar1131 + (1'h1)))
            begin
              reg1132 <= $signed((((^reg1108) ?
                  $unsigned(reg375[(4'hd):(4'h9)]) : reg294[(1'h0):(1'h0)]) <<< $signed($signed((~&reg1116)))));
              reg1133 = (|(&reg322[(4'hd):(1'h1)]));
            end
          for (forvar1134 = (1'h0); (forvar1134 < (3'h4)); forvar1134 = (forvar1134 + (1'h1)))
            begin
              reg1135 <= (reg1119[(4'h9):(2'h2)] ?
                  ((8'hb7) | $signed(((8'hb5) ^ ((8'hbd) & reg1126)))) : reg368[(4'hf):(4'hb)]);
            end
        end
      if (reg1101)
        begin
          reg1136 <= $signed($signed(reg377));
          for (forvar1137 = (1'h0); (forvar1137 < (2'h2)); forvar1137 = (forvar1137 + (1'h1)))
            begin
              reg1138 <= $signed(reg391[(4'ha):(4'h9)]);
              reg1139 <= ((~^(^{reg326[(5'h10):(3'h4)],
                  {reg1114, reg347}})) ~^ ((reg1120 != ($signed(reg325) ?
                  (reg469 ? reg301 : reg377) : $signed((8'ha1)))) >= (wire199 ?
                  ((8'ha1) | reg347[(5'h10):(5'h10)]) : $signed(forvar1122[(3'h7):(2'h2)]))));
              reg1140 = forvar1123[(3'h4):(1'h1)];
              reg1141 <= (^reg380[(4'hf):(3'h4)]);
              reg1142 <= $unsigned($unsigned((reg298[(1'h1):(1'h0)] ?
                  reg445 : reg1115[(3'h6):(1'h1)])));
            end
          for (forvar1143 = (1'h0); (forvar1143 < (2'h2)); forvar1143 = (forvar1143 + (1'h1)))
            begin
              reg1144 = reg374;
              reg1145 = (reg1118 == $signed(reg377));
              reg1146 <= (^~$signed((+((forvar1123 & reg1140) ?
                  (8'hb1) : $signed(reg462)))));
              reg1147 = ($unsigned((~&$signed(reg410))) ?
                  reg1120[(4'hf):(4'h8)] : (^~(reg294[(3'h7):(3'h6)] ?
                      reg409 : $unsigned($signed(reg377)))));
            end
          reg1148 <= $unsigned(reg362);
          if ($signed((^$unsigned((8'ha0)))))
            begin
              reg1149 <= reg466[(3'h5):(1'h0)];
              reg1150 <= $unsigned(($unsigned({$signed(reg1130)}) != ((((8'hb4) & (7'h47)) ?
                      {reg415, (8'haa)} : {reg457}) ?
                  $unsigned(forvar1123) : (reg394 >> $signed((7'h4a))))));
              reg1151 <= $signed(reg1127[(1'h0):(1'h0)]);
            end
          else
            begin
              reg1149 <= wire291;
              reg1150 <= reg317;
              reg1151 <= (7'h40);
              reg1152 <= $signed((($signed(reg374) ~^ (((8'hbf) * reg1145) ?
                  (+reg365) : (wire436 ?
                      reg381 : reg1129))) < $unsigned((^$signed(reg1128)))));
              reg1153 <= ($unsigned({$unsigned(reg1145)}) * $signed(reg327));
            end
        end
      else
        begin
          reg1136 <= $signed(reg398);
          reg1137 <= $signed($signed(reg327));
        end
    end
endmodule
