(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param1768 = ((~{(((7'h46) ? (8'ha1) : (8'ha7)) ? (~|(8'h9f)) : ((7'h4a) ^~ (8'hae)))}) ? ((-(&((8'hb5) == (8'haf)))) & (!(-(|(7'h46))))) : ({((~&(7'h43)) ? (^~(8'hbc)) : ((8'hb9) != (8'hb3))), {(~(7'h48)), ((7'h42) ? (7'h42) : (8'hb1))}} >>> ((~{(8'hb9)}) ? ((8'haa) >>> ((7'h42) ? (8'hb0) : (7'h44))) : (&(~(7'h40)))))))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h75e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire3;
  input wire [(5'h18):(1'h0)] wire2;
  input wire [(2'h3):(1'h0)] wire1;
  input wire [(3'h6):(1'h0)] wire0;
  wire signed [(4'h9):(1'h0)] wire1720;
  wire [(4'hf):(1'h0)] wire77;
  wire signed [(5'h12):(1'h0)] wire32;
  reg [(3'h6):(1'h0)] reg1767 = (1'h0);
  reg [(4'he):(1'h0)] reg1766 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1763 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1761 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1760 = (1'h0);
  reg [(4'h9):(1'h0)] reg1750 = (1'h0);
  reg [(3'h6):(1'h0)] reg1757 = (1'h0);
  reg [(2'h2):(1'h0)] reg1754 = (1'h0);
  reg [(5'h13):(1'h0)] reg1753 = (1'h0);
  reg [(4'hd):(1'h0)] reg1752 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1747 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1744 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1743 = (1'h0);
  reg [(4'h9):(1'h0)] reg1740 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1738 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1737 = (1'h0);
  reg [(5'h18):(1'h0)] reg1736 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1734 = (1'h0);
  reg [(5'h14):(1'h0)] reg1733 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1732 = (1'h0);
  reg [(3'h7):(1'h0)] reg1727 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg93 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg92 = (1'h0);
  reg [(5'h11):(1'h0)] reg91 = (1'h0);
  reg [(5'h17):(1'h0)] reg87 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg83 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg82 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg76 = (1'h0);
  reg [(4'h8):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg74 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg67 = (1'h0);
  reg [(5'h12):(1'h0)] reg66 = (1'h0);
  reg [(4'he):(1'h0)] reg58 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg56 = (1'h0);
  reg [(5'h13):(1'h0)] reg54 = (1'h0);
  reg [(5'h12):(1'h0)] reg53 = (1'h0);
  reg [(4'ha):(1'h0)] reg47 = (1'h0);
  reg [(4'h9):(1'h0)] reg43 = (1'h0);
  reg [(3'h6):(1'h0)] reg41 = (1'h0);
  reg [(5'h14):(1'h0)] reg38 = (1'h0);
  reg [(4'h8):(1'h0)] reg36 = (1'h0);
  reg [(5'h13):(1'h0)] reg35 = (1'h0);
  reg [(5'h13):(1'h0)] reg34 = (1'h0);
  reg [(4'h8):(1'h0)] reg29 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg28 = (1'h0);
  reg [(2'h2):(1'h0)] reg24 = (1'h0);
  reg [(4'hd):(1'h0)] reg23 = (1'h0);
  reg signed [(4'he):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg15 = (1'h0);
  reg [(2'h3):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg11 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg9 = (1'h0);
  reg [(5'h11):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1765 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1764 = (1'h0);
  reg [(5'h11):(1'h0)] reg1762 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1759 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1758 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1756 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1755 = (1'h0);
  reg [(3'h6):(1'h0)] reg1751 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1750 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1749 = (1'h0);
  reg [(4'h9):(1'h0)] reg1748 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1746 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1745 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1742 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1741 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1739 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1735 = (1'h0);
  reg [(5'h13):(1'h0)] reg1735 = (1'h0);
  reg [(4'hf):(1'h0)] reg1731 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1730 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1729 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1728 = (1'h0);
  reg [(5'h12):(1'h0)] reg1726 = (1'h0);
  reg [(5'h18):(1'h0)] reg1725 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1724 = (1'h0);
  reg [(5'h13):(1'h0)] reg1723 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1722 = (1'h0);
  reg [(5'h17):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg90 = (1'h0);
  reg [(5'h12):(1'h0)] forvar89 = (1'h0);
  reg [(5'h17):(1'h0)] reg88 = (1'h0);
  reg signed [(4'he):(1'h0)] reg86 = (1'h0);
  reg [(5'h16):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar83 = (1'h0);
  reg [(4'h8):(1'h0)] reg78 = (1'h0);
  reg [(4'hd):(1'h0)] reg84 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg81 = (1'h0);
  reg [(3'h6):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg79 = (1'h0);
  reg [(5'h18):(1'h0)] forvar78 = (1'h0);
  reg [(5'h18):(1'h0)] reg72 = (1'h0);
  reg [(5'h14):(1'h0)] reg71 = (1'h0);
  reg [(4'hb):(1'h0)] reg70 = (1'h0);
  reg [(5'h12):(1'h0)] reg69 = (1'h0);
  reg [(5'h11):(1'h0)] reg68 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg65 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg64 = (1'h0);
  reg [(4'hc):(1'h0)] reg63 = (1'h0);
  reg [(4'hd):(1'h0)] reg62 = (1'h0);
  reg [(2'h3):(1'h0)] reg61 = (1'h0);
  reg [(4'he):(1'h0)] forvar60 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar59 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg57 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg55 = (1'h0);
  reg [(4'hb):(1'h0)] reg52 = (1'h0);
  reg [(4'h9):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar50 = (1'h0);
  reg [(5'h12):(1'h0)] reg49 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg48 = (1'h0);
  reg [(3'h5):(1'h0)] reg46 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar45 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar44 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar42 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg40 = (1'h0);
  reg [(2'h3):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg37 = (1'h0);
  reg [(5'h10):(1'h0)] forvar33 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg31 = (1'h0);
  reg [(4'hc):(1'h0)] reg30 = (1'h0);
  reg [(5'h16):(1'h0)] reg27 = (1'h0);
  reg [(4'h8):(1'h0)] reg26 = (1'h0);
  reg [(4'h9):(1'h0)] reg25 = (1'h0);
  reg [(5'h13):(1'h0)] forvar22 = (1'h0);
  reg [(4'hf):(1'h0)] reg21 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg20 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg18 = (1'h0);
  reg [(5'h17):(1'h0)] forvar17 = (1'h0);
  reg [(3'h6):(1'h0)] reg16 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4 = (1'h0);
  assign y = {wire1720,
                 wire77,
                 wire32,
                 reg1767,
                 reg1766,
                 reg1763,
                 reg1761,
                 reg1760,
                 reg1750,
                 reg1757,
                 reg1754,
                 reg1753,
                 reg1752,
                 reg1747,
                 reg1744,
                 reg1743,
                 reg1740,
                 reg1738,
                 reg1737,
                 reg1736,
                 reg1734,
                 reg1733,
                 reg1732,
                 reg1727,
                 reg93,
                 reg92,
                 reg91,
                 reg87,
                 reg83,
                 reg82,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg67,
                 reg66,
                 reg58,
                 reg56,
                 reg54,
                 reg53,
                 reg47,
                 reg43,
                 reg41,
                 reg38,
                 reg36,
                 reg35,
                 reg34,
                 reg29,
                 reg28,
                 reg24,
                 reg23,
                 reg17,
                 reg15,
                 reg14,
                 reg13,
                 reg11,
                 reg9,
                 reg8,
                 reg1765,
                 forvar1764,
                 reg1762,
                 forvar1759,
                 forvar1758,
                 forvar1756,
                 reg1755,
                 reg1751,
                 forvar1750,
                 reg1749,
                 reg1748,
                 reg1746,
                 reg1745,
                 reg1742,
                 reg1741,
                 reg1739,
                 forvar1735,
                 reg1735,
                 reg1731,
                 reg1730,
                 forvar1729,
                 reg1728,
                 reg1726,
                 reg1725,
                 reg1724,
                 reg1723,
                 forvar1722,
                 reg94,
                 reg90,
                 forvar89,
                 reg88,
                 reg86,
                 reg85,
                 forvar83,
                 reg78,
                 reg84,
                 reg81,
                 reg80,
                 reg79,
                 forvar78,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 forvar60,
                 forvar59,
                 reg57,
                 reg55,
                 reg52,
                 reg51,
                 forvar50,
                 reg49,
                 reg48,
                 reg46,
                 forvar45,
                 forvar44,
                 forvar42,
                 reg40,
                 reg39,
                 reg37,
                 forvar33,
                 reg31,
                 reg30,
                 reg27,
                 reg26,
                 reg25,
                 forvar22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 forvar17,
                 reg16,
                 reg12,
                 reg10,
                 forvar7,
                 reg6,
                 reg5,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (1'h0)); forvar4 = (forvar4 + (1'h1)))
        begin
          reg5 = wire0[(3'h4):(2'h3)];
          reg6 = wire0[(3'h5):(1'h1)];
        end
      for (forvar7 = (1'h0); (forvar7 < (2'h2)); forvar7 = (forvar7 + (1'h1)))
        begin
          reg8 <= $signed(reg5[(2'h3):(1'h0)]);
          reg9 <= $signed(wire1[(1'h1):(1'h1)]);
          reg10 = ($signed($signed(reg9)) >= (reg6[(3'h6):(3'h6)] > wire2[(5'h15):(4'hd)]));
          reg11 <= $unsigned(((wire1 ?
              (^(reg8 && forvar7)) : ((wire3 ? (7'h46) : forvar7) ?
                  (forvar7 ?
                      wire0 : wire3) : ((8'ha1) || (8'ha2)))) >= (+{$unsigned(wire3)})));
          if (reg11[(4'hc):(3'h7)])
            begin
              reg12 = ($unsigned(wire2[(5'h14):(1'h1)]) ? (+(&reg9)) : reg5);
            end
          else
            begin
              reg13 <= wire1[(1'h0):(1'h0)];
              reg14 <= ({wire2[(3'h7):(3'h6)], {$signed((wire2 ^ reg8))}} ?
                  reg8 : $unsigned(reg11[(3'h4):(3'h4)]));
              reg15 <= (($signed((&(reg5 ? reg5 : reg12))) ? forvar4 : reg14) ?
                  ((8'hb0) || $signed((!(-forvar4)))) : $unsigned(reg13[(1'h0):(1'h0)]));
              reg16 = {$signed($signed((~&$signed(reg14))))};
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg14[(2'h2):(1'h1)])
        begin
          reg17 <= wire2[(3'h6):(2'h3)];
        end
      else
        begin
          for (forvar17 = (1'h0); (forvar17 < (1'h1)); forvar17 = (forvar17 + (1'h1)))
            begin
              reg18 = $unsigned(($unsigned(reg17[(4'hd):(3'h6)]) ?
                  (reg15 < ({reg13,
                      wire0} & (~^wire1))) : $signed((^(wire0 ^ wire3)))));
              reg19 = wire2[(4'hd):(3'h6)];
              reg20 = (($unsigned((~^$signed(reg8))) ?
                  (wire0[(2'h2):(1'h0)] ?
                      (~$unsigned(reg9)) : $unsigned((&(8'hbd)))) : $unsigned(reg8[(4'he):(4'hc)])) << (+reg9[(1'h1):(1'h1)]));
              reg21 = wire3[(2'h2):(1'h1)];
            end
          for (forvar22 = (1'h0); (forvar22 < (1'h0)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 <= reg20;
              reg24 <= $unsigned((!$unsigned($signed((8'hbd)))));
              reg25 = $unsigned($signed(reg21));
              reg26 = $unsigned((^~$unsigned((8'h9d))));
              reg27 = $unsigned($signed(((+$signed((7'h48))) >= {(wire3 ^ reg20),
                  {(8'hb6), wire0}})));
            end
          reg28 <= reg13[(1'h1):(1'h1)];
          if ((|$unsigned($signed(reg14))))
            begin
              reg29 <= ($signed($unsigned((reg19[(4'hb):(4'hb)] >> (reg25 ?
                      reg20 : reg11)))) ?
                  $unsigned(wire1) : {$unsigned(reg24), reg25});
            end
          else
            begin
              reg30 = (reg15[(5'h16):(2'h3)] >> (^~{forvar17}));
            end
        end
      reg31 = ($unsigned($signed(reg30[(4'hb):(1'h0)])) ?
          $signed((~|$unsigned($signed(reg25)))) : reg17);
    end
  assign wire32 = reg11[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar33 = (1'h0); (forvar33 < (1'h0)); forvar33 = (forvar33 + (1'h1)))
        begin
          if (reg17[(4'hb):(4'h8)])
            begin
              reg34 <= reg23[(1'h1):(1'h1)];
              reg35 <= $unsigned(($signed(reg24[(1'h1):(1'h0)]) ?
                  (|$signed($signed(reg9))) : $signed(wire3)));
              reg36 <= (($unsigned(reg23[(3'h6):(3'h4)]) < (($signed(reg34) ?
                  (reg29 ?
                      reg14 : forvar33) : $signed(wire3)) >> $unsigned((forvar33 < reg14)))) << wire3);
              reg37 = (reg11 && {$signed((~&(~|reg13))),
                  (((reg11 >> reg29) ? (reg17 >> reg23) : {reg24, (8'hbf)}) ?
                      reg14 : (reg28[(3'h5):(3'h4)] ?
                          wire3[(1'h0):(1'h0)] : {(7'h42)}))});
              reg38 <= $signed(((&reg13[(1'h0):(1'h0)]) >= reg17[(3'h5):(3'h4)]));
            end
          else
            begin
              reg34 <= $unsigned({(-wire0[(2'h2):(1'h1)]),
                  $signed((-(!wire2)))});
              reg37 = $unsigned(reg17);
              reg38 <= (&$signed((reg28[(3'h5):(1'h0)] ?
                  reg35 : $signed($signed(reg8)))));
              reg39 = ({$unsigned(($unsigned((7'h43)) ? (~^wire32) : reg29))} ?
                  wire2[(4'he):(2'h3)] : reg15[(4'hd):(3'h6)]);
            end
          reg40 = $unsigned($signed(reg14[(2'h3):(1'h1)]));
        end
      reg41 <= reg38[(5'h11):(5'h10)];
      for (forvar42 = (1'h0); (forvar42 < (1'h0)); forvar42 = (forvar42 + (1'h1)))
        begin
          reg43 <= ($unsigned((~|$unsigned((7'h41)))) - {reg13,
              $signed(((^reg28) ? forvar42 : $signed((7'h47))))});
        end
    end
  always
    @(posedge clk) begin
      for (forvar44 = (1'h0); (forvar44 < (2'h2)); forvar44 = (forvar44 + (1'h1)))
        begin
          for (forvar45 = (1'h0); (forvar45 < (2'h3)); forvar45 = (forvar45 + (1'h1)))
            begin
              reg46 = $unsigned(((8'haf) ?
                  ((!reg9[(1'h1):(1'h1)]) ?
                      (+$signed((8'hb6))) : ((reg9 ^~ reg41) ?
                          $signed(wire1) : reg28[(3'h5):(2'h2)])) : $unsigned((((8'hb6) ?
                      wire0 : reg11) != (^reg38)))));
              reg47 <= reg28;
              reg48 = ((|((|(reg41 ^~ wire32)) ?
                  ($signed((8'hb9)) ?
                      $unsigned((7'h42)) : (wire0 == reg9)) : wire1[(1'h0):(1'h0)])) ^~ reg41[(1'h0):(1'h0)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg49 = (&({$unsigned(((8'hb8) ? wire1 : reg35)), $unsigned((|(8'hbd)))} ?
          ($signed($signed(reg28)) ?
              {reg14, reg23} : ($unsigned(reg43) ?
                  (reg9 | reg9) : (~reg23))) : (wire32[(1'h0):(1'h0)] ?
              reg17[(4'hd):(4'hc)] : $signed(reg29[(2'h2):(1'h0)]))));
      for (forvar50 = (1'h0); (forvar50 < (2'h3)); forvar50 = (forvar50 + (1'h1)))
        begin
          if ((!((reg23 ? reg23[(1'h0):(1'h0)] : reg11[(4'ha):(1'h1)]) ?
              (!reg13) : (wire0 == (reg49[(4'h9):(4'h9)] | reg11)))))
            begin
              reg51 = $signed(wire1[(1'h0):(1'h0)]);
              reg52 = (reg14 * (!(reg38[(3'h4):(2'h3)] >>> (-(~^reg28)))));
              reg53 <= $unsigned(wire3[(1'h1):(1'h0)]);
              reg54 <= ((reg13 ?
                  (reg35 ?
                      $signed(wire32[(4'h9):(1'h1)]) : $unsigned($unsigned((7'h45)))) : (8'hb2)) <= (reg13[(1'h1):(1'h1)] < ((((8'ha3) ?
                  (8'hb0) : wire0) >>> reg29) ~^ (^~$signed((8'hac))))));
              reg55 = (((7'h45) < reg28[(4'h9):(1'h1)]) ~^ $unsigned(reg14[(2'h2):(1'h0)]));
            end
          else
            begin
              reg53 <= reg51;
              reg55 = $signed(({{wire32[(4'h9):(2'h3)], $signed(reg13)},
                      reg29} ?
                  $unsigned($unsigned((wire2 >> wire3))) : wire2));
              reg56 <= $signed(((reg17 ?
                      reg34[(1'h1):(1'h0)] : $unsigned((-reg38))) ?
                  (((reg47 <= (8'h9e)) + (&reg28)) + $unsigned((reg49 ?
                      reg24 : forvar50))) : (|((reg38 ?
                      reg47 : reg9) == (!reg11)))));
              reg57 = reg17;
            end
          reg58 <= (|(~^($signed(reg43) && (8'h9c))));
        end
      for (forvar59 = (1'h0); (forvar59 < (3'h4)); forvar59 = (forvar59 + (1'h1)))
        begin
          for (forvar60 = (1'h0); (forvar60 < (2'h2)); forvar60 = (forvar60 + (1'h1)))
            begin
              reg61 = (8'hab);
            end
          reg62 = ($unsigned((~&(-$unsigned(reg52)))) || ({wire0} ?
              reg55 : reg49[(4'he):(4'hb)]));
          if ($unsigned($unsigned((~&{(reg52 ? reg28 : reg24)}))))
            begin
              reg63 = {$unsigned(wire3)};
              reg64 = ((((forvar50 ? reg29 : (7'h41)) >= (~(reg29 ?
                      reg51 : (8'hbd)))) ?
                  reg29[(3'h5):(1'h0)] : $signed(wire32[(4'hd):(4'hb)])) ^~ ((~^$signed((reg34 + forvar50))) ?
                  reg23 : (((~^reg51) << {(8'hae)}) ?
                      $unsigned(reg43[(3'h4):(3'h4)]) : $unsigned(reg51[(3'h4):(2'h2)]))));
              reg65 = (reg41 <<< (~|(!$unsigned(wire3))));
            end
          else
            begin
              reg66 <= reg53;
              reg67 <= reg24[(1'h1):(1'h1)];
              reg68 = ($signed(wire1[(1'h0):(1'h0)]) ? reg11 : $signed(reg62));
            end
          reg69 = ({$unsigned(((^~reg11) ?
                  (reg34 ? reg62 : reg63) : (reg17 ?
                      reg41 : (8'h9d))))} > $signed((reg63 ?
              reg67[(2'h2):(1'h0)] : $signed($unsigned(reg58)))));
          if (((~(+forvar50[(3'h4):(3'h4)])) ?
              $signed(reg54[(3'h4):(2'h2)]) : {$unsigned($unsigned(reg55))}))
            begin
              reg70 = (reg43 ?
                  ((^~((reg41 ? reg62 : reg66) ?
                      $unsigned(wire1) : reg11[(3'h4):(2'h3)])) - $unsigned({wire2[(3'h4):(1'h0)],
                      (reg41 ? (8'hb7) : reg66)})) : reg64);
              reg71 = (wire2[(1'h1):(1'h1)] ?
                  $signed((wire32 ~^ $signed(wire3))) : (~($unsigned($signed(reg49)) ^~ $signed({reg47,
                      (8'hb7)}))));
              reg72 = reg43[(1'h1):(1'h0)];
              reg73 <= reg70;
            end
          else
            begin
              reg73 <= (($unsigned($signed((8'ha6))) ?
                      reg23[(2'h2):(2'h2)] : $signed((~^(7'h46)))) ?
                  {reg9} : reg67[(4'h9):(1'h1)]);
              reg74 <= $signed((&$unsigned(reg53)));
              reg75 <= ($unsigned($signed($signed($unsigned(reg24)))) ?
                  wire1[(1'h1):(1'h1)] : (^~$signed($unsigned($signed((8'ha9))))));
            end
        end
      reg76 <= ((({reg53} ?
                  $unsigned($signed(reg14)) : ((reg53 & reg65) ?
                      reg34[(5'h11):(4'he)] : $signed((7'h41)))) ?
              $unsigned(forvar60[(3'h6):(1'h0)]) : {(-$unsigned(wire3))}) ?
          ((^~($unsigned(reg74) * (~&reg14))) + (+reg56[(4'hf):(1'h1)])) : $signed($signed(wire3[(1'h0):(1'h0)])));
    end
  assign wire77 = ($signed($unsigned($signed($signed(reg35)))) >>> reg75[(2'h3):(1'h0)]);
  always
    @(posedge clk) begin
      if (reg47)
        begin
          for (forvar78 = (1'h0); (forvar78 < (1'h0)); forvar78 = (forvar78 + (1'h1)))
            begin
              reg79 = {$signed(((~^(reg58 ? wire1 : reg41)) ?
                      reg13[(1'h1):(1'h1)] : reg13[(3'h5):(3'h5)]))};
              reg80 = reg11[(3'h6):(1'h1)];
            end
          if (((forvar78[(4'h8):(2'h3)] ?
              $signed($signed((^~forvar78))) : (((&reg9) ?
                      wire0 : ((8'hb1) ? reg73 : reg56)) ?
                  (reg43[(3'h4):(2'h2)] == reg76[(3'h5):(3'h4)]) : {(^reg56),
                      (|reg73)})) & $signed($unsigned((reg80[(3'h4):(1'h1)] ?
              $unsigned((8'hba)) : (~^reg56))))))
            begin
              reg81 = ((reg58[(1'h1):(1'h1)] ?
                      ((((8'hac) ? reg56 : reg67) & {reg54,
                          reg58}) & reg58) : reg54) ?
                  (!$unsigned(($signed(reg53) ?
                      (wire1 ?
                          reg11 : reg41) : (~(8'h9c))))) : {(-reg34[(5'h13):(3'h5)])});
              reg82 <= ((&($signed($unsigned(reg79)) <= reg11[(4'hf):(2'h3)])) || (reg41 ?
                  ((+$signed(wire77)) ?
                      (reg38[(3'h7):(3'h4)] == $unsigned(wire3)) : $unsigned($signed(reg17))) : (^$signed(reg54[(2'h3):(1'h1)]))));
              reg83 <= (!reg28);
            end
          else
            begin
              reg81 = $signed((reg80[(1'h0):(1'h0)] ?
                  (^~$signed((wire2 - reg11))) : $signed($signed({reg73}))));
              reg84 = wire77;
            end
        end
      else
        begin
          if (reg17[(4'ha):(2'h2)])
            begin
              reg78 = (~^{reg76, (7'h49)});
              reg79 = ($unsigned(reg8) ?
                  ($unsigned((((8'hbd) ? wire0 : reg58) ?
                          reg29[(3'h7):(1'h0)] : (reg43 ? reg47 : reg34))) ?
                      reg41[(2'h3):(1'h1)] : reg29[(3'h7):(1'h1)]) : ($unsigned(reg24[(1'h1):(1'h0)]) + $signed(forvar78[(4'hf):(4'hd)])));
            end
          else
            begin
              reg78 = reg54;
              reg79 = (reg8 ?
                  $signed($unsigned($signed($unsigned(reg23)))) : (reg41[(3'h6):(1'h0)] ?
                      {{$signed(reg17), reg15}, reg82} : $unsigned(reg56)));
              reg82 <= reg9;
            end
          for (forvar83 = (1'h0); (forvar83 < (2'h2)); forvar83 = (forvar83 + (1'h1)))
            begin
              reg84 = $signed(reg38);
            end
          reg85 = $unsigned(reg58[(2'h2):(2'h2)]);
        end
      reg86 = $unsigned(reg53[(3'h6):(1'h0)]);
      reg87 <= (!reg9);
      reg88 = reg85;
    end
  always
    @(posedge clk) begin
      for (forvar89 = (1'h0); (forvar89 < (3'h4)); forvar89 = (forvar89 + (1'h1)))
        begin
          reg90 = (8'hba);
        end
      reg91 <= (reg24[(1'h0):(1'h0)] ?
          {$unsigned($signed({reg66}))} : ((!(^~$unsigned(reg56))) ?
              ((reg43[(3'h5):(1'h1)] && $signed(reg47)) <<< $signed(wire3)) : (|(forvar89 ?
                  $signed(reg28) : wire1[(1'h1):(1'h0)]))));
      reg92 <= (|(8'hbd));
      reg93 <= reg92;
      reg94 = $signed(wire32);
    end
  module95 #() modinst1721 (wire1720, clk, reg83, reg54, reg73, reg38);
  always
    @(posedge clk) begin
      for (forvar1722 = (1'h0); (forvar1722 < (3'h4)); forvar1722 = (forvar1722 + (1'h1)))
        begin
          if ((7'h43))
            begin
              reg1723 = ((8'hb5) >> {wire77});
              reg1724 = reg41[(1'h0):(1'h0)];
              reg1725 = (|reg82[(1'h1):(1'h0)]);
              reg1726 = $signed({$signed((reg36[(3'h6):(3'h4)] ?
                      reg82[(1'h0):(1'h0)] : {reg17}))});
              reg1727 <= (+((-((reg91 | (8'h9e)) <= (reg76 != reg35))) ^ $unsigned((&(reg13 > reg83)))));
            end
          else
            begin
              reg1727 <= ((~&(!reg15[(3'h4):(1'h1)])) & $signed(wire3));
              reg1728 = $signed($unsigned((reg91 > (+(reg11 ?
                  reg56 : reg54)))));
            end
          for (forvar1729 = (1'h0); (forvar1729 < (1'h1)); forvar1729 = (forvar1729 + (1'h1)))
            begin
              reg1730 = forvar1722[(2'h2):(1'h1)];
              reg1731 = (($signed($signed(reg74)) ? (~|(~^reg29)) : (8'hb5)) ?
                  ((!(reg76[(2'h2):(1'h1)] ?
                          reg92 : ((7'h41) ? reg43 : forvar1729))) ?
                      reg66[(4'h9):(3'h4)] : (+(+(reg24 || reg13)))) : ($signed({$unsigned(reg47)}) ~^ $unsigned((^~reg75[(4'h8):(2'h2)]))));
              reg1732 <= $signed((8'hab));
            end
        end
      reg1733 <= (-reg36);
      reg1734 <= wire1720;
      if ($signed($signed({({reg1725} != (reg1730 ? reg58 : wire32)),
          $unsigned(reg93[(2'h2):(1'h1)])})))
        begin
          if ($signed(($unsigned($signed($unsigned(reg82))) < $unsigned((~&(reg13 >= (7'h43)))))))
            begin
              reg1735 = reg1728[(3'h4):(1'h0)];
            end
          else
            begin
              reg1735 = ({($unsigned((^~reg47)) > ($signed((8'hbd)) & $signed(reg35)))} ^~ (~&$signed((^~reg1734))));
              reg1736 <= $unsigned(((~reg93) ?
                  reg56 : (reg8[(4'hf):(4'he)] >= ((reg8 ?
                      wire0 : (8'hbb)) <= ((7'h4a) <= wire2)))));
              reg1737 <= (|reg15[(5'h12):(5'h11)]);
              reg1738 <= (7'h44);
            end
        end
      else
        begin
          for (forvar1735 = (1'h0); (forvar1735 < (1'h0)); forvar1735 = (forvar1735 + (1'h1)))
            begin
              reg1736 <= $signed(($unsigned($signed(reg1727)) ?
                  (wire1720 ^ (^~{reg87})) : (&(wire3 >> $unsigned(wire3)))));
              reg1737 <= ((&$unsigned((wire1[(2'h3):(1'h0)] << ((7'h48) + reg24)))) <<< reg1724[(4'he):(2'h3)]);
              reg1739 = reg67[(3'h6):(3'h5)];
            end
          if ((~&reg93[(2'h2):(1'h1)]))
            begin
              reg1740 <= (reg1728[(4'h8):(3'h6)] - (^~({(reg1735 | reg1737),
                      $unsigned(reg53)} ?
                  (reg1738[(1'h1):(1'h0)] ?
                      ((8'hbf) ?
                          reg29 : reg35) : $unsigned(reg14)) : (8'ha7))));
              reg1741 = reg35[(3'h6):(1'h0)];
              reg1742 = ($signed(reg1723[(3'h4):(2'h3)]) ?
                  (|$unsigned((~$signed(reg56)))) : ((({(8'hbc)} & (wire2 ?
                      (8'ha4) : forvar1722)) ^~ (reg1740 || wire0[(3'h6):(1'h1)])) >>> ($signed(reg87[(5'h10):(2'h3)]) | forvar1735)));
              reg1743 <= $unsigned((forvar1722 <<< reg1736));
            end
          else
            begin
              reg1740 <= (^$unsigned((reg29 ?
                  {$signed(forvar1735)} : ($unsigned(reg1737) != reg28[(4'ha):(1'h1)]))));
            end
          if ((reg1725 ? wire3 : reg17[(2'h2):(2'h2)]))
            begin
              reg1744 <= $unsigned((+$unsigned(reg43)));
              reg1745 = {$unsigned(({$unsigned((8'hb3))} < ((&reg15) | (forvar1735 | reg1738)))),
                  reg14[(2'h3):(1'h0)]};
              reg1746 = (^(!(+((~|reg1741) > reg1735))));
              reg1747 <= $signed(reg91);
              reg1748 = {(reg1735[(4'h9):(1'h0)] || (|$signed((7'h43)))),
                  $signed((reg1747 + $unsigned((reg1745 ? reg91 : reg47))))};
            end
          else
            begin
              reg1744 <= ($signed(reg34[(4'ha):(1'h1)]) >>> ((^$unsigned($unsigned(reg87))) ?
                  reg1745 : $signed((^~forvar1729))));
            end
          reg1749 = reg91;
        end
    end
  always
    @(posedge clk) begin
      if (reg1747)
        begin
          for (forvar1750 = (1'h0); (forvar1750 < (1'h1)); forvar1750 = (forvar1750 + (1'h1)))
            begin
              reg1751 = $signed($signed($unsigned(reg1732[(4'h8):(3'h6)])));
              reg1752 <= $signed(reg1747[(2'h2):(1'h0)]);
              reg1753 <= $signed(((~&(((8'hbd) ^~ reg54) + (forvar1750 * (8'had)))) <<< (reg1751[(2'h2):(2'h2)] ?
                  $unsigned($signed(reg17)) : reg1727)));
              reg1754 <= $unsigned((+(~^((-reg28) ?
                  {reg53} : ((7'h41) ? (7'h43) : reg43)))));
            end
          reg1755 = $unsigned(reg36[(2'h2):(1'h0)]);
          for (forvar1756 = (1'h0); (forvar1756 < (1'h0)); forvar1756 = (forvar1756 + (1'h1)))
            begin
              reg1757 <= (^(((reg13[(1'h0):(1'h0)] - {wire3}) ?
                      $unsigned(reg56[(2'h2):(1'h0)]) : (reg76[(4'h8):(3'h6)] ?
                          (8'hbb) : $unsigned(reg92))) ?
                  forvar1756 : (reg75 ?
                      ({reg47} != reg93[(2'h2):(1'h0)]) : reg1734[(5'h14):(4'he)])));
            end
        end
      else
        begin
          reg1750 <= forvar1756;
          reg1751 = reg14[(1'h0):(1'h0)];
        end
      for (forvar1758 = (1'h0); (forvar1758 < (3'h4)); forvar1758 = (forvar1758 + (1'h1)))
        begin
          for (forvar1759 = (1'h0); (forvar1759 < (1'h1)); forvar1759 = (forvar1759 + (1'h1)))
            begin
              reg1760 <= wire2[(5'h17):(4'hf)];
              reg1761 <= (~&({(reg23[(4'h9):(1'h0)] ?
                      (reg91 ? forvar1759 : reg1740) : (wire1 ?
                          reg1738 : reg1734))} + reg1751[(1'h0):(1'h0)]));
              reg1762 = reg36;
            end
          reg1763 <= ((reg1760[(2'h2):(2'h2)] & (+$signed((reg1732 ?
              reg1738 : reg58)))) || reg1734);
        end
      for (forvar1764 = (1'h0); (forvar1764 < (3'h4)); forvar1764 = (forvar1764 + (1'h1)))
        begin
          reg1765 = $unsigned(reg1732[(4'h9):(2'h2)]);
          reg1766 <= reg1757;
        end
      reg1767 <= $signed((reg17 ? reg58[(3'h6):(1'h1)] : wire2));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module95
#(parameter param1718 = {(({((8'ha1) >= (8'ha0))} ? {((8'hb9) ^ (8'hb4)), ((8'ha5) || (8'hac))} : (((8'h9e) ? (8'haa) : (7'h4a)) ? ((8'h9f) ? (7'h41) : (8'hbd)) : ((8'hbb) <= (8'hac)))) ? ((((8'hb4) ? (8'h9d) : (7'h4a)) ? (8'hb9) : ((7'h49) ^~ (8'ha4))) ? (((7'h42) ? (7'h46) : (8'hb7)) ^ ((8'ha6) ? (7'h46) : (8'ha6))) : (~|{(7'h40)})) : (+{{(8'hb8), (8'ha7)}, (^(7'h44))})), (((((8'hba) ~^ (8'hac)) ? {(8'hb4), (8'hbe)} : ((7'h47) ? (8'hab) : (8'haf))) * (((8'h9c) ? (8'ha9) : (7'h4a)) ? ((8'hb7) ? (8'hbf) : (8'ha4)) : (7'h41))) ~^ ((((8'hba) ? (7'h48) : (8'haa)) != ((8'hbf) ? (8'hb4) : (8'hab))) - (((8'hb2) ? (8'h9d) : (8'hbe)) ? ((8'ha0) & (8'ha5)) : ((8'had) ? (7'h44) : (7'h46)))))}, 
parameter param1719 = (+((((param1718 ~^ param1718) << (param1718 && param1718)) ? (^(-(7'h4a))) : ((~^param1718) || (+param1718))) ? param1718 : param1718)))
(y, clk, wire99, wire98, wire97, wire96);
  output wire [(32'ha3a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire99;
  input wire [(5'h13):(1'h0)] wire98;
  input wire signed [(4'h9):(1'h0)] wire97;
  input wire [(5'h10):(1'h0)] wire96;
  wire signed [(4'hc):(1'h0)] wire1717;
  wire signed [(4'hb):(1'h0)] wire1669;
  wire signed [(5'h13):(1'h0)] wire1619;
  wire signed [(5'h14):(1'h0)] wire802;
  wire [(4'hb):(1'h0)] wire800;
  wire signed [(5'h16):(1'h0)] wire102;
  wire [(5'h14):(1'h0)] wire101;
  wire signed [(5'h11):(1'h0)] wire100;
  wire [(5'h10):(1'h0)] wire1621;
  wire [(4'ha):(1'h0)] wire1664;
  wire signed [(5'h17):(1'h0)] wire1665;
  wire [(3'h4):(1'h0)] wire1666;
  reg [(4'hd):(1'h0)] reg1707 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1716 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1711 = (1'h0);
  reg [(4'hd):(1'h0)] reg1708 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1705 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1704 = (1'h0);
  reg [(5'h10):(1'h0)] reg1701 = (1'h0);
  reg [(5'h10):(1'h0)] reg1700 = (1'h0);
  reg [(4'ha):(1'h0)] reg1697 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1696 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1693 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1692 = (1'h0);
  reg [(4'hc):(1'h0)] reg1689 = (1'h0);
  reg [(4'hb):(1'h0)] reg1688 = (1'h0);
  reg [(4'hf):(1'h0)] reg1687 = (1'h0);
  reg [(2'h2):(1'h0)] reg1682 = (1'h0);
  reg [(4'hc):(1'h0)] reg1677 = (1'h0);
  reg [(5'h14):(1'h0)] reg1676 = (1'h0);
  reg [(5'h12):(1'h0)] reg1674 = (1'h0);
  reg [(4'hf):(1'h0)] reg1673 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1662 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1661 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1660 = (1'h0);
  reg [(5'h14):(1'h0)] reg1659 = (1'h0);
  reg [(4'hd):(1'h0)] reg1655 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1654 = (1'h0);
  reg [(3'h5):(1'h0)] reg1650 = (1'h0);
  reg [(3'h4):(1'h0)] reg1649 = (1'h0);
  reg [(5'h12):(1'h0)] reg1648 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1644 = (1'h0);
  reg [(5'h15):(1'h0)] reg1638 = (1'h0);
  reg [(4'h8):(1'h0)] reg1640 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1639 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1636 = (1'h0);
  reg [(5'h15):(1'h0)] reg1633 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1630 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1627 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1626 = (1'h0);
  reg [(5'h11):(1'h0)] reg1624 = (1'h0);
  reg [(4'he):(1'h0)] reg1623 = (1'h0);
  reg [(5'h12):(1'h0)] reg804 = (1'h0);
  reg [(4'ha):(1'h0)] reg805 = (1'h0);
  reg [(5'h10):(1'h0)] reg806 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg807 = (1'h0);
  reg [(3'h6):(1'h0)] reg810 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg811 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg812 = (1'h0);
  reg [(4'h8):(1'h0)] reg813 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg817 = (1'h0);
  reg [(4'hf):(1'h0)] reg819 = (1'h0);
  reg [(3'h4):(1'h0)] reg821 = (1'h0);
  reg [(5'h18):(1'h0)] reg826 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg829 = (1'h0);
  reg [(2'h2):(1'h0)] reg830 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg832 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg840 = (1'h0);
  reg [(4'h8):(1'h0)] reg843 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg846 = (1'h0);
  reg [(3'h4):(1'h0)] reg847 = (1'h0);
  reg [(5'h14):(1'h0)] reg849 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg851 = (1'h0);
  reg [(3'h7):(1'h0)] reg852 = (1'h0);
  reg [(5'h14):(1'h0)] reg853 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg854 = (1'h0);
  reg [(5'h16):(1'h0)] reg855 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg858 = (1'h0);
  reg [(5'h10):(1'h0)] reg859 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg861 = (1'h0);
  reg [(4'h8):(1'h0)] reg863 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg865 = (1'h0);
  reg [(2'h3):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg869 = (1'h0);
  reg [(5'h11):(1'h0)] reg874 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg875 = (1'h0);
  reg [(5'h14):(1'h0)] reg876 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg877 = (1'h0);
  reg [(5'h18):(1'h0)] reg878 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg883 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg885 = (1'h0);
  reg [(4'he):(1'h0)] reg886 = (1'h0);
  reg [(5'h12):(1'h0)] reg888 = (1'h0);
  reg [(5'h12):(1'h0)] reg889 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg890 = (1'h0);
  reg [(2'h2):(1'h0)] reg891 = (1'h0);
  reg [(2'h3):(1'h0)] reg892 = (1'h0);
  reg [(4'hd):(1'h0)] reg893 = (1'h0);
  reg [(4'hb):(1'h0)] reg887 = (1'h0);
  reg [(4'hd):(1'h0)] reg1712 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1709 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1715 = (1'h0);
  reg [(3'h5):(1'h0)] reg1714 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1713 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1712 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1710 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1709 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1707 = (1'h0);
  reg [(5'h11):(1'h0)] reg1706 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1703 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1702 = (1'h0);
  reg [(4'hf):(1'h0)] reg1699 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1692 = (1'h0);
  reg [(5'h17):(1'h0)] reg1691 = (1'h0);
  reg [(3'h5):(1'h0)] reg1698 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1695 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1694 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1691 = (1'h0);
  reg [(5'h11):(1'h0)] reg1690 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1686 = (1'h0);
  reg [(5'h14):(1'h0)] reg1685 = (1'h0);
  reg [(4'hc):(1'h0)] reg1684 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1683 = (1'h0);
  reg [(5'h11):(1'h0)] reg1681 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1680 = (1'h0);
  reg [(2'h2):(1'h0)] reg1679 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1678 = (1'h0);
  reg [(4'h8):(1'h0)] reg1675 = (1'h0);
  reg [(5'h11):(1'h0)] reg1672 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1671 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1670 = (1'h0);
  reg [(2'h3):(1'h0)] reg1668 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1663 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1658 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1657 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1656 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1653 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1652 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1651 = (1'h0);
  reg [(4'ha):(1'h0)] reg1647 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1647 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1646 = (1'h0);
  reg [(4'hb):(1'h0)] reg1645 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1637 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1643 = (1'h0);
  reg [(3'h5):(1'h0)] reg1642 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1641 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1638 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1637 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1622 = (1'h0);
  reg [(5'h14):(1'h0)] reg1635 = (1'h0);
  reg [(3'h7):(1'h0)] reg1634 = (1'h0);
  reg [(5'h14):(1'h0)] reg1632 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1631 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1629 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1628 = (1'h0);
  reg [(5'h17):(1'h0)] reg1625 = (1'h0);
  reg [(5'h15):(1'h0)] reg1622 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg895 = (1'h0);
  reg [(3'h4):(1'h0)] reg894 = (1'h0);
  reg [(5'h17):(1'h0)] forvar887 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg884 = (1'h0);
  reg [(4'hb):(1'h0)] forvar882 = (1'h0);
  reg [(3'h6):(1'h0)] reg881 = (1'h0);
  reg [(4'h9):(1'h0)] reg880 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg879 = (1'h0);
  reg [(4'hb):(1'h0)] reg873 = (1'h0);
  reg [(3'h5):(1'h0)] forvar872 = (1'h0);
  reg [(4'hf):(1'h0)] reg871 = (1'h0);
  reg [(2'h2):(1'h0)] reg870 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg867 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg866 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg862 = (1'h0);
  reg [(5'h15):(1'h0)] forvar860 = (1'h0);
  reg [(3'h4):(1'h0)] forvar847 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg857 = (1'h0);
  reg [(5'h11):(1'h0)] reg856 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg850 = (1'h0);
  reg [(3'h6):(1'h0)] reg848 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg845 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg844 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg842 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg841 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg839 = (1'h0);
  reg [(3'h6):(1'h0)] reg838 = (1'h0);
  reg [(4'he):(1'h0)] forvar837 = (1'h0);
  reg [(2'h3):(1'h0)] reg836 = (1'h0);
  reg [(3'h7):(1'h0)] reg835 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar834 = (1'h0);
  reg [(5'h12):(1'h0)] reg833 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg831 = (1'h0);
  reg [(4'he):(1'h0)] forvar825 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg828 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg827 = (1'h0);
  reg [(5'h11):(1'h0)] reg825 = (1'h0);
  reg [(2'h2):(1'h0)] reg824 = (1'h0);
  reg [(5'h14):(1'h0)] reg823 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar822 = (1'h0);
  reg [(3'h6):(1'h0)] reg820 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg818 = (1'h0);
  reg [(4'hd):(1'h0)] reg816 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar815 = (1'h0);
  reg [(5'h11):(1'h0)] forvar814 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg809 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg808 = (1'h0);
  reg [(3'h7):(1'h0)] forvar803 = (1'h0);
  assign y = {wire1717,
                 wire1669,
                 wire1619,
                 wire802,
                 wire800,
                 wire102,
                 wire101,
                 wire100,
                 wire1621,
                 wire1664,
                 wire1665,
                 wire1666,
                 reg1707,
                 reg1716,
                 reg1711,
                 reg1708,
                 reg1705,
                 reg1704,
                 reg1701,
                 reg1700,
                 reg1697,
                 reg1696,
                 reg1693,
                 reg1692,
                 reg1689,
                 reg1688,
                 reg1687,
                 reg1682,
                 reg1677,
                 reg1676,
                 reg1674,
                 reg1673,
                 reg1662,
                 reg1661,
                 reg1660,
                 reg1659,
                 reg1655,
                 reg1654,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1644,
                 reg1638,
                 reg1640,
                 reg1639,
                 reg1636,
                 reg1633,
                 reg1630,
                 reg1627,
                 reg1626,
                 reg1624,
                 reg1623,
                 reg804,
                 reg805,
                 reg806,
                 reg807,
                 reg810,
                 reg811,
                 reg812,
                 reg813,
                 reg817,
                 reg819,
                 reg821,
                 reg826,
                 reg829,
                 reg830,
                 reg832,
                 reg840,
                 reg843,
                 reg846,
                 reg847,
                 reg849,
                 reg851,
                 reg852,
                 reg853,
                 reg854,
                 reg855,
                 reg858,
                 reg859,
                 reg861,
                 reg863,
                 reg865,
                 reg868,
                 reg869,
                 reg874,
                 reg875,
                 reg876,
                 reg877,
                 reg878,
                 reg883,
                 reg885,
                 reg886,
                 reg888,
                 reg889,
                 reg890,
                 reg891,
                 reg892,
                 reg893,
                 reg887,
                 reg1712,
                 reg1709,
                 reg1715,
                 reg1714,
                 reg1713,
                 forvar1712,
                 reg1710,
                 forvar1709,
                 forvar1707,
                 reg1706,
                 forvar1703,
                 reg1702,
                 reg1699,
                 forvar1692,
                 reg1691,
                 reg1698,
                 reg1695,
                 reg1694,
                 forvar1691,
                 reg1690,
                 reg1686,
                 reg1685,
                 reg1684,
                 reg1683,
                 reg1681,
                 reg1680,
                 reg1679,
                 forvar1678,
                 reg1675,
                 reg1672,
                 forvar1671,
                 reg1670,
                 reg1668,
                 reg1663,
                 reg1658,
                 reg1657,
                 reg1656,
                 reg1653,
                 forvar1652,
                 reg1651,
                 reg1647,
                 forvar1647,
                 reg1646,
                 reg1645,
                 forvar1637,
                 reg1643,
                 reg1642,
                 reg1641,
                 forvar1638,
                 reg1637,
                 forvar1622,
                 reg1635,
                 reg1634,
                 reg1632,
                 forvar1631,
                 reg1629,
                 reg1628,
                 reg1625,
                 reg1622,
                 reg895,
                 reg894,
                 forvar887,
                 reg884,
                 forvar882,
                 reg881,
                 reg880,
                 reg879,
                 reg873,
                 forvar872,
                 reg871,
                 reg870,
                 reg867,
                 reg866,
                 reg864,
                 reg862,
                 forvar860,
                 forvar847,
                 reg857,
                 reg856,
                 reg850,
                 reg848,
                 reg845,
                 reg844,
                 reg842,
                 reg841,
                 reg839,
                 reg838,
                 forvar837,
                 reg836,
                 reg835,
                 forvar834,
                 reg833,
                 reg831,
                 forvar825,
                 reg828,
                 reg827,
                 reg825,
                 reg824,
                 reg823,
                 forvar822,
                 reg820,
                 reg818,
                 reg816,
                 forvar815,
                 forvar814,
                 reg809,
                 reg808,
                 forvar803,
                 (1'h0)};
  assign wire100 = (($signed($signed((wire96 ?
                       wire99 : wire98))) < {wire97[(3'h7):(3'h7)]}) || wire98[(4'hb):(3'h4)]);
  assign wire101 = $unsigned((!$unsigned(wire99)));
  assign wire102 = $unsigned((~^wire96[(3'h7):(3'h6)]));
  module103 #() modinst801 (.wire104(wire98), .wire106(wire101), .clk(clk), .wire107(wire96), .wire105(wire99), .y(wire800));
  assign wire802 = ($unsigned(($unsigned(wire97) ?
                       wire96[(2'h3):(2'h3)] : $signed((wire96 ^~ wire800)))) | $signed(($signed((^~wire98)) ?
                       ({wire800, wire97} ?
                           $unsigned((8'hb4)) : $signed(wire96)) : (^$signed(wire98)))));
  always
    @(posedge clk) begin
      for (forvar803 = (1'h0); (forvar803 < (2'h3)); forvar803 = (forvar803 + (1'h1)))
        begin
          reg804 <= ($unsigned($unsigned((^~{wire100}))) >> ({$signed($unsigned(wire96))} ?
              wire800 : wire96[(1'h0):(1'h0)]));
          if ({wire802[(5'h14):(4'hf)],
              $unsigned({(!(wire102 ? wire96 : wire96)), wire802})})
            begin
              reg805 <= ((~wire98[(4'hd):(4'ha)]) ?
                  $unsigned($unsigned(wire96)) : $unsigned({(^~(8'hb8))}));
              reg806 <= (~|(($unsigned($signed(forvar803)) < (+wire97[(1'h1):(1'h1)])) ~^ {(wire98 ~^ $unsigned(wire99))}));
              reg807 <= reg804[(5'h12):(3'h7)];
              reg808 = (~^{$signed((wire102 ? (wire101 ~^ (8'ha6)) : (8'ha1))),
                  reg806});
              reg809 = reg807;
            end
          else
            begin
              reg805 <= wire97;
              reg806 <= $unsigned({reg805[(4'h9):(2'h2)]});
              reg807 <= wire800[(4'h8):(1'h1)];
              reg810 <= (+(+(&$signed($signed(wire100)))));
              reg811 <= reg808;
            end
        end
      reg812 <= reg808[(4'ha):(2'h2)];
      reg813 <= $unsigned($signed(reg810[(3'h5):(1'h0)]));
      for (forvar814 = (1'h0); (forvar814 < (3'h4)); forvar814 = (forvar814 + (1'h1)))
        begin
          for (forvar815 = (1'h0); (forvar815 < (2'h3)); forvar815 = (forvar815 + (1'h1)))
            begin
              reg816 = $unsigned($signed($signed((reg808 ~^ (reg804 ^~ wire102)))));
            end
          if ((wire101[(4'hd):(3'h7)] ~^ (^((~&(wire800 ?
              reg809 : (8'hbc))) > wire800[(1'h0):(1'h0)]))))
            begin
              reg817 <= ((((reg804[(3'h7):(1'h0)] ?
                      $signed(wire100) : (&reg806)) != {wire96[(4'hb):(2'h2)]}) ?
                  (7'h41) : {(wire99[(3'h6):(3'h6)] && $signed(forvar803)),
                      wire96[(3'h6):(2'h3)]}) >= $signed({wire97}));
              reg818 = reg811;
              reg819 <= reg804;
              reg820 = $unsigned((!forvar803));
            end
          else
            begin
              reg817 <= ((8'had) ?
                  {((^$unsigned(reg819)) ? (^(reg807 > wire99)) : {wire98}),
                      $signed(reg818)} : wire99);
              reg819 <= reg807[(5'h10):(5'h10)];
              reg821 <= reg811;
            end
          for (forvar822 = (1'h0); (forvar822 < (2'h2)); forvar822 = (forvar822 + (1'h1)))
            begin
              reg823 = (reg812 ?
                  $signed(reg821[(2'h3):(2'h3)]) : {(wire100[(1'h1):(1'h0)] || reg805[(1'h1):(1'h0)])});
            end
          reg824 = (($signed((~((8'hb6) ? reg808 : reg823))) ?
                  (forvar814 ?
                      $unsigned(((8'haf) ?
                          wire99 : reg811)) : reg811) : (reg808[(4'hc):(3'h4)] - ((^~wire101) ?
                      reg819[(4'ha):(1'h1)] : $unsigned(wire802)))) ?
              $unsigned($signed($signed($unsigned(reg811)))) : (((wire96[(4'ha):(3'h4)] ^ $unsigned(reg804)) ?
                  (^~(&reg806)) : $signed({reg813, wire102})) < wire800));
        end
    end
  always
    @(posedge clk) begin
      if ((((^~$unsigned((reg810 - reg806))) && $signed(($unsigned(reg817) & reg810))) ?
          wire102 : $unsigned($signed(((reg821 ? (8'hbf) : wire102) ?
              $signed(reg810) : ((7'h45) ? wire800 : (8'hbe)))))))
        begin
          reg825 = $signed((!$signed((8'hab))));
          reg826 <= ((reg811[(2'h3):(1'h0)] ?
              $signed(reg825) : reg807[(3'h6):(3'h4)]) ~^ $unsigned({reg817[(1'h1):(1'h0)]}));
          reg827 = (8'hb9);
          reg828 = {{$unsigned({(reg819 ? reg825 : wire96)}),
                  $signed({$unsigned(reg807), (reg827 ? wire800 : reg819)})},
              ((+(8'hbb)) >> (reg804 ?
                  reg813[(1'h0):(1'h0)] : wire97[(4'h9):(1'h1)]))};
        end
      else
        begin
          for (forvar825 = (1'h0); (forvar825 < (3'h4)); forvar825 = (forvar825 + (1'h1)))
            begin
              reg827 = wire97[(1'h0):(1'h0)];
              reg829 <= {$signed({($unsigned(reg817) ?
                          $unsigned(forvar825) : $unsigned((7'h46)))}),
                  ($signed(((reg811 ? wire102 : reg827) ?
                      (|wire98) : $unsigned(wire97))) < reg828[(1'h0):(1'h0)])};
              reg830 <= wire98;
              reg831 = reg825;
              reg832 <= reg826;
            end
        end
      reg833 = (^($signed(({reg810} > (wire100 ? (8'ha2) : wire101))) ?
          (reg827[(4'h9):(3'h6)] >= {reg804[(2'h2):(2'h2)],
              reg812[(5'h11):(2'h3)]}) : (reg810 * (reg828 ?
              reg813 : (reg827 || (8'hb9))))));
      for (forvar834 = (1'h0); (forvar834 < (1'h1)); forvar834 = (forvar834 + (1'h1)))
        begin
          reg835 = {wire98};
          reg836 = (!$signed((+reg811[(1'h0):(1'h0)])));
          for (forvar837 = (1'h0); (forvar837 < (1'h1)); forvar837 = (forvar837 + (1'h1)))
            begin
              reg838 = {($unsigned((!$unsigned(forvar825))) ?
                      {(&(7'h48)),
                          wire102[(2'h2):(1'h0)]} : $unsigned($signed((^reg819)))),
                  {(reg830[(1'h1):(1'h0)] ? forvar837 : wire100[(4'h9):(3'h6)]),
                      reg831[(2'h3):(2'h2)]}};
              reg839 = (reg838 <= (-reg828[(4'ha):(3'h5)]));
              reg840 <= (!reg806[(4'ha):(4'ha)]);
              reg841 = (|(reg819 ?
                  ((-wire97[(4'h9):(1'h1)]) ?
                      wire99[(4'h9):(4'h9)] : ((wire99 | reg825) ?
                          reg807[(3'h5):(3'h5)] : $signed(forvar834))) : $signed($signed($signed(reg831)))));
              reg842 = (!reg826);
            end
          reg843 <= {$unsigned(reg806[(3'h5):(2'h2)])};
        end
    end
  always
    @(posedge clk) begin
      reg844 = (~^($unsigned($unsigned(reg807[(4'h8):(3'h7)])) ?
          reg840 : ((~(&(8'ha3))) ? (8'h9d) : {(wire96 != wire98)})));
    end
  always
    @(posedge clk) begin
      if ($unsigned($signed(reg821)))
        begin
          reg845 = (reg805 ?
              {$signed({reg805}),
                  (-reg830)} : (((-(reg832 << reg830)) ^~ reg826) ^~ $unsigned(($unsigned(wire102) ?
                  (^~reg812) : $signed(wire800)))));
          if ((($unsigned($unsigned({wire101, wire101})) * {((wire102 ?
                      reg821 : reg811) | reg813),
                  wire100[(2'h2):(2'h2)]}) ?
              reg807 : ((~|$signed($unsigned(wire100))) ?
                  (|$unsigned({wire100, wire100})) : ((|$unsigned(reg811)) ?
                      reg810 : {$signed(reg817)}))))
            begin
              reg846 <= $signed((~((^$unsigned(reg832)) != (^~{wire98}))));
              reg847 <= {{({$signed(reg819)} & (reg832 <<< (&(7'h45)))),
                      $signed(($signed(reg805) ~^ reg805))}};
              reg848 = reg826;
              reg849 <= reg829[(1'h1):(1'h0)];
            end
          else
            begin
              reg848 = wire100;
              reg850 = $signed((8'hbe));
              reg851 <= reg846;
              reg852 <= $unsigned({(^~$unsigned((reg851 ? wire802 : reg846))),
                  wire98});
              reg853 <= (&$signed((reg830 == $unsigned($signed(reg852)))));
            end
          reg854 <= $signed(((wire102[(1'h1):(1'h1)] <<< ((reg807 || wire97) ?
              reg821[(2'h2):(1'h0)] : (+reg805))) + reg811));
          if ((|reg840[(3'h4):(3'h4)]))
            begin
              reg855 <= (~&wire102[(4'h9):(2'h3)]);
              reg856 = reg811[(2'h3):(2'h2)];
              reg857 = $signed(((8'ha6) ? reg819[(4'hc):(2'h2)] : reg830));
              reg858 <= ((~&$signed($unsigned(reg826[(3'h6):(1'h1)]))) >> $unsigned($unsigned({reg840[(3'h5):(1'h0)]})));
              reg859 <= (~|reg807[(3'h4):(1'h0)]);
            end
          else
            begin
              reg855 <= $signed(((^~wire102) ?
                  {reg840,
                      $signed((reg843 ?
                          reg858 : reg845))} : $signed((|reg830))));
              reg856 = (((~|reg851) && reg813) != (reg854 <<< (((|reg806) ?
                  ((8'hb6) <<< reg812) : $signed(reg821)) >= $signed(reg851))));
              reg857 = (~^$unsigned($unsigned((reg840 ?
                  (~^reg840) : $unsigned((8'ha7))))));
              reg858 <= $unsigned((~((^~$unsigned(wire96)) | $signed((reg819 >= (8'hae))))));
            end
        end
      else
        begin
          reg845 = $signed((^~$unsigned((~$unsigned(wire800)))));
          reg846 <= reg854;
          for (forvar847 = (1'h0); (forvar847 < (3'h4)); forvar847 = (forvar847 + (1'h1)))
            begin
              reg848 = (~|(wire101 + ($unsigned((wire100 ? reg829 : wire97)) ?
                  $signed($unsigned(reg845)) : reg810[(2'h2):(1'h1)])));
              reg850 = reg804[(2'h3):(2'h2)];
              reg856 = reg840[(4'hf):(4'hc)];
              reg857 = {$unsigned((!(~&wire99[(2'h2):(1'h0)])))};
            end
        end
      for (forvar860 = (1'h0); (forvar860 < (1'h1)); forvar860 = (forvar860 + (1'h1)))
        begin
          if ((!$unsigned(((~^((8'h9f) ? (7'h49) : reg849)) ?
              $signed((reg804 ? reg821 : reg829)) : {(reg817 | reg806),
                  (+reg840)}))))
            begin
              reg861 <= $unsigned($signed(($unsigned($signed(reg847)) & (reg807 ?
                  (&forvar847) : (reg830 ? reg846 : reg830)))));
              reg862 = wire102[(5'h14):(4'hc)];
              reg863 <= reg855;
              reg864 = ($unsigned((reg861[(2'h2):(2'h2)] == $signed($unsigned(reg843)))) ?
                  $signed(reg847[(3'h4):(2'h2)]) : wire101);
              reg865 <= reg853[(1'h0):(1'h0)];
            end
          else
            begin
              reg862 = {{reg857, ((&wire102) <= {reg821[(2'h3):(2'h3)]})},
                  ((reg857 ?
                          reg811[(1'h0):(1'h0)] : (reg855[(2'h2):(1'h1)] + (&reg829))) ?
                      $signed(((reg859 ^ reg812) ^~ $signed(wire98))) : reg865[(1'h1):(1'h0)])};
              reg863 <= reg853[(4'h8):(3'h5)];
              reg865 <= $signed(wire96);
            end
          if ((reg849[(2'h2):(1'h0)] ?
              ((reg819 ?
                  reg805[(2'h3):(1'h0)] : ((reg830 <<< reg817) ?
                      $unsigned(reg829) : $signed(reg832))) || reg854) : (^$unsigned($unsigned((reg811 ?
                  reg865 : reg855))))))
            begin
              reg866 = $signed($unsigned({reg804}));
              reg867 = reg806;
            end
          else
            begin
              reg866 = $signed((&{$unsigned($signed((7'h40))),
                  (reg821[(2'h3):(1'h0)] >>> (^~(8'hb7)))}));
              reg868 <= reg805;
              reg869 <= wire102[(5'h11):(2'h2)];
              reg870 = reg859[(4'h9):(3'h6)];
              reg871 = $unsigned($signed(({(&reg817)} < ($signed(reg850) <= (^~reg869)))));
            end
          for (forvar872 = (1'h0); (forvar872 < (1'h0)); forvar872 = (forvar872 + (1'h1)))
            begin
              reg873 = $unsigned($signed((^~$unsigned($signed(wire101)))));
              reg874 <= $signed((+({reg856[(2'h2):(1'h1)],
                  $signed(forvar847)} >>> (+$signed(wire802)))));
              reg875 <= $unsigned({{$signed(reg846[(2'h2):(1'h0)]),
                      {reg855[(3'h7):(1'h0)], reg861}},
                  ($unsigned((reg861 & reg845)) + reg854)});
              reg876 <= reg851[(4'he):(2'h2)];
              reg877 <= $signed((wire800 + ((~^reg847[(2'h3):(1'h1)]) == reg852)));
            end
          reg878 <= ($unsigned(({(reg840 ? reg867 : (8'h9f)), $signed(reg850)} ?
                  $signed((~|wire800)) : $unsigned($signed((8'hae))))) ?
              (|(8'ha0)) : ((wire102 ?
                  wire97[(4'h9):(3'h6)] : ($signed(reg819) ?
                      reg821[(1'h1):(1'h1)] : {reg846})) - reg832));
        end
      reg879 = $signed((reg830 < $unsigned((reg874 ?
          (reg819 ? (8'had) : reg826) : (reg873 <<< reg821)))));
      if ((-reg876))
        begin
          reg880 = reg877;
        end
      else
        begin
          reg880 = reg879;
          reg881 = (~(reg871[(4'hb):(2'h3)] ?
              reg807 : $unsigned(($signed((8'hae)) ?
                  (!reg852) : ((8'ha0) + reg804)))));
          for (forvar882 = (1'h0); (forvar882 < (3'h4)); forvar882 = (forvar882 + (1'h1)))
            begin
              reg883 <= ($unsigned((!$signed((forvar860 ?
                  reg866 : reg810)))) * reg868[(1'h1):(1'h0)]);
              reg884 = (~reg852[(1'h1):(1'h1)]);
            end
          reg885 <= {((reg857[(3'h5):(3'h4)] || reg868) * reg880),
              (~|$unsigned((wire100[(3'h4):(1'h0)] ?
                  $signed(wire802) : {reg810, reg870})))};
        end
      if ((|$signed(reg856)))
        begin
          reg886 <= reg881;
          for (forvar887 = (1'h0); (forvar887 < (1'h0)); forvar887 = (forvar887 + (1'h1)))
            begin
              reg888 <= $unsigned(reg807[(3'h7):(1'h0)]);
              reg889 <= reg879;
            end
          if ($signed(reg876))
            begin
              reg890 <= $signed((~&$unsigned(($signed(wire800) ?
                  (~^reg830) : $unsigned((8'ha0))))));
              reg891 <= wire800[(3'h7):(3'h7)];
              reg892 <= (-$signed((wire99[(1'h0):(1'h0)] * $signed($signed(reg829)))));
              reg893 <= reg806;
            end
          else
            begin
              reg894 = ((reg813[(3'h4):(3'h4)] ?
                  (~reg819[(4'ha):(3'h7)]) : ($signed((~reg866)) - ({reg846} ?
                      $unsigned(reg819) : wire802))) == {$signed(($signed(reg862) ?
                      reg829[(2'h2):(1'h1)] : $unsigned(reg871)))});
              reg895 = ($unsigned(($unsigned({(7'h40)}) ?
                  ($signed((8'hbe)) ?
                      $signed(reg889) : $signed(reg864)) : reg806)) & ((reg810[(1'h1):(1'h0)] ?
                  (~&reg874[(4'h9):(2'h2)]) : reg812) * reg873));
            end
        end
      else
        begin
          reg886 <= ($signed(wire97) ?
              (((^reg877) && reg806[(4'hb):(2'h3)]) <= reg804[(5'h11):(3'h7)]) : $signed((reg810 ?
                  (((8'hac) ^~ reg894) ?
                      (~(8'haf)) : reg843) : ((^~wire102) <= (&(8'hb2))))));
          reg887 <= (~|(reg806[(3'h4):(3'h4)] ?
              reg804 : $signed((~|((8'hbe) | reg853)))));
          reg888 <= $unsigned((((8'ha7) ? reg854[(4'h8):(1'h0)] : reg811) ?
              (reg879 ?
                  reg868[(2'h2):(1'h1)] : ($signed(reg871) ~^ (reg857 ?
                      (8'h9e) : (7'h41)))) : (($signed(reg874) ?
                      {(8'h9d)} : reg850[(1'h0):(1'h0)]) ?
                  (reg850 ?
                      $signed(reg881) : $signed(wire101)) : $unsigned((-forvar872)))));
        end
    end
  module896 #() modinst1620 (.wire900(wire96), .clk(clk), .wire898(reg887), .wire897(reg829), .y(wire1619), .wire899(reg812));
  assign wire1621 = (&($signed(reg805) ?
                        ({$unsigned(reg849)} ?
                            $signed((8'haa)) : reg883) : $signed(reg863)));
  always
    @(posedge clk) begin
      if (((^~($unsigned(reg830) != ({reg888} <= reg886))) - ((^~reg853) << ($signed($unsigned(reg819)) >= (reg854 ?
          (wire99 * (8'hb5)) : $unsigned(reg876))))))
        begin
          if ((reg883 + reg874))
            begin
              reg1622 = wire102[(5'h12):(1'h1)];
              reg1623 <= (^reg886);
              reg1624 <= (-{(((reg1623 < (7'h42)) ?
                      (reg811 <= reg861) : (reg874 >= reg819)) ^~ $unsigned(reg855[(4'h8):(3'h7)])),
                  reg885});
              reg1625 = {wire97, $unsigned($unsigned(reg868))};
            end
          else
            begin
              reg1623 <= ($unsigned((reg832 - ($unsigned(wire96) ?
                      reg846[(1'h1):(1'h1)] : $signed((8'hb3))))) ?
                  $unsigned($signed(reg829[(5'h11):(3'h7)])) : ($unsigned(({reg807} ?
                      (reg1622 | reg875) : $signed(reg885))) != $unsigned($unsigned($unsigned(reg854)))));
              reg1625 = ((~reg875) ?
                  reg891 : (((^reg886) >= $signed((~&reg855))) ?
                      $signed(((reg819 >= reg832) || $signed(reg1623))) : $unsigned(reg805)));
              reg1626 <= $signed(reg819);
            end
          if ($signed((reg1623[(2'h3):(2'h2)] + reg849[(5'h12):(3'h7)])))
            begin
              reg1627 <= ((reg885 < ((^~(reg847 ?
                      wire102 : reg859)) <<< $unsigned((reg1626 + reg1622)))) ?
                  (&$unsigned((reg1626[(3'h5):(2'h2)] <<< (reg878 == reg877)))) : (~&($unsigned(reg888[(4'h9):(3'h4)]) ?
                      ($signed(reg851) <= $signed(reg810)) : reg806)));
              reg1628 = wire99;
              reg1629 = ((+$signed((-(reg851 >> (8'hab))))) ?
                  {{(|$unsigned(wire800))}} : $unsigned((~&$signed(reg1624[(5'h11):(3'h7)]))));
              reg1630 <= (($signed(((reg1629 <= wire97) ?
                          {reg829, (8'hb4)} : (wire96 ? (8'hbd) : reg891))) ?
                      {((^~reg810) <<< {reg1625})} : reg810[(2'h2):(1'h0)]) ?
                  reg1625[(1'h0):(1'h0)] : (reg840 ? reg1623 : reg806));
            end
          else
            begin
              reg1628 = ($signed(((^~$unsigned(reg889)) ?
                  reg821[(1'h0):(1'h0)] : reg877[(4'ha):(3'h7)])) ^~ ($signed((reg875 ?
                      (reg874 == reg883) : ((8'hbd) ? reg830 : reg859))) ?
                  (~&$signed($unsigned(reg851))) : $signed($unsigned(wire800))));
              reg1630 <= (8'h9e);
            end
          for (forvar1631 = (1'h0); (forvar1631 < (2'h3)); forvar1631 = (forvar1631 + (1'h1)))
            begin
              reg1632 = ((^$signed((!(reg863 ?
                  reg1623 : reg886)))) - (^(&$signed($unsigned(reg853)))));
              reg1633 <= (|(+(8'ha8)));
              reg1634 = $signed(((~&reg859[(3'h5):(1'h1)]) + reg892));
              reg1635 = (reg851 ^~ $unsigned((~^$signed({reg830}))));
              reg1636 <= (($unsigned((reg821 ~^ reg829[(4'he):(4'hd)])) & reg1635[(5'h13):(2'h2)]) * ($unsigned(((reg855 > reg826) >> (wire101 > reg805))) != {(reg859 >> reg829),
                  reg829[(5'h10):(3'h6)]}));
            end
        end
      else
        begin
          for (forvar1622 = (1'h0); (forvar1622 < (3'h4)); forvar1622 = (forvar1622 + (1'h1)))
            begin
              reg1623 <= ((+{(^$unsigned(reg876)), wire100}) ?
                  reg877 : $unsigned(forvar1631[(4'h9):(4'h8)]));
              reg1624 <= wire102;
            end
        end
      if (reg1625)
        begin
          reg1637 = reg893;
          for (forvar1638 = (1'h0); (forvar1638 < (2'h2)); forvar1638 = (forvar1638 + (1'h1)))
            begin
              reg1639 <= {reg886[(4'hb):(4'hb)], wire802[(3'h6):(2'h2)]};
              reg1640 <= (($signed((|$unsigned(wire800))) ?
                      (|$signed(((7'h40) ?
                          (7'h47) : (7'h41)))) : reg843[(3'h4):(1'h0)]) ?
                  reg813 : ($unsigned((8'ha8)) | (^~((reg1633 & reg888) && reg810))));
            end
          reg1641 = (^$signed($unsigned($signed($signed(reg826)))));
          reg1642 = $signed($unsigned(({(7'h45)} ?
              (-(wire97 ? reg812 : (8'ha0))) : ((wire800 || wire1619) ?
                  (^~reg810) : (~reg813)))));
          reg1643 = $signed(reg887[(4'ha):(4'h9)]);
        end
      else
        begin
          for (forvar1637 = (1'h0); (forvar1637 < (1'h1)); forvar1637 = (forvar1637 + (1'h1)))
            begin
              reg1638 <= ((wire100[(4'hc):(4'hb)] ?
                  forvar1631[(5'h10):(1'h0)] : {($unsigned(reg878) ~^ ((8'hbe) || reg830)),
                      reg859}) <= ((8'hae) ?
                  ($unsigned($signed(reg817)) ?
                      $unsigned($unsigned(reg840)) : ($unsigned(reg868) ?
                          $signed(reg1640) : (~|wire99))) : {{$unsigned(reg829)},
                      ((8'ha9) >> wire1621)}));
              reg1639 <= {(((8'hb8) ?
                          {(reg851 ? reg865 : reg1626),
                              $signed(reg846)} : ((~|reg811) + (+reg1636))) ?
                      $unsigned((~((8'ha4) ?
                          reg885 : wire1621))) : (reg1643 >> reg853[(3'h6):(1'h1)])),
                  (+$unsigned(reg811))};
              reg1641 = reg812[(3'h7):(3'h6)];
              reg1644 <= $signed(($signed(wire98[(1'h0):(1'h0)]) ?
                  reg807[(5'h13):(5'h12)] : reg1633[(3'h5):(3'h4)]));
              reg1645 = ({reg1630} ?
                  $unsigned(reg865[(1'h1):(1'h1)]) : ($signed(((!reg806) ?
                      reg893 : {reg810,
                          reg1639})) || $unsigned(($unsigned((8'haa)) ?
                      (forvar1637 ? reg877 : reg1632) : {wire102, (8'hb4)}))));
            end
          reg1646 = (~|$signed((((wire97 ^~ reg1645) ?
              $signed(reg812) : (|reg847)) + {$unsigned(reg840),
              ((7'h41) ? reg1633 : reg843)})));
        end
      if ($unsigned((^(~reg1643))))
        begin
          for (forvar1647 = (1'h0); (forvar1647 < (2'h2)); forvar1647 = (forvar1647 + (1'h1)))
            begin
              reg1648 <= reg807[(4'hc):(3'h4)];
              reg1649 <= ((((|(reg852 ? reg819 : wire98)) ?
                          (8'ha4) : ((~|reg810) != {reg840})) ?
                      ({$unsigned(reg806), reg1625[(5'h13):(5'h13)]} ?
                          wire800 : reg1645) : reg855) ?
                  reg830[(2'h2):(1'h0)] : $signed(reg892));
              reg1650 <= $signed(reg886[(2'h3):(1'h0)]);
            end
        end
      else
        begin
          reg1647 = $unsigned(($unsigned($unsigned((reg1629 >= reg830))) ?
              $signed(reg1632) : (^((^~reg1635) ?
                  $signed(reg887) : $unsigned(reg812)))));
          reg1648 <= (~&reg883);
          reg1651 = (8'hb9);
          for (forvar1652 = (1'h0); (forvar1652 < (3'h4)); forvar1652 = (forvar1652 + (1'h1)))
            begin
              reg1653 = $unsigned(reg853);
              reg1654 <= {(^(^~$signed(reg893[(1'h1):(1'h1)])))};
              reg1655 <= $unsigned(((((~|reg1647) >> {(8'had)}) + reg855[(4'hd):(4'hc)]) ?
                  wire96 : $unsigned(($unsigned(wire98) ?
                      reg826 : $signed(wire101)))));
            end
          if (wire99[(4'h8):(3'h7)])
            begin
              reg1656 = (&((reg1627 & $signed((-reg889))) ?
                  {$unsigned(reg854[(3'h6):(2'h3)]),
                      (reg843[(3'h6):(3'h6)] ?
                          reg893[(3'h6):(2'h3)] : reg832[(3'h5):(2'h3)])} : reg892));
              reg1657 = {reg1623,
                  $unsigned(($signed((reg1651 ?
                      reg1622 : reg893)) == (+$unsigned(wire97))))};
              reg1658 = reg849;
            end
          else
            begin
              reg1659 <= reg1624;
              reg1660 <= $unsigned($signed({((wire1619 >= reg1645) >> (reg804 ?
                      reg853 : (8'hb3)))}));
              reg1661 <= ((~&reg812) ?
                  (reg878 - (({(8'had)} ?
                          (reg1624 && reg1660) : (reg1639 ?
                              reg1643 : reg1654)) ?
                      (8'hba) : (reg854[(3'h7):(3'h7)] >>> (reg811 ?
                          wire100 : reg1626)))) : (reg1635 >> reg1642[(2'h3):(2'h2)]));
              reg1662 <= $unsigned(reg868);
              reg1663 = (((8'ha0) || (8'hb4)) ?
                  $signed(reg843) : $signed((^~$signed((|reg1656)))));
            end
        end
    end
  assign wire1664 = (((8'ha3) != (reg1661[(4'h9):(3'h6)] ?
                        $signed(reg849) : wire99)) == ((reg817 ?
                            $signed($unsigned(reg829)) : ($unsigned(wire1621) ?
                                $unsigned(wire98) : (reg1644 == (8'hbd)))) ?
                        $unsigned($signed({reg865,
                            wire97})) : (wire98 <<< reg806)));
  assign wire1665 = reg874[(3'h5):(3'h4)];
  module1227 #() modinst1667 (wire1666, clk, reg826, reg865, reg874, wire100, reg861);
  always
    @(posedge clk) begin
      reg1668 = (^{{$unsigned(reg1660[(1'h1):(1'h1)]),
              ((7'h40) ? $unsigned(reg807) : wire98[(1'h0):(1'h0)])}});
    end
  assign wire1669 = {wire1664[(2'h2):(1'h0)]};
  always
    @(posedge clk) begin
      reg1670 = (8'ha2);
      if (((~^$signed($signed(reg1640[(1'h1):(1'h0)]))) ?
          $unsigned(reg890) : wire98[(4'ha):(3'h7)]))
        begin
          for (forvar1671 = (1'h0); (forvar1671 < (1'h0)); forvar1671 = (forvar1671 + (1'h1)))
            begin
              reg1672 = ((reg1670 ^~ (8'hb5)) ?
                  wire96[(3'h6):(2'h3)] : $unsigned(((-$signed(wire102)) & (!(reg861 * reg1624)))));
              reg1673 <= $unsigned(reg1661[(4'hb):(4'hb)]);
              reg1674 <= ($unsigned(reg840) ? reg1640 : reg852[(1'h1):(1'h1)]);
              reg1675 = (reg885[(1'h1):(1'h1)] ?
                  reg874[(4'hf):(4'ha)] : ($unsigned(reg1673) + $signed($signed($signed((8'hb4))))));
              reg1676 <= ((-{$unsigned((reg806 ?
                      forvar1671 : wire102))}) >>> $unsigned((($signed((7'h44)) - $unsigned(wire98)) <<< (reg854 ?
                  $unsigned((8'ha8)) : (~reg1662)))));
            end
          reg1677 <= $unsigned({(reg853 || (8'hb4)), reg832});
        end
      else
        begin
          for (forvar1671 = (1'h0); (forvar1671 < (1'h0)); forvar1671 = (forvar1671 + (1'h1)))
            begin
              reg1672 = (^~($unsigned(((reg887 ^ reg876) ?
                  (reg1624 ^ wire97) : (8'hb6))) ^~ {reg886}));
              reg1673 <= wire802;
            end
          reg1674 <= $signed((reg1662 ?
              (reg888[(4'he):(3'h6)] ?
                  $unsigned((~|reg810)) : {((7'h49) - reg804),
                      $unsigned((8'ha2))}) : $signed($unsigned(reg1676[(4'hd):(4'h9)]))));
        end
      for (forvar1678 = (1'h0); (forvar1678 < (3'h4)); forvar1678 = (forvar1678 + (1'h1)))
        begin
          if ((({reg804} ?
                  (((!(8'hb3)) >= $signed(wire802)) ?
                      $unsigned(reg887) : $unsigned((~&reg1674))) : ({(reg832 ?
                              (7'h4a) : (8'hbf))} ?
                      (8'ha8) : reg847[(2'h3):(1'h1)])) ?
              wire1619[(4'hb):(3'h6)] : (-$unsigned((reg1675 ?
                  $unsigned(reg1650) : (!reg829))))))
            begin
              reg1679 = (($signed((((8'hac) < reg887) ?
                          $unsigned(reg819) : ((8'ha6) ? wire1621 : reg876))) ?
                      $signed(($unsigned(reg1638) ?
                          $unsigned(reg1640) : ((8'h9e) - reg853))) : reg1649) ?
                  reg1638[(2'h3):(1'h1)] : reg888[(4'ha):(3'h7)]);
              reg1680 = (~|(|reg1662[(3'h4):(2'h2)]));
              reg1681 = (($signed((((8'haf) <<< reg811) - reg805)) | $unsigned($unsigned($unsigned(reg804)))) ~^ $signed(({(7'h45),
                  reg869[(1'h0):(1'h0)]} && ((reg869 ?
                  reg1673 : reg1677) || reg878))));
              reg1682 <= ((+((7'h48) | ($unsigned(reg829) ?
                  reg811[(2'h3):(1'h1)] : reg829))) - $signed(reg878[(4'ha):(4'ha)]));
              reg1683 = (&reg858[(1'h0):(1'h0)]);
            end
          else
            begin
              reg1679 = $unsigned(reg1626);
              reg1682 <= {reg1661[(4'he):(2'h2)], (~forvar1671[(1'h1):(1'h1)])};
            end
          reg1684 = reg1674;
          if (reg874)
            begin
              reg1685 = (|(!(reg878[(2'h3):(1'h1)] ?
                  ($signed(reg869) ?
                      (!reg1679) : (reg875 >> reg1679)) : $unsigned($signed(reg821)))));
              reg1686 = ($signed($unsigned(((reg1676 >> reg1683) || {reg854,
                  (7'h49)}))) << reg1659);
            end
          else
            begin
              reg1687 <= $signed(wire97);
              reg1688 <= $signed($unsigned(reg851[(4'hd):(2'h3)]));
              reg1689 <= (^~{$unsigned((^~reg852))});
              reg1690 = $unsigned((~(&(reg1675 <<< (~reg804)))));
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed((~^(~^$signed($unsigned(reg892))))))
        begin
          for (forvar1691 = (1'h0); (forvar1691 < (3'h4)); forvar1691 = (forvar1691 + (1'h1)))
            begin
              reg1692 <= $unsigned((reg1654 ?
                  $unsigned(wire800[(3'h6):(3'h6)]) : ({$signed(forvar1691)} ?
                      $unsigned(reg852[(3'h7):(3'h6)]) : $signed({reg876}))));
              reg1693 <= (|(($unsigned($unsigned((8'haf))) ?
                  (~&$signed(reg876)) : (+$unsigned(reg813))) >>> $signed(($signed((8'hbd)) ?
                  (reg859 ? wire1666 : reg1659) : (reg840 != reg849)))));
              reg1694 = ((7'h45) ?
                  (reg1623 ^ (reg807 || ((^~reg847) << $unsigned(reg889)))) : $unsigned({reg1649,
                      (~(~^reg875))}));
              reg1695 = $signed(reg855);
              reg1696 <= ((~&$signed(reg1640[(4'h8):(1'h0)])) ?
                  reg887[(1'h1):(1'h0)] : wire1664);
            end
          reg1697 <= ((~^((-(reg846 != wire1621)) && (reg1636[(2'h2):(1'h0)] ?
                  {reg1649, reg877} : reg1650[(2'h3):(2'h3)]))) ?
              $signed($signed((reg810 == $signed(reg1644)))) : ((~&$unsigned({wire800,
                      reg1623})) ?
                  (reg883 ?
                      (~|$unsigned(reg893)) : $signed($signed(reg1689))) : ($signed($signed((8'had))) ?
                      $signed($unsigned(reg821)) : $unsigned(reg810))));
          reg1698 = ($signed(reg863) + (8'h9d));
        end
      else
        begin
          reg1691 = $unsigned(($signed(($signed(wire1619) >= {reg891,
              reg875})) ~^ $signed(wire97)));
          for (forvar1692 = (1'h0); (forvar1692 < (1'h0)); forvar1692 = (forvar1692 + (1'h1)))
            begin
              reg1694 = reg817;
              reg1695 = $signed((|(-reg876[(5'h13):(5'h13)])));
              reg1698 = reg1689[(1'h0):(1'h0)];
              reg1699 = wire96[(3'h5):(3'h5)];
              reg1700 <= $unsigned((reg807 >> $signed(((wire98 && reg847) >>> reg874[(4'hf):(1'h1)]))));
            end
          reg1701 <= $signed({$unsigned(({wire102} ?
                  ((8'hab) | reg874) : ((8'haf) >= (7'h46)))),
              $unsigned(reg1682)});
          reg1702 = ($unsigned(reg829) <= $signed({({reg889} ~^ $unsigned(wire802))}));
          for (forvar1703 = (1'h0); (forvar1703 < (2'h2)); forvar1703 = (forvar1703 + (1'h1)))
            begin
              reg1704 <= $signed((^(((wire802 ? reg1633 : reg1698) | (7'h47)) ?
                  (7'h40) : $unsigned(reg893[(4'hd):(3'h4)]))));
              reg1705 <= $signed((!(((~|reg1698) | $unsigned(reg1687)) * $signed((7'h40)))));
            end
        end
      if ((8'had))
        begin
          reg1706 = reg1705;
          for (forvar1707 = (1'h0); (forvar1707 < (1'h0)); forvar1707 = (forvar1707 + (1'h1)))
            begin
              reg1708 <= {$unsigned($signed($unsigned(reg889)))};
            end
          for (forvar1709 = (1'h0); (forvar1709 < (1'h0)); forvar1709 = (forvar1709 + (1'h1)))
            begin
              reg1710 = $unsigned(($signed($unsigned(forvar1692[(2'h2):(1'h0)])) ?
                  $signed($signed(reg877[(3'h4):(3'h4)])) : ((reg1677 ?
                          wire1665[(5'h16):(5'h10)] : $signed(reg1673)) ?
                      reg1689 : (+{reg832, reg1697}))));
            end
          reg1711 <= {reg1623};
          for (forvar1712 = (1'h0); (forvar1712 < (1'h0)); forvar1712 = (forvar1712 + (1'h1)))
            begin
              reg1713 = $unsigned($unsigned(((reg878 * (reg1702 ?
                  (8'ha3) : reg1700)) <<< ({reg1649} ?
                  $unsigned(reg890) : {reg1706}))));
              reg1714 = (~&(8'ha3));
              reg1715 = (~^($unsigned(($unsigned(reg1700) ?
                      $signed(reg1708) : $signed(reg1654))) ?
                  (reg807 ?
                      (reg1662 ?
                          reg804 : (reg1662 ?
                              wire97 : reg1660)) : reg1699) : ($signed((reg1702 >>> reg1688)) ?
                      reg865[(4'h9):(3'h6)] : reg869[(4'h9):(3'h4)])));
              reg1716 <= $unsigned((reg807 ^ (^({reg1661} ?
                  reg1689 : $unsigned(reg1714)))));
            end
        end
      else
        begin
          reg1707 <= reg1676[(3'h5):(1'h1)];
          reg1709 = ($signed(reg877[(3'h5):(2'h2)]) << ((~^(reg886[(4'he):(3'h5)] ?
                  (~&reg805) : $unsigned(reg1716))) ?
              (reg1654 > reg832[(3'h4):(2'h2)]) : (&($signed(reg1715) ?
                  $signed((8'hbb)) : {reg805, reg1699}))));
          reg1710 = ((reg1689 <<< reg1640[(3'h7):(2'h3)]) ?
              $unsigned(($unsigned((reg1714 ?
                  reg805 : reg806)) || $unsigned((reg1640 | wire800)))) : $signed(reg1698[(2'h3):(2'h3)]));
          if (((($signed((~reg865)) >> (reg812 ^~ (&reg843))) ?
                  (!(~&reg886)) : reg1638) ?
              {$signed((reg1716 ? $unsigned(reg1649) : reg840)),
                  (|(((8'h9f) ? reg887 : reg876) ?
                      (~&(8'hab)) : $signed(reg804)))} : ({$unsigned(reg1626),
                      {(reg849 + reg1633)}} ?
                  (reg1702 ?
                      $unsigned(reg1709[(3'h5):(1'h1)]) : $signed((!reg1654))) : ((8'h9e) & (^(reg876 ?
                      reg810 : reg1711))))))
            begin
              reg1712 = (~(-reg876));
            end
          else
            begin
              reg1712 = $signed(($unsigned((wire100 ?
                  reg1662 : {reg1655})) >> $signed($unsigned((reg891 ~^ reg1688)))));
            end
          reg1713 = reg1677[(4'hc):(4'hb)];
        end
    end
  assign wire1717 = ($unsigned($unsigned(reg1649)) && $unsigned((reg1638[(5'h14):(3'h6)] ?
                        ({reg1697, reg868} ?
                            (reg1644 ?
                                (8'hb1) : reg847) : wire1664) : ((reg830 && wire101) ?
                            ((8'hac) ?
                                wire802 : reg861) : $unsigned(reg1687)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module896  (y, clk, wire897, wire898, wire899, wire900);
  output wire [(32'hd2b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h18):(1'h0)] wire897;
  input wire [(4'ha):(1'h0)] wire898;
  input wire signed [(4'he):(1'h0)] wire899;
  input wire [(5'h10):(1'h0)] wire900;
  wire signed [(5'h12):(1'h0)] wire1617;
  wire [(5'h11):(1'h0)] wire1526;
  wire [(4'hd):(1'h0)] wire1494;
  wire [(4'hd):(1'h0)] wire1492;
  wire [(4'h9):(1'h0)] wire901;
  wire signed [(4'hd):(1'h0)] wire902;
  wire [(5'h15):(1'h0)] wire1066;
  wire [(5'h18):(1'h0)] wire1069;
  wire signed [(5'h18):(1'h0)] wire1087;
  wire [(4'hb):(1'h0)] wire1088;
  wire [(2'h3):(1'h0)] wire1089;
  wire signed [(4'hb):(1'h0)] wire1212;
  wire signed [(4'hb):(1'h0)] wire1213;
  wire [(2'h3):(1'h0)] wire1226;
  wire signed [(4'hd):(1'h0)] wire1453;
  reg signed [(5'h12):(1'h0)] reg1524 = (1'h0);
  reg [(5'h16):(1'h0)] reg1523 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1522 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1520 = (1'h0);
  reg [(3'h5):(1'h0)] reg1519 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1517 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1511 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1516 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1515 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1513 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1512 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1508 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1506 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1503 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1502 = (1'h0);
  reg [(5'h18):(1'h0)] reg1501 = (1'h0);
  reg [(2'h3):(1'h0)] reg1499 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1496 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1490 = (1'h0);
  reg [(4'hc):(1'h0)] reg1489 = (1'h0);
  reg [(5'h15):(1'h0)] reg1487 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1486 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1480 = (1'h0);
  reg [(2'h3):(1'h0)] reg1478 = (1'h0);
  reg [(4'hc):(1'h0)] reg1477 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1476 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1474 = (1'h0);
  reg [(5'h15):(1'h0)] reg1472 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1471 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1470 = (1'h0);
  reg [(3'h4):(1'h0)] reg1467 = (1'h0);
  reg [(2'h3):(1'h0)] reg1464 = (1'h0);
  reg [(2'h3):(1'h0)] reg1462 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1458 = (1'h0);
  reg [(5'h17):(1'h0)] reg1225 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1223 = (1'h0);
  reg [(5'h18):(1'h0)] reg1222 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1221 = (1'h0);
  reg [(5'h18):(1'h0)] reg1218 = (1'h0);
  reg [(4'hb):(1'h0)] reg1217 = (1'h0);
  reg [(5'h10):(1'h0)] reg1214 = (1'h0);
  reg [(4'hf):(1'h0)] reg1210 = (1'h0);
  reg [(3'h6):(1'h0)] reg1207 = (1'h0);
  reg [(3'h4):(1'h0)] reg1203 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1199 = (1'h0);
  reg [(2'h2):(1'h0)] reg1198 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1197 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1195 = (1'h0);
  reg [(5'h17):(1'h0)] reg1192 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1196 = (1'h0);
  reg [(4'h9):(1'h0)] reg1190 = (1'h0);
  reg [(5'h15):(1'h0)] reg1189 = (1'h0);
  reg [(5'h15):(1'h0)] reg1187 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1186 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1185 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1183 = (1'h0);
  reg [(5'h11):(1'h0)] reg1181 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1180 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1179 = (1'h0);
  reg [(5'h15):(1'h0)] reg1178 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1175 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1174 = (1'h0);
  reg [(4'h8):(1'h0)] reg1172 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1168 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1167 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1164 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1161 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1159 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1158 = (1'h0);
  reg [(3'h5):(1'h0)] reg1156 = (1'h0);
  reg [(5'h16):(1'h0)] reg1154 = (1'h0);
  reg [(3'h5):(1'h0)] reg1153 = (1'h0);
  reg [(5'h14):(1'h0)] reg1143 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1138 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1137 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1135 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1134 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1133 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1129 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1128 = (1'h0);
  reg [(3'h4):(1'h0)] reg1123 = (1'h0);
  reg [(5'h11):(1'h0)] reg1122 = (1'h0);
  reg [(4'hf):(1'h0)] reg1118 = (1'h0);
  reg [(5'h17):(1'h0)] reg1117 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1115 = (1'h0);
  reg [(5'h16):(1'h0)] reg1113 = (1'h0);
  reg [(5'h16):(1'h0)] reg1112 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1107 = (1'h0);
  reg [(4'hc):(1'h0)] reg1106 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1104 = (1'h0);
  reg [(4'hc):(1'h0)] reg1103 = (1'h0);
  reg [(4'h9):(1'h0)] reg1101 = (1'h0);
  reg [(4'hd):(1'h0)] reg1099 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1098 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1095 = (1'h0);
  reg [(3'h4):(1'h0)] reg1093 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1092 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1091 = (1'h0);
  reg [(5'h10):(1'h0)] reg1086 = (1'h0);
  reg [(4'hc):(1'h0)] reg1085 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1084 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1083 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1076 = (1'h0);
  reg [(5'h16):(1'h0)] reg1072 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1068 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1525 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1521 = (1'h0);
  reg [(5'h16):(1'h0)] reg1518 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1514 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1511 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1510 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1509 = (1'h0);
  reg [(5'h16):(1'h0)] reg1507 = (1'h0);
  reg [(4'hd):(1'h0)] reg1505 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1504 = (1'h0);
  reg [(3'h6):(1'h0)] reg1500 = (1'h0);
  reg [(4'he):(1'h0)] reg1498 = (1'h0);
  reg [(5'h16):(1'h0)] reg1497 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1495 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1493 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1491 = (1'h0);
  reg [(5'h12):(1'h0)] reg1488 = (1'h0);
  reg [(4'hc):(1'h0)] reg1485 = (1'h0);
  reg [(2'h2):(1'h0)] reg1484 = (1'h0);
  reg [(2'h3):(1'h0)] reg1483 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1482 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1481 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1479 = (1'h0);
  reg [(5'h17):(1'h0)] reg1475 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1473 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1469 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1468 = (1'h0);
  reg [(3'h4):(1'h0)] reg1466 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1465 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1463 = (1'h0);
  reg [(5'h16):(1'h0)] reg1461 = (1'h0);
  reg [(5'h16):(1'h0)] reg1460 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1459 = (1'h0);
  reg [(5'h15):(1'h0)] reg1457 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1456 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1455 = (1'h0);
  reg [(5'h17):(1'h0)] reg1224 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1220 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1220 = (1'h0);
  reg [(5'h10):(1'h0)] reg1219 = (1'h0);
  reg [(4'h9):(1'h0)] reg1216 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1215 = (1'h0);
  reg [(5'h14):(1'h0)] reg1211 = (1'h0);
  reg [(2'h2):(1'h0)] reg1209 = (1'h0);
  reg [(5'h18):(1'h0)] reg1208 = (1'h0);
  reg [(4'h8):(1'h0)] reg1206 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1205 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1204 = (1'h0);
  reg [(5'h13):(1'h0)] reg1202 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1201 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1200 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1185 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1195 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1194 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1193 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1192 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1191 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1188 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1184 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1182 = (1'h0);
  reg [(4'he):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1177 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1176 = (1'h0);
  reg [(5'h16):(1'h0)] reg1173 = (1'h0);
  reg [(4'hf):(1'h0)] reg1171 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1170 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1160 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1169 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1166 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1165 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1163 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1162 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1160 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1157 = (1'h0);
  reg [(4'hc):(1'h0)] reg1155 = (1'h0);
  reg [(5'h11):(1'h0)] reg1152 = (1'h0);
  reg [(5'h14):(1'h0)] reg1151 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1150 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1149 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1148 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1147 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1146 = (1'h0);
  reg [(3'h6):(1'h0)] reg1145 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1144 = (1'h0);
  reg [(4'hb):(1'h0)] reg1142 = (1'h0);
  reg [(4'hc):(1'h0)] reg1141 = (1'h0);
  reg [(4'hf):(1'h0)] reg1140 = (1'h0);
  reg [(3'h4):(1'h0)] reg1139 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1122 = (1'h0);
  reg [(5'h10):(1'h0)] reg1136 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1132 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1131 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1130 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1127 = (1'h0);
  reg [(4'hb):(1'h0)] reg1126 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1125 = (1'h0);
  reg [(4'hb):(1'h0)] reg1124 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1121 = (1'h0);
  reg [(5'h10):(1'h0)] reg1120 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1119 = (1'h0);
  reg [(4'hd):(1'h0)] reg1116 = (1'h0);
  reg [(5'h10):(1'h0)] reg1114 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1110 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1106 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1104 = (1'h0);
  reg [(4'h9):(1'h0)] reg1111 = (1'h0);
  reg [(4'h9):(1'h0)] reg1110 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1109 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1108 = (1'h0);
  reg [(5'h14):(1'h0)] reg1105 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1102 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1100 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1097 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1094 = (1'h0);
  reg [(5'h17):(1'h0)] reg1090 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1082 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1081 = (1'h0);
  reg [(5'h16):(1'h0)] reg1080 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1079 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1078 = (1'h0);
  reg [(2'h2):(1'h0)] reg1077 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1075 = (1'h0);
  reg [(4'he):(1'h0)] reg1074 = (1'h0);
  reg [(3'h7):(1'h0)] reg1073 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1071 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1070 = (1'h0);
  assign y = {wire1617,
                 wire1526,
                 wire1494,
                 wire1492,
                 wire901,
                 wire902,
                 wire1066,
                 wire1069,
                 wire1087,
                 wire1088,
                 wire1089,
                 wire1212,
                 wire1213,
                 wire1226,
                 wire1453,
                 reg1524,
                 reg1523,
                 reg1522,
                 reg1520,
                 reg1519,
                 reg1517,
                 reg1511,
                 reg1516,
                 reg1515,
                 reg1513,
                 reg1512,
                 reg1508,
                 reg1506,
                 reg1503,
                 reg1502,
                 reg1501,
                 reg1499,
                 reg1496,
                 reg1490,
                 reg1489,
                 reg1487,
                 reg1486,
                 reg1480,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1474,
                 reg1472,
                 reg1471,
                 reg1470,
                 reg1467,
                 reg1464,
                 reg1462,
                 reg1458,
                 reg1225,
                 reg1223,
                 reg1222,
                 reg1221,
                 reg1218,
                 reg1217,
                 reg1214,
                 reg1210,
                 reg1207,
                 reg1203,
                 reg1199,
                 reg1198,
                 reg1197,
                 reg1195,
                 reg1192,
                 reg1196,
                 reg1190,
                 reg1189,
                 reg1187,
                 reg1186,
                 reg1185,
                 reg1183,
                 reg1181,
                 reg1180,
                 reg1179,
                 reg1178,
                 reg1175,
                 reg1174,
                 reg1172,
                 reg1168,
                 reg1167,
                 reg1164,
                 reg1161,
                 reg1159,
                 reg1158,
                 reg1156,
                 reg1154,
                 reg1153,
                 reg1143,
                 reg1138,
                 reg1137,
                 reg1135,
                 reg1134,
                 reg1133,
                 reg1129,
                 reg1128,
                 reg1123,
                 reg1122,
                 reg1118,
                 reg1117,
                 reg1115,
                 reg1113,
                 reg1112,
                 reg1107,
                 reg1106,
                 reg1104,
                 reg1103,
                 reg1101,
                 reg1099,
                 reg1098,
                 reg1095,
                 reg1093,
                 reg1092,
                 reg1091,
                 reg1086,
                 reg1085,
                 reg1084,
                 reg1083,
                 reg1076,
                 reg1072,
                 reg1068,
                 reg1525,
                 reg1521,
                 reg1518,
                 reg1514,
                 forvar1511,
                 reg1510,
                 reg1509,
                 reg1507,
                 reg1505,
                 reg1504,
                 reg1500,
                 reg1498,
                 reg1497,
                 forvar1495,
                 reg1493,
                 reg1491,
                 reg1488,
                 reg1485,
                 reg1484,
                 reg1483,
                 reg1482,
                 forvar1481,
                 reg1479,
                 reg1475,
                 reg1473,
                 reg1469,
                 forvar1468,
                 reg1466,
                 reg1465,
                 reg1463,
                 reg1461,
                 reg1460,
                 reg1459,
                 reg1457,
                 forvar1456,
                 forvar1455,
                 reg1224,
                 forvar1220,
                 reg1220,
                 reg1219,
                 reg1216,
                 reg1215,
                 reg1211,
                 reg1209,
                 reg1208,
                 reg1206,
                 forvar1205,
                 forvar1204,
                 reg1202,
                 forvar1201,
                 forvar1200,
                 forvar1185,
                 forvar1195,
                 reg1194,
                 reg1193,
                 forvar1192,
                 reg1191,
                 reg1188,
                 reg1184,
                 reg1182,
                 reg1176,
                 reg1177,
                 forvar1176,
                 reg1173,
                 reg1171,
                 forvar1170,
                 reg1160,
                 reg1169,
                 forvar1166,
                 reg1165,
                 reg1163,
                 reg1162,
                 forvar1160,
                 forvar1157,
                 reg1155,
                 reg1152,
                 reg1151,
                 reg1150,
                 reg1149,
                 forvar1148,
                 forvar1147,
                 reg1146,
                 reg1145,
                 reg1144,
                 reg1142,
                 reg1141,
                 reg1140,
                 reg1139,
                 forvar1122,
                 reg1136,
                 reg1132,
                 reg1131,
                 reg1130,
                 reg1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1121,
                 reg1120,
                 reg1119,
                 reg1116,
                 reg1114,
                 forvar1110,
                 forvar1106,
                 forvar1104,
                 reg1111,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1105,
                 reg1102,
                 forvar1100,
                 reg1097,
                 reg1096,
                 reg1094,
                 reg1090,
                 reg1082,
                 reg1081,
                 reg1080,
                 reg1079,
                 forvar1078,
                 reg1077,
                 reg1075,
                 reg1074,
                 reg1073,
                 forvar1071,
                 reg1070,
                 (1'h0)};
  assign wire901 = ((~|((~^wire897[(2'h3):(2'h3)]) != ($unsigned(wire898) >> (wire899 - wire898)))) ?
                       {$unsigned((wire899[(3'h7):(3'h4)] ?
                               $signed((7'h48)) : $unsigned((8'hb6)))),
                           wire897} : {((-$unsigned(wire898)) + (wire898[(1'h1):(1'h0)] ?
                               (^wire897) : $unsigned(wire897))),
                           $signed(($unsigned(wire898) ?
                               wire897 : (wire898 ? wire899 : wire897)))});
  assign wire902 = wire899;
  module903 #() modinst1067 (wire1066, clk, wire902, wire899, wire897, wire898);
  always
    @(posedge clk) begin
      reg1068 <= ((+$unsigned((((8'hb1) < (8'h9f)) && wire899))) ?
          $signed(wire897[(1'h1):(1'h0)]) : (~|$signed(wire898)));
    end
  assign wire1069 = $signed($unsigned(($signed(wire897[(4'h8):(1'h1)]) ?
                        ((wire900 ? wire1066 : wire900) ?
                            (wire898 ?
                                wire897 : wire902) : $unsigned(wire899)) : ($signed((7'h42)) ?
                            (&reg1068) : (|(8'hab))))));
  always
    @(posedge clk) begin
      reg1070 = ((&(((reg1068 ? wire902 : reg1068) != (-wire1069)) ?
              ($signed(wire898) ?
                  $unsigned(reg1068) : (wire1069 && wire897)) : $unsigned({wire899}))) ?
          (^~$signed($signed($unsigned(wire902)))) : $unsigned(wire902));
      for (forvar1071 = (1'h0); (forvar1071 < (3'h4)); forvar1071 = (forvar1071 + (1'h1)))
        begin
          if ((wire898[(2'h3):(1'h1)] ?
              ((!(~|((8'hb1) ~^ wire899))) ~^ {wire902[(4'hd):(3'h6)],
                  reg1070[(4'hb):(4'hb)]}) : $signed((wire901 ?
                  $unsigned($signed(wire1069)) : $signed(wire1069[(4'hf):(3'h7)])))))
            begin
              reg1072 <= (wire1069[(3'h5):(1'h1)] ?
                  (reg1068[(2'h2):(2'h2)] ?
                      (~|($signed(wire900) ?
                          wire1069[(3'h7):(3'h5)] : $unsigned(wire1066))) : (wire899 ?
                          $unsigned(wire1069[(5'h15):(3'h4)]) : (!wire899[(4'hc):(4'ha)]))) : $signed(((^$unsigned(wire901)) <<< ($signed(forvar1071) ?
                      $signed(wire897) : (reg1070 ? wire900 : (7'h49))))));
            end
          else
            begin
              reg1073 = (forvar1071[(4'hd):(2'h2)] ?
                  (wire902 ?
                      reg1070 : wire898[(4'ha):(2'h3)]) : {(|((wire901 >= (8'ha4)) == (reg1068 ?
                          wire899 : reg1068))),
                      (~|$unsigned(forvar1071))});
            end
          reg1074 = ($unsigned($unsigned(reg1070[(5'h10):(4'he)])) ?
              {wire899} : ($unsigned((((7'h43) > wire901) >>> wire899)) >> (((!reg1072) ?
                      wire897 : (^wire1069)) ?
                  (wire900[(4'ha):(2'h3)] ^ {wire899}) : {$unsigned(wire899)})));
          if ((^$unsigned(wire1069)))
            begin
              reg1075 = wire901;
              reg1076 <= $signed(reg1068);
            end
          else
            begin
              reg1075 = wire900;
            end
        end
      reg1077 = $signed((($unsigned($signed(reg1072)) == {(wire900 == wire902)}) ?
          ({$signed((8'hb4)), wire897[(4'hc):(4'hb)]} ?
              (((8'h9e) << wire901) ?
                  $unsigned(reg1070) : reg1068) : $signed(wire899)) : {$unsigned((wire902 << wire1069)),
              $unsigned((reg1068 > reg1075))}));
      for (forvar1078 = (1'h0); (forvar1078 < (2'h3)); forvar1078 = (forvar1078 + (1'h1)))
        begin
          reg1079 = $unsigned({((~^(^~forvar1078)) ?
                  {reg1072} : reg1073[(1'h1):(1'h1)])});
          if (((^{wire899[(4'h8):(3'h7)],
              ((wire1069 ?
                  reg1079 : reg1068) > reg1079)}) * $unsigned(wire902[(2'h2):(1'h1)])))
            begin
              reg1080 = reg1068[(1'h0):(1'h0)];
              reg1081 = ((($unsigned(wire899) ?
                  {$unsigned((8'ha3))} : ((reg1074 ?
                      reg1079 : reg1070) - (8'hb0))) || reg1076[(3'h4):(1'h0)]) | $signed(reg1077[(2'h2):(1'h1)]));
              reg1082 = wire902;
            end
          else
            begin
              reg1083 <= $unsigned({(^~(^~{wire900})),
                  ($unsigned((forvar1071 ? (8'hba) : reg1082)) ?
                      wire900[(3'h6):(3'h5)] : ((reg1073 ? reg1074 : reg1070) ?
                          reg1075 : (reg1075 >= (8'hb7))))});
              reg1084 <= $unsigned((($signed((&reg1079)) >= $signed($signed(wire898))) ?
                  wire902[(3'h5):(3'h5)] : {($signed(reg1068) * wire1066[(4'hd):(3'h5)]),
                      {$signed(reg1070)}}));
              reg1085 <= ($signed((-$signed(reg1079))) ?
                  reg1079[(2'h2):(2'h2)] : (~&wire902));
              reg1086 <= {reg1076[(2'h2):(1'h0)],
                  $unsigned(wire898[(4'h8):(3'h4)])};
            end
        end
    end
  assign wire1087 = $unsigned($unsigned(((~|(&reg1072)) & (wire901[(3'h7):(1'h0)] <<< (~|reg1072)))));
  assign wire1088 = (((~^reg1072) ? reg1083 : $signed(reg1076)) ?
                        $signed($signed($unsigned((8'ha4)))) : ({{wire1069,
                                (wire1069 ?
                                    reg1076 : wire897)}} >>> (|({wire902,
                                (8'haa)} ?
                            reg1068 : (wire1087 > reg1084)))));
  assign wire1089 = (reg1083 >> $unsigned(reg1086));
  always
    @(posedge clk) begin
      if (($unsigned(($signed(wire901[(4'h8):(3'h7)]) ?
              reg1076 : {$signed(wire902)})) ?
          wire898[(3'h6):(3'h6)] : ($unsigned({wire1066[(4'he):(4'hc)],
              (+reg1086)}) <= $unsigned($signed((+(8'h9d)))))))
        begin
          reg1090 = {($unsigned($unsigned((reg1076 ? wire1069 : reg1086))) ?
                  $unsigned(((+wire899) ^ ((7'h49) & wire900))) : (wire901[(1'h0):(1'h0)] == ($unsigned(wire1066) || (+wire902)))),
              $signed(($unsigned((reg1076 != (8'h9e))) ?
                  ((reg1068 <<< wire902) <<< {(8'hbc)}) : ({wire901} - $unsigned(reg1085))))};
        end
      else
        begin
          reg1091 <= (8'h9d);
          reg1092 <= ({((~&(8'hba)) <<< {$signed(wire897)})} <<< wire897);
          reg1093 <= ((~^wire1088[(1'h0):(1'h0)]) <<< (reg1092 ?
              reg1085[(2'h3):(1'h0)] : $signed(wire900)));
          if (($unsigned($unsigned({(wire902 ? wire899 : wire1066),
              ((8'h9c) > reg1084)})) ~^ $signed(wire897[(5'h11):(4'he)])))
            begin
              reg1094 = reg1084[(5'h13):(3'h4)];
              reg1095 <= $unsigned($unsigned(reg1083));
              reg1096 = wire899[(4'h9):(3'h6)];
              reg1097 = (8'hb2);
            end
          else
            begin
              reg1095 <= $signed($signed((($signed(reg1097) ?
                  reg1090[(3'h5):(2'h3)] : reg1084[(5'h17):(4'hc)]) >> (-{wire897}))));
              reg1096 = (^~{wire1088[(4'hb):(1'h0)], wire1066[(3'h4):(1'h0)]});
              reg1098 <= (^~(7'h4a));
              reg1099 <= wire899;
            end
        end
      for (forvar1100 = (1'h0); (forvar1100 < (3'h4)); forvar1100 = (forvar1100 + (1'h1)))
        begin
          reg1101 <= (~^reg1083);
          reg1102 = reg1097;
          reg1103 <= ($signed($signed($signed(reg1091))) ?
              reg1072[(5'h10):(4'hf)] : (&((~|(~^reg1096)) <= {$unsigned((8'h9c))})));
        end
      if ((~^reg1101))
        begin
          if ((reg1101[(2'h3):(2'h3)] ?
              (^$signed(wire1069)) : {{(!(~reg1093))}}))
            begin
              reg1104 <= reg1086[(4'hf):(4'hf)];
              reg1105 = $unsigned((8'ha9));
              reg1106 <= $unsigned((~|(reg1068 ?
                  ($signed(reg1093) ^ (reg1093 << reg1104)) : {$unsigned((7'h48)),
                      reg1076})));
              reg1107 <= ($signed(reg1096[(4'hc):(4'ha)]) ?
                  $unsigned(((~&(reg1106 && (8'hab))) + (+wire1087[(3'h6):(3'h6)]))) : (~$signed($signed($unsigned(reg1083)))));
            end
          else
            begin
              reg1104 <= $signed(({(reg1068 ?
                      $signed(wire1069) : $signed(wire899)),
                  $signed($signed(reg1076))} * (reg1083[(2'h2):(1'h0)] ?
                  ((reg1105 | wire899) >= $signed(reg1105)) : reg1107)));
              reg1105 = (($unsigned(reg1083[(4'hb):(4'h8)]) > $unsigned({(reg1068 ?
                          reg1099 : reg1091),
                      $unsigned(wire899)})) ?
                  (reg1102[(4'hb):(4'h9)] | ($signed((reg1092 != (7'h46))) ^~ reg1099[(4'ha):(1'h0)])) : ((reg1068[(2'h3):(2'h3)] > (reg1090 << $signed(wire900))) ?
                      (^~(~&(forvar1100 ?
                          wire902 : wire1087))) : $signed((wire899[(3'h4):(3'h4)] ?
                          wire1066 : reg1091))));
              reg1108 = {$unsigned(($signed((reg1092 == reg1098)) & (((8'ha2) ?
                          reg1084 : reg1076) ?
                      $unsigned(reg1101) : $signed(forvar1100))))};
              reg1109 = reg1098[(1'h0):(1'h0)];
            end
          reg1110 = (($unsigned($unsigned((8'ha3))) * $unsigned($signed((reg1109 || reg1093)))) && (({reg1090[(3'h7):(3'h6)],
                  (-wire898)} ?
              $signed({reg1107}) : ((^reg1099) == forvar1100)) < (~&wire1089[(2'h3):(2'h2)])));
          reg1111 = ($signed($signed((~$unsigned(reg1097)))) << $unsigned((~^reg1091)));
          reg1112 <= ($unsigned($unsigned((^forvar1100))) ?
              (^~(((reg1093 ? reg1102 : reg1103) ^ (reg1096 <<< reg1093)) ?
                  (reg1110 & reg1085) : reg1102[(2'h2):(1'h0)])) : $signed(reg1094));
          reg1113 <= (wire901 ?
              reg1093[(1'h1):(1'h0)] : (($unsigned($signed(reg1090)) ?
                      {reg1072,
                          (wire1087 >> (8'ha2))} : ((8'hb3) <<< (^~reg1093))) ?
                  reg1068[(4'h8):(1'h1)] : wire1066));
        end
      else
        begin
          for (forvar1104 = (1'h0); (forvar1104 < (1'h0)); forvar1104 = (forvar1104 + (1'h1)))
            begin
              reg1105 = $unsigned((($unsigned((~|wire1066)) ?
                  ($unsigned(reg1090) ?
                      $unsigned(wire901) : reg1090[(4'h9):(3'h7)]) : ($signed(reg1095) & (~^wire1087))) >>> $unsigned((^(!reg1085)))));
            end
          for (forvar1106 = (1'h0); (forvar1106 < (3'h4)); forvar1106 = (forvar1106 + (1'h1)))
            begin
              reg1108 = $unsigned(wire1089);
              reg1109 = (&((($signed(reg1113) ?
                      $unsigned(wire897) : $unsigned(reg1109)) ?
                  (^~(forvar1104 ?
                      wire1089 : forvar1100)) : $unsigned($signed(reg1093))) > (!reg1068[(1'h1):(1'h0)])));
            end
          for (forvar1110 = (1'h0); (forvar1110 < (1'h1)); forvar1110 = (forvar1110 + (1'h1)))
            begin
              reg1112 <= {$signed({(^(reg1101 | reg1106)),
                      ((wire897 ? wire1069 : reg1103) <<< $unsigned(reg1091))}),
                  $signed($unsigned(((wire897 + wire1088) ?
                      (|(7'h47)) : reg1093[(2'h2):(2'h2)])))};
              reg1113 <= $signed($unsigned(($signed((8'hb7)) ?
                  ({wire1069, reg1083} ?
                      $signed(reg1101) : $unsigned(reg1095)) : ($unsigned(reg1096) ?
                      (~&reg1107) : (wire899 ? reg1097 : wire1089)))));
              reg1114 = reg1110[(4'h9):(4'h8)];
              reg1115 <= (wire1066 >> $unsigned(({reg1099[(3'h6):(3'h6)],
                      (reg1104 + wire1087)} ?
                  $unsigned((wire1069 ?
                      reg1112 : reg1099)) : wire1089[(2'h2):(2'h2)])));
            end
          if (($unsigned(reg1105[(4'he):(4'h8)]) ?
              {$signed($unsigned($signed(wire1087))),
                  (reg1114[(4'hb):(2'h2)] > reg1098[(2'h3):(2'h3)])} : $unsigned(wire899)))
            begin
              reg1116 = wire897[(5'h17):(3'h5)];
              reg1117 <= reg1072[(4'hc):(2'h2)];
              reg1118 <= $unsigned(((^~(~^$signed(reg1076))) >= (+(7'h41))));
            end
          else
            begin
              reg1116 = (($signed(reg1084[(4'h9):(2'h2)]) ?
                      (^reg1113) : ({(-reg1102)} != $unsigned((reg1118 < forvar1106)))) ?
                  ((reg1076 ?
                          $signed((reg1097 ?
                              (8'ha5) : reg1113)) : $unsigned(reg1072)) ?
                      (((~|reg1113) ?
                          (^~reg1111) : (reg1118 ?
                              wire1087 : reg1112)) == $unsigned({reg1103,
                          reg1107})) : (($signed(reg1112) ?
                              (reg1107 != reg1105) : reg1104[(4'hf):(2'h2)]) ?
                          reg1113 : $unsigned(forvar1100))) : $unsigned(forvar1100));
              reg1119 = reg1118[(3'h5):(3'h5)];
              reg1120 = $unsigned($signed(wire899));
            end
          reg1121 = (|$unsigned(($unsigned(reg1109) - $unsigned((reg1083 * (8'ha7))))));
        end
      if ($signed(($unsigned((^~$unsigned(reg1121))) ?
          reg1112[(3'h4):(1'h0)] : ((reg1110 <= reg1119) ~^ ({(8'haa),
              reg1118} * $unsigned(wire1069))))))
        begin
          if (wire1089)
            begin
              reg1122 <= (((($unsigned(wire899) >> reg1072[(3'h4):(2'h3)]) ?
                      (~&$signed((8'hbf))) : forvar1106[(3'h5):(2'h2)]) ?
                  ($signed({reg1068}) ?
                      $signed(reg1112) : reg1092) : ((reg1121 || ((8'ha1) ?
                      (8'hb3) : reg1096)) * (&(~(8'hac))))) | ($signed((8'ha3)) || $unsigned($unsigned((forvar1106 ?
                  reg1076 : wire1066)))));
              reg1123 <= (&forvar1100);
            end
          else
            begin
              reg1124 = $signed(forvar1100[(3'h5):(3'h4)]);
              reg1125 = $unsigned((reg1124[(4'ha):(3'h4)] ?
                  {(reg1113 ? wire1089 : {reg1096}),
                      $unsigned((reg1113 & reg1120))} : ({$unsigned(reg1083),
                      wire901} != {(reg1122 * reg1098)})));
              reg1126 = ((reg1106[(4'h9):(1'h1)] ?
                  (((reg1072 * (8'hbb)) + reg1104[(1'h0):(1'h0)]) ?
                      reg1072 : $signed((-wire900))) : reg1121) * ((-({(8'haf),
                          reg1076} ?
                      $signed(reg1104) : (^~reg1096))) ?
                  wire1089[(1'h1):(1'h0)] : ((reg1119[(3'h5):(2'h2)] ^~ (reg1118 ?
                      (8'h9f) : wire1089)) - $unsigned((+reg1115)))));
              reg1127 = reg1083;
            end
          reg1128 <= (reg1090 * $signed(reg1096));
          reg1129 <= reg1126[(4'hb):(4'h8)];
          reg1130 = $signed($signed(reg1094[(3'h4):(1'h0)]));
          if ((~|$unsigned((+($unsigned(reg1068) - (&reg1111))))))
            begin
              reg1131 = reg1118[(3'h4):(2'h2)];
              reg1132 = reg1124[(3'h5):(3'h5)];
              reg1133 <= (7'h4a);
              reg1134 <= $unsigned({$signed(($unsigned(wire1088) + {reg1097,
                      (8'ha7)})),
                  $unsigned(($signed(reg1083) ^ (wire1089 | wire897)))});
            end
          else
            begin
              reg1133 <= $signed($signed(({$unsigned(reg1104)} ?
                  $signed({wire899, (8'h9c)}) : reg1129[(3'h7):(3'h7)])));
              reg1134 <= forvar1100[(4'h9):(3'h7)];
              reg1135 <= ($signed($unsigned(((^(8'hb1)) >> reg1107))) && $signed({reg1076[(2'h2):(1'h0)],
                  ($unsigned(reg1098) >>> (wire1069 >= (8'ha8)))}));
              reg1136 = wire1066;
            end
        end
      else
        begin
          for (forvar1122 = (1'h0); (forvar1122 < (3'h4)); forvar1122 = (forvar1122 + (1'h1)))
            begin
              reg1123 <= $unsigned(reg1095);
              reg1128 <= reg1111[(4'h9):(3'h4)];
              reg1130 = $signed(wire902);
              reg1133 <= forvar1106[(1'h1):(1'h1)];
              reg1134 <= $unsigned((-((^reg1106) || (~^reg1099))));
            end
          if ($signed(($unsigned($unsigned(reg1122)) ?
              reg1103 : (~^$signed((reg1112 & reg1076))))))
            begin
              reg1136 = ($unsigned(wire901[(3'h7):(3'h6)]) | (|$signed((reg1118 ?
                  $unsigned(reg1098) : $signed(reg1107)))));
              reg1137 <= {forvar1104[(3'h4):(1'h0)]};
              reg1138 <= ($unsigned((^wire899)) ~^ reg1120[(1'h1):(1'h1)]);
              reg1139 = ({($signed((reg1135 & reg1086)) ?
                      wire902 : ((|reg1084) != (reg1127 | reg1137))),
                  $unsigned(reg1091)} >= $unsigned(({$unsigned(reg1103)} ?
                  forvar1110 : {$signed((7'h41))})));
              reg1140 = ($signed((^~$unsigned((wire1069 ?
                  reg1084 : reg1112)))) * $signed($unsigned(wire1089)));
            end
          else
            begin
              reg1136 = ((^~$unsigned($signed($unsigned(forvar1122)))) & reg1129[(2'h3):(1'h0)]);
              reg1139 = $unsigned(reg1130);
              reg1140 = (!{$unsigned({$signed((7'h4a))}),
                  $signed({$unsigned(reg1122)})});
            end
          if ($signed({(((reg1134 > reg1111) ^~ (~|reg1112)) ?
                  reg1125 : ((8'hb1) != reg1092)),
              reg1136}))
            begin
              reg1141 = wire899;
              reg1142 = {wire898};
            end
          else
            begin
              reg1141 = ($signed(reg1138) >= $unsigned($unsigned(((8'ha3) ?
                  {reg1110} : ((8'ha7) >>> reg1085)))));
            end
          if (({reg1106[(3'h4):(3'h4)], reg1068} >>> (reg1091[(1'h1):(1'h1)] ?
              {$unsigned((~|reg1109))} : (~^$unsigned($signed(forvar1110))))))
            begin
              reg1143 <= $unsigned((8'hbf));
              reg1144 = {$signed($signed({(~&reg1091)}))};
            end
          else
            begin
              reg1144 = $signed((~^(&$unsigned($unsigned(wire900)))));
              reg1145 = (forvar1106 < reg1134[(4'ha):(4'h9)]);
            end
        end
      reg1146 = (-reg1127[(2'h3):(1'h0)]);
    end
  always
    @(posedge clk) begin
      for (forvar1147 = (1'h0); (forvar1147 < (1'h1)); forvar1147 = (forvar1147 + (1'h1)))
        begin
          for (forvar1148 = (1'h0); (forvar1148 < (1'h0)); forvar1148 = (forvar1148 + (1'h1)))
            begin
              reg1149 = wire900;
              reg1150 = ($signed($unsigned((8'ha6))) > (wire899 ~^ $signed($signed((wire901 ~^ reg1086)))));
              reg1151 = {(reg1129[(2'h3):(2'h3)] ?
                      ((~&wire897[(4'he):(4'h9)]) ?
                          reg1123[(1'h0):(1'h0)] : {(forvar1148 ?
                                  (8'hb6) : reg1086)}) : (^$unsigned((&reg1095)))),
                  ((~|($unsigned(forvar1148) ?
                      (reg1098 << wire900) : (~&(7'h41)))) > $unsigned((~^(reg1091 ?
                      reg1068 : reg1103))))};
              reg1152 = wire898;
              reg1153 <= {$signed($unsigned(((wire898 ? forvar1148 : reg1104) ?
                      $signed(reg1134) : (+reg1085))))};
            end
          reg1154 <= (wire1087[(1'h1):(1'h0)] >>> (({$unsigned(wire1066)} ?
              $signed((8'hac)) : reg1095[(1'h0):(1'h0)]) || $signed($signed(reg1112[(2'h3):(2'h2)]))));
          reg1155 = wire902;
          reg1156 <= ((~(^(|reg1129[(3'h5):(1'h0)]))) >> $signed(reg1068[(3'h7):(3'h6)]));
        end
      for (forvar1157 = (1'h0); (forvar1157 < (2'h2)); forvar1157 = (forvar1157 + (1'h1)))
        begin
          reg1158 <= ($unsigned((reg1101 ?
              $signed({(8'hb2),
                  reg1156}) : $signed((^reg1115)))) << reg1098[(2'h3):(2'h2)]);
        end
    end
  always
    @(posedge clk) begin
      if ($signed($unsigned((~&reg1106[(1'h1):(1'h0)]))))
        begin
          reg1159 <= (-((^~$signed({reg1129})) ?
              ($unsigned(wire1088) ?
                  reg1158[(2'h2):(1'h0)] : reg1113[(3'h5):(1'h0)]) : (((~|(8'ha8)) ?
                      wire1088[(2'h2):(2'h2)] : reg1107) ?
                  ($signed(reg1153) ?
                      reg1135[(4'h9):(2'h2)] : ((8'hb2) < reg1083)) : $signed(((7'h48) ?
                      reg1137 : (8'hb2))))));
          for (forvar1160 = (1'h0); (forvar1160 < (1'h1)); forvar1160 = (forvar1160 + (1'h1)))
            begin
              reg1161 <= {{(~|(~|(!reg1159)))}};
              reg1162 = $signed($unsigned(reg1129));
              reg1163 = $signed((&(~reg1161[(5'h13):(5'h13)])));
              reg1164 <= $signed((^~(reg1134[(2'h2):(2'h2)] ?
                  {reg1098, (reg1093 ^~ reg1129)} : wire899)));
              reg1165 = reg1156[(3'h4):(1'h0)];
            end
          for (forvar1166 = (1'h0); (forvar1166 < (1'h0)); forvar1166 = (forvar1166 + (1'h1)))
            begin
              reg1167 <= $signed(($unsigned(reg1128) <<< $unsigned({(wire1069 <<< reg1076),
                  (wire900 <<< reg1091)})));
              reg1168 <= $signed($signed(((8'ha8) ?
                  reg1072[(4'h9):(3'h4)] : reg1133[(3'h5):(1'h1)])));
              reg1169 = (($unsigned(($signed(reg1101) ? reg1113 : {reg1161})) ?
                  $signed(reg1163) : (^~reg1084[(5'h10):(4'he)])) >= reg1156);
            end
        end
      else
        begin
          reg1159 <= (~|($signed(($signed(reg1159) + $signed((8'hb9)))) ?
              reg1128[(3'h6):(1'h1)] : $unsigned($unsigned(reg1161[(2'h2):(1'h1)]))));
          reg1160 = $signed((($unsigned((~^reg1113)) ?
                  reg1085[(4'ha):(4'ha)] : {reg1084[(4'ha):(2'h3)],
                      $unsigned(reg1113)}) ?
              (~&(!(-(7'h4a)))) : wire900));
          reg1162 = (~^$unsigned($signed(((+reg1161) ?
              reg1107 : (reg1085 ? reg1153 : (8'ha1))))));
        end
      if ($unsigned((&{($unsigned(reg1168) ^~ reg1135[(4'ha):(4'h9)])})))
        begin
          for (forvar1170 = (1'h0); (forvar1170 < (1'h0)); forvar1170 = (forvar1170 + (1'h1)))
            begin
              reg1171 = (-reg1168[(2'h2):(2'h2)]);
              reg1172 <= $unsigned(reg1086);
              reg1173 = {(&($unsigned(((8'h9f) << (8'haa))) ^~ $signed($unsigned(wire1088)))),
                  $unsigned(reg1128)};
              reg1174 <= $signed((8'hb6));
            end
          reg1175 <= $signed(($signed({wire899[(4'hb):(4'hb)]}) ?
              {$unsigned({reg1143, forvar1166}),
                  (^{wire1069, wire1069})} : reg1083[(3'h6):(3'h5)]));
          for (forvar1176 = (1'h0); (forvar1176 < (1'h1)); forvar1176 = (forvar1176 + (1'h1)))
            begin
              reg1177 = ((((wire899[(4'hc):(2'h2)] >> reg1162) >> wire900) >> ((+$unsigned(reg1167)) ?
                  (&(reg1129 ?
                      reg1129 : wire1066)) : reg1143)) < $signed(reg1106));
              reg1178 <= $signed(((($unsigned((8'h9f)) ?
                          (reg1072 ?
                              forvar1176 : reg1085) : ((8'had) <= forvar1176)) ?
                      {$signed(reg1153)} : $unsigned((reg1154 - wire901))) ?
                  $unsigned($unsigned((~reg1118))) : $unsigned(reg1115)));
              reg1179 <= reg1076;
              reg1180 <= reg1128[(2'h3):(2'h2)];
              reg1181 <= ((~(~|(reg1156[(3'h5):(2'h2)] ?
                  ((7'h42) < reg1143) : reg1138))) != {(8'ha2)});
            end
        end
      else
        begin
          for (forvar1170 = (1'h0); (forvar1170 < (2'h3)); forvar1170 = (forvar1170 + (1'h1)))
            begin
              reg1171 = $unsigned((~|forvar1170[(3'h5):(3'h5)]));
              reg1172 <= $signed(reg1093);
              reg1173 = reg1104[(3'h6):(3'h6)];
              reg1176 = (~^(reg1093 ?
                  (8'had) : $unsigned($unsigned(((8'ha3) ?
                      reg1115 : reg1162)))));
            end
          if (forvar1160)
            begin
              reg1177 = ((wire1087 ?
                      ($unsigned((8'hbf)) ^ wire899[(4'hb):(3'h5)]) : $unsigned(reg1153[(2'h2):(1'h0)])) ?
                  $signed($unsigned($unsigned(reg1168[(2'h3):(1'h0)]))) : wire899);
            end
          else
            begin
              reg1178 <= (&(reg1123[(3'h4):(1'h0)] == $unsigned(($signed(reg1118) ?
                  wire898 : (reg1076 * reg1163)))));
              reg1182 = reg1084;
              reg1183 <= reg1163[(2'h2):(1'h1)];
              reg1184 = $unsigned(reg1163);
            end
        end
      if (reg1134[(4'he):(4'ha)])
        begin
          reg1185 <= wire902;
          reg1186 <= (+($signed(reg1168[(2'h2):(1'h1)]) + (!$unsigned(((7'h41) & reg1159)))));
          if ((+(!(+reg1179[(5'h14):(4'hb)]))))
            begin
              reg1187 <= reg1169;
              reg1188 = (8'hb1);
            end
          else
            begin
              reg1187 <= reg1093;
              reg1188 = wire899;
              reg1189 <= ($unsigned($signed(reg1085[(3'h7):(3'h4)])) ^~ (($unsigned((reg1167 <<< reg1138)) ?
                  (~reg1129) : $signed((^reg1138))) != (^~reg1187)));
              reg1190 <= ((8'ha2) ?
                  $signed(wire902[(3'h5):(1'h0)]) : $unsigned($unsigned(forvar1160)));
              reg1191 = $signed(((8'hb0) ?
                  $unsigned(((reg1104 >> reg1093) ?
                      $unsigned(reg1169) : $unsigned(reg1162))) : $signed(((-reg1107) * (reg1068 ?
                      wire1089 : wire1088)))));
            end
          for (forvar1192 = (1'h0); (forvar1192 < (2'h2)); forvar1192 = (forvar1192 + (1'h1)))
            begin
              reg1193 = {wire897[(4'h8):(3'h6)]};
              reg1194 = (|reg1128[(2'h2):(1'h1)]);
            end
          for (forvar1195 = (1'h0); (forvar1195 < (2'h3)); forvar1195 = (forvar1195 + (1'h1)))
            begin
              reg1196 <= (+(!((~^$signed(reg1137)) ?
                  forvar1195[(5'h11):(4'hf)] : $signed((~reg1101)))));
            end
        end
      else
        begin
          for (forvar1185 = (1'h0); (forvar1185 < (2'h3)); forvar1185 = (forvar1185 + (1'h1)))
            begin
              reg1188 = reg1103[(4'ha):(3'h4)];
              reg1189 <= $signed($unsigned(reg1186[(2'h3):(2'h2)]));
              reg1191 = (+$signed((({(8'hab)} <<< reg1115[(1'h0):(1'h0)]) ^ (&reg1185))));
              reg1192 <= ((&(({reg1138} != (8'hb8)) ? reg1174 : forvar1160)) ?
                  $signed($signed($unsigned((reg1183 ?
                      reg1181 : reg1161)))) : $signed($unsigned((+{reg1185}))));
              reg1195 <= $signed($signed(reg1168[(2'h2):(1'h1)]));
            end
        end
      reg1197 <= reg1188[(4'h9):(3'h4)];
    end
  always
    @(posedge clk) begin
      reg1198 <= (reg1099 || (^wire900[(4'hc):(2'h2)]));
    end
  always
    @(posedge clk) begin
      reg1199 <= (($signed((^reg1174[(2'h3):(1'h1)])) <<< $unsigned(((^~reg1185) == $unsigned(reg1156)))) ?
          (^~$signed({(8'hbf)})) : (~|((8'haa) ?
              reg1164[(5'h16):(4'h9)] : (+(reg1086 ? reg1172 : reg1086)))));
      for (forvar1200 = (1'h0); (forvar1200 < (3'h4)); forvar1200 = (forvar1200 + (1'h1)))
        begin
          for (forvar1201 = (1'h0); (forvar1201 < (1'h1)); forvar1201 = (forvar1201 + (1'h1)))
            begin
              reg1202 = ((((~|(&reg1158)) > $unsigned($signed((8'hb8)))) ?
                  (((~|reg1192) << (reg1190 ? reg1158 : reg1192)) ?
                      ((8'hbe) ?
                          reg1164[(4'hd):(3'h5)] : reg1129[(3'h4):(3'h4)]) : (reg1167[(1'h1):(1'h1)] << $unsigned(reg1199))) : forvar1201[(2'h2):(2'h2)]) > ((((reg1084 >= reg1099) > {wire897}) ?
                  reg1112 : {$unsigned(reg1186)}) >> reg1117));
            end
          reg1203 <= {{(((reg1084 <<< (8'ha8)) ?
                      {wire1087} : wire901[(1'h0):(1'h0)]) >>> (^wire900)),
                  $unsigned((reg1199 >>> (reg1154 || wire902)))},
              {(|reg1107[(4'h8):(4'h8)]), forvar1201}};
        end
      for (forvar1204 = (1'h0); (forvar1204 < (2'h2)); forvar1204 = (forvar1204 + (1'h1)))
        begin
          for (forvar1205 = (1'h0); (forvar1205 < (2'h3)); forvar1205 = (forvar1205 + (1'h1)))
            begin
              reg1206 = (|$signed((!reg1068)));
              reg1207 <= {($signed(reg1084[(5'h16):(4'he)]) | reg1164)};
              reg1208 = $unsigned(reg1164);
              reg1209 = reg1101[(1'h0):(1'h0)];
            end
          reg1210 <= $signed($unsigned((-$unsigned((reg1118 ?
              reg1154 : reg1099)))));
          reg1211 = wire902;
        end
    end
  assign wire1212 = (~&(&reg1153[(3'h4):(2'h2)]));
  assign wire1213 = reg1181;
  always
    @(posedge clk) begin
      reg1214 <= reg1112[(4'hc):(2'h2)];
      reg1215 = ((($signed((wire900 ?
          reg1156 : reg1068)) - (^~reg1086)) || $unsigned((^$signed(reg1207)))) || ((~(reg1086 << (wire1213 & reg1164))) ?
          $signed($signed((reg1086 ^ reg1107))) : $unsigned($signed({reg1107}))));
      reg1216 = reg1156;
      if ((-reg1174))
        begin
          reg1217 <= (^({(reg1133 ? (+wire1087) : (reg1084 != reg1128)),
              (reg1190[(3'h6):(2'h3)] != (reg1158 << reg1076))} & $signed($unsigned(reg1135[(4'he):(4'h9)]))));
          if (($unsigned({wire902[(2'h2):(1'h1)]}) ?
              (8'hb9) : ({$signed((~^(8'haa))),
                      ((reg1123 ?
                          reg1118 : (8'ha2)) * reg1179[(5'h12):(4'h9)])} ?
                  $signed((!reg1091)) : $unsigned({(8'hbe), reg1101}))))
            begin
              reg1218 <= {(reg1153[(2'h2):(1'h0)] * $unsigned({$signed((7'h45))}))};
              reg1219 = wire1089[(2'h2):(1'h1)];
              reg1220 = reg1099[(2'h3):(1'h0)];
            end
          else
            begin
              reg1219 = reg1156[(3'h5):(3'h5)];
              reg1221 <= ((reg1123[(1'h1):(1'h1)] >> ($unsigned((~wire902)) ?
                  ((&reg1099) ?
                      (reg1128 != wire902) : (reg1175 < reg1084)) : ((reg1084 ?
                          reg1215 : wire900) ?
                      (~|reg1174) : (~reg1134)))) < $signed(reg1091[(3'h7):(1'h1)]));
              reg1222 <= (8'hb0);
            end
        end
      else
        begin
          reg1217 <= $unsigned({{($unsigned((8'h9e)) >> reg1175[(3'h4):(2'h3)])},
              (reg1129 ~^ (~^(reg1168 >= reg1178)))});
          reg1219 = reg1217[(3'h7):(3'h7)];
          for (forvar1220 = (1'h0); (forvar1220 < (1'h1)); forvar1220 = (forvar1220 + (1'h1)))
            begin
              reg1221 <= ($signed($unsigned(($signed(reg1195) <= $unsigned(reg1159)))) >> reg1123[(2'h2):(1'h0)]);
              reg1222 <= wire1089;
              reg1223 <= reg1123;
              reg1224 = (reg1076 ?
                  reg1113 : $unsigned((~|($unsigned((8'hb2)) * $unsigned(wire1087)))));
              reg1225 <= (8'haf);
            end
        end
    end
  assign wire1226 = (~&(reg1168 >> (~($unsigned(reg1106) ?
                        reg1179 : (reg1168 | reg1185)))));
  module1227 #() modinst1454 (wire1453, clk, reg1167, reg1113, wire1069, reg1189, reg1143);
  always
    @(posedge clk) begin
      for (forvar1455 = (1'h0); (forvar1455 < (1'h0)); forvar1455 = (forvar1455 + (1'h1)))
        begin
          for (forvar1456 = (1'h0); (forvar1456 < (1'h1)); forvar1456 = (forvar1456 + (1'h1)))
            begin
              reg1457 = {(~&(^~$unsigned($signed(reg1159)))), reg1183};
              reg1458 <= $unsigned(($unsigned($signed($signed(reg1091))) ?
                  ({(7'h46)} ?
                      {(~reg1133)} : (~&$unsigned(wire897))) : reg1196));
              reg1459 = $signed($unsigned($signed(wire899)));
            end
          reg1460 = reg1196;
          reg1461 = $unsigned(reg1210[(1'h0):(1'h0)]);
          if (reg1085[(4'ha):(2'h2)])
            begin
              reg1462 <= (8'h9d);
              reg1463 = {$signed((((reg1123 != (8'h9e)) <<< (reg1129 ?
                          forvar1455 : (7'h44))) ?
                      (&(reg1135 ?
                          reg1167 : reg1190)) : (wire1089 + reg1181[(2'h2):(1'h0)]))),
                  ((~&$signed(reg1122[(4'ha):(3'h6)])) ?
                      wire897 : reg1180[(5'h10):(4'hc)])};
              reg1464 <= (reg1460[(4'ha):(2'h3)] ?
                  {$unsigned($signed(reg1217))} : ((reg1463 > reg1203[(1'h1):(1'h0)]) ?
                      (reg1076 ?
                          reg1192[(5'h14):(3'h7)] : (reg1457 == (&(8'ha9)))) : $signed($unsigned((^reg1190)))));
            end
          else
            begin
              reg1462 <= (^((($unsigned(wire1087) | (forvar1456 ?
                      reg1196 : reg1086)) + ($unsigned((8'hbe)) ?
                      $unsigned(reg1135) : {reg1118, reg1214})) ?
                  $signed($unsigned(wire1066)) : (($unsigned(reg1129) ?
                          (reg1159 || (8'ha2)) : reg1196[(3'h6):(2'h2)]) ?
                      {wire897, wire1212[(3'h6):(1'h1)]} : reg1168)));
              reg1464 <= (~|(!reg1183[(1'h1):(1'h1)]));
              reg1465 = $unsigned(wire902);
              reg1466 = ((^(((wire1069 ~^ (8'hac)) >> (^reg1134)) <<< reg1180[(4'h9):(4'h8)])) ?
                  ($unsigned($signed(reg1460)) ~^ ($signed($unsigned(wire1226)) ?
                      reg1161 : $signed($unsigned(reg1459)))) : {(wire899[(3'h7):(3'h4)] ?
                          $unsigned((reg1128 ~^ reg1113)) : (((8'hab) != reg1217) ?
                              $unsigned(wire897) : $signed(reg1156))),
                      ((~&(reg1143 ?
                          reg1106 : reg1072)) ^ $unsigned(reg1083))});
              reg1467 <= (~reg1117);
            end
          for (forvar1468 = (1'h0); (forvar1468 < (1'h1)); forvar1468 = (forvar1468 + (1'h1)))
            begin
              reg1469 = ({(8'haa)} ?
                  (reg1186[(3'h6):(3'h5)] != reg1112) : (($signed((reg1458 - reg1093)) ?
                          (reg1159 ?
                              (reg1467 ? reg1467 : reg1198) : (reg1068 ?
                                  reg1180 : reg1183)) : $unsigned($signed(reg1115))) ?
                      reg1107 : (!($unsigned((7'h45)) ?
                          reg1068[(3'h6):(2'h2)] : (reg1091 << reg1164)))));
            end
        end
      reg1470 <= ((~&(wire902 < (reg1225 ?
          reg1464[(2'h3):(2'h3)] : (~wire1087)))) ^ (~(!({reg1196, wire1212} ?
          reg1134[(4'hc):(4'h8)] : {reg1134, reg1076}))));
      if ($unsigned(wire1213[(4'ha):(4'h9)]))
        begin
          if ((reg1222 + $unsigned(reg1225)))
            begin
              reg1471 <= reg1134[(5'h10):(3'h4)];
              reg1472 <= $unsigned(reg1104[(3'h6):(3'h4)]);
            end
          else
            begin
              reg1473 = $signed($signed(((reg1179[(3'h5):(1'h1)] >> (forvar1468 ~^ reg1084)) ?
                  $unsigned({reg1207, reg1465}) : {$signed(reg1179)})));
              reg1474 <= (~&$signed((^~(((7'h43) && reg1167) * (8'ha6)))));
              reg1475 = $unsigned((reg1192[(4'h9):(3'h7)] ?
                  (reg1470 | {(-forvar1468)}) : ($signed($signed((8'hbe))) * $signed(reg1099[(4'hd):(4'hd)]))));
              reg1476 <= (!reg1137);
              reg1477 <= ($unsigned(($unsigned((~&reg1467)) >= ((reg1473 ?
                  (8'hbb) : reg1122) | (&reg1210)))) << ((((reg1466 & reg1113) ?
                      $unsigned(reg1203) : reg1174[(5'h10):(4'hd)]) ?
                  $signed({reg1466}) : ((reg1203 << forvar1455) ?
                      forvar1456[(3'h4):(1'h1)] : reg1117[(5'h11):(4'he)])) <= ({wire897[(1'h0):(1'h0)]} ?
                  $unsigned(reg1153[(3'h4):(1'h1)]) : $signed((|reg1161)))));
            end
          reg1478 <= $signed($signed((!reg1159)));
          reg1479 = $signed($signed(wire902[(3'h5):(3'h5)]));
        end
      else
        begin
          reg1471 <= reg1175;
          reg1473 = (reg1223 ?
              reg1135 : ($signed(reg1115[(4'ha):(2'h2)]) ?
                  (+$unsigned((reg1112 ^ wire1089))) : (((reg1164 + reg1159) && (^forvar1468)) & (8'hb5))));
          reg1475 = reg1199[(3'h6):(3'h5)];
        end
      reg1480 <= reg1134[(3'h6):(2'h3)];
      for (forvar1481 = (1'h0); (forvar1481 < (3'h4)); forvar1481 = (forvar1481 + (1'h1)))
        begin
          reg1482 = forvar1456;
          if (reg1092)
            begin
              reg1483 = ((-(reg1465 || (|(!reg1474)))) ?
                  {reg1135, reg1183} : (|reg1218));
            end
          else
            begin
              reg1483 = $unsigned(reg1128[(3'h7):(3'h7)]);
              reg1484 = ($unsigned((^~reg1472)) ?
                  ({({reg1469} ? (+reg1178) : {reg1192, reg1092}),
                      reg1190} << (reg1092 ?
                      $signed($signed(reg1480)) : (-(reg1473 - reg1092)))) : {(~^reg1477[(4'h9):(1'h1)]),
                      reg1104[(4'he):(4'hd)]});
              reg1485 = (|($signed({$unsigned(reg1153),
                  (reg1469 ? forvar1455 : reg1091)}) ^ (8'hbd)));
            end
          if ((reg1460[(4'ha):(3'h7)] ?
              ((-$unsigned(((7'h49) == reg1129))) ?
                  reg1458[(2'h3):(1'h1)] : forvar1456) : {reg1458}))
            begin
              reg1486 <= (($unsigned((reg1479[(3'h6):(3'h5)] ?
                  reg1460[(4'hf):(1'h1)] : $signed(reg1113))) >= ($unsigned((reg1217 * reg1133)) ?
                  reg1098 : {$signed(reg1464),
                      (reg1095 ?
                          reg1112 : reg1068)})) * reg1099[(1'h1):(1'h1)]);
              reg1487 <= ((((|{reg1217}) ?
                      wire899 : reg1192[(2'h3):(1'h1)]) <= (~^((reg1474 != (8'ha1)) ?
                      $signed((7'h48)) : reg1186[(4'h9):(4'h9)]))) ?
                  (reg1106[(3'h4):(1'h0)] < {(|(reg1135 ? reg1135 : reg1156)),
                      $unsigned((reg1474 <= reg1158))}) : $unsigned({$signed((wire898 == wire900)),
                      forvar1468[(2'h2):(2'h2)]}));
              reg1488 = ((^wire1066) ?
                  ((((reg1464 && reg1185) >= (~|reg1198)) | (^~(^reg1107))) ^~ {reg1178[(5'h10):(5'h10)]}) : reg1190[(3'h5):(2'h2)]);
            end
          else
            begin
              reg1488 = $signed($signed(($unsigned(reg1084) ~^ reg1483)));
              reg1489 <= ((~^(($unsigned((7'h45)) ?
                          reg1103[(4'h8):(4'h8)] : (~&(7'h49))) ?
                      reg1128[(2'h3):(1'h1)] : $signed(reg1180))) ?
                  reg1175[(2'h3):(1'h1)] : (-(!(7'h40))));
              reg1490 <= (~|((($unsigned(reg1461) + (reg1178 - reg1172)) & ($unsigned(reg1207) >>> reg1104[(4'hd):(3'h4)])) <= {$unsigned($unsigned((8'hb3))),
                  ((reg1178 <= wire1087) ?
                      (reg1187 >>> reg1207) : $unsigned((8'ha8)))}));
            end
          reg1491 = $unsigned((8'hb4));
        end
    end
  assign wire1492 = reg1153;
  always
    @(posedge clk) begin
      reg1493 = {$signed(({$unsigned((8'haa))} >= (reg1091 | reg1476[(3'h5):(3'h5)])))};
    end
  assign wire1494 = ($unsigned({wire902}) * $unsigned($unsigned($unsigned(reg1072))));
  always
    @(posedge clk) begin
      for (forvar1495 = (1'h0); (forvar1495 < (3'h4)); forvar1495 = (forvar1495 + (1'h1)))
        begin
          if ((|reg1217[(3'h6):(3'h5)]))
            begin
              reg1496 <= reg1198[(1'h1):(1'h0)];
              reg1497 = (($unsigned((reg1118[(4'hc):(2'h3)] + {reg1153})) ?
                      ($signed($signed(reg1106)) ?
                          (^~$signed(reg1093)) : ($signed(reg1156) & $unsigned(reg1478))) : reg1159) ?
                  reg1134 : ($unsigned((8'hb8)) ? reg1496 : {reg1112}));
              reg1498 = (($unsigned({(wire900 ? wire1069 : reg1072),
                      (reg1085 ? reg1128 : wire1087)}) ?
                  (~&(reg1138[(4'hf):(2'h3)] != reg1159[(3'h7):(3'h4)])) : (wire1069[(3'h6):(1'h1)] | reg1476)) & $signed($unsigned($signed(wire1226))));
              reg1499 <= reg1467;
              reg1500 = reg1190;
            end
          else
            begin
              reg1497 = $unsigned(reg1085);
              reg1498 = reg1497[(1'h0):(1'h0)];
            end
        end
      if (reg1085[(3'h6):(3'h4)])
        begin
          if ((!$unsigned((^~reg1137[(1'h0):(1'h0)]))))
            begin
              reg1501 <= (|wire1212[(2'h2):(1'h1)]);
              reg1502 <= forvar1495;
              reg1503 <= $unsigned(reg1174[(4'ha):(4'h8)]);
            end
          else
            begin
              reg1504 = $unsigned((8'haa));
              reg1505 = (-reg1135);
              reg1506 <= reg1092[(1'h0):(1'h0)];
              reg1507 = reg1185;
            end
          reg1508 <= $signed(reg1472);
          reg1509 = $signed(($unsigned(((^wire900) ?
              (|reg1210) : reg1467)) + (wire900[(5'h10):(2'h3)] ?
              {reg1168} : reg1106)));
          reg1510 = {reg1506,
              {$signed(($unsigned(reg1143) ?
                      (reg1161 ? reg1499 : (8'ha5)) : $signed(reg1128))),
                  reg1503[(4'h8):(1'h1)]}};
        end
      else
        begin
          reg1501 <= reg1185[(3'h6):(1'h0)];
        end
      if (reg1498)
        begin
          for (forvar1511 = (1'h0); (forvar1511 < (1'h1)); forvar1511 = (forvar1511 + (1'h1)))
            begin
              reg1512 <= reg1198;
              reg1513 <= $signed({(((~&reg1158) | $signed((7'h47))) & ($unsigned((8'hb4)) & (7'h46)))});
              reg1514 = ((+($signed((reg1098 ? (8'hb9) : reg1478)) ?
                      ($unsigned((8'hac)) ^~ reg1084[(4'ha):(3'h5)]) : {(|reg1207),
                          (reg1084 ^~ reg1159)})) ?
                  $signed($signed($unsigned($signed(reg1085)))) : reg1138[(5'h14):(3'h5)]);
              reg1515 <= reg1221;
              reg1516 <= wire897;
            end
        end
      else
        begin
          if ($unsigned(($unsigned(reg1106) - $signed((!$unsigned(reg1472))))))
            begin
              reg1511 <= (&$signed($signed($signed((-reg1501)))));
              reg1514 = ((~&$unsigned((reg1158[(2'h2):(2'h2)] ~^ $unsigned(reg1196)))) ?
                  wire900[(1'h1):(1'h0)] : $unsigned((&(reg1128[(1'h1):(1'h0)] ?
                      reg1474 : $unsigned((7'h4a))))));
              reg1515 <= {reg1476[(2'h3):(1'h1)],
                  {((reg1076 ? reg1214 : (7'h41)) ?
                          ((|reg1210) ?
                              reg1172 : (reg1158 ?
                                  reg1496 : reg1512)) : {(reg1505 << wire899)}),
                      (^~reg1091[(4'hf):(1'h1)])}};
              reg1516 <= $signed($signed((~reg1503[(1'h0):(1'h0)])));
              reg1517 <= reg1504[(2'h3):(1'h0)];
            end
          else
            begin
              reg1514 = $signed($signed(($unsigned((reg1190 ?
                      reg1203 : reg1517)) ?
                  $unsigned((wire1492 >= reg1174)) : wire1213)));
              reg1515 <= (({wire1492} ~^ ((!reg1195) ^ reg1129[(3'h6):(1'h0)])) ?
                  (8'haa) : reg1129[(1'h0):(1'h0)]);
              reg1518 = reg1112[(3'h7):(2'h3)];
            end
          if ((-$signed(reg1192)))
            begin
              reg1519 <= $unsigned(($unsigned($signed($signed(reg1486))) ?
                  (~^reg1092[(2'h3):(1'h0)]) : reg1092[(1'h1):(1'h0)]));
              reg1520 <= ($unsigned($unsigned(reg1187)) * reg1156);
            end
          else
            begin
              reg1521 = reg1181[(4'hf):(3'h5)];
            end
          reg1522 <= (^~$unsigned((reg1113[(3'h6):(3'h4)] ?
              wire1069[(5'h16):(3'h5)] : $unsigned($signed(reg1118)))));
        end
      if ((^(~|((reg1198[(1'h0):(1'h0)] ?
          (reg1508 ^ reg1478) : reg1504) | reg1175))))
        begin
          reg1523 <= reg1174[(5'h14):(2'h2)];
          reg1524 <= reg1093;
        end
      else
        begin
          reg1525 = $unsigned(($signed($unsigned(reg1474)) ?
              ({$signed(reg1198)} ?
                  (7'h4a) : {(reg1478 ?
                          reg1500 : reg1156)}) : {$signed($unsigned(reg1223))}));
        end
    end
  assign wire1526 = $unsigned((reg1107[(3'h4):(1'h1)] == (($unsigned(reg1499) ?
                            $unsigned(wire1088) : ((8'ha9) == (7'h45))) ?
                        (((8'hb9) >= reg1158) ?
                            (reg1519 && (7'h49)) : $signed(reg1129)) : (~reg1181))));
  module1527 #() modinst1618 (wire1617, clk, reg1104, reg1476, reg1099, reg1143);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module103
#(parameter param798 = (~^(^~((((8'ha4) & (8'hb2)) ? ((8'hb1) >>> (8'ha0)) : (-(8'hbf))) ? ((-(8'ha6)) ? ((8'ha3) < (8'ha3)) : ((7'h41) >>> (8'ha6))) : ((^~(8'hbf)) ? {(8'hb9), (7'h44)} : (8'haa))))), 
parameter param799 = (param798 << ((8'hb7) ? param798 : (^~{(param798 ? param798 : param798), (+param798)}))))
(y, clk, wire107, wire106, wire105, wire104);
  output wire [(32'hdc2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire107;
  input wire [(4'hf):(1'h0)] wire106;
  input wire signed [(4'hb):(1'h0)] wire105;
  input wire signed [(5'h13):(1'h0)] wire104;
  wire signed [(5'h18):(1'h0)] wire764;
  wire signed [(3'h6):(1'h0)] wire642;
  wire [(3'h6):(1'h0)] wire496;
  wire signed [(5'h14):(1'h0)] wire480;
  wire [(2'h2):(1'h0)] wire479;
  wire [(5'h13):(1'h0)] wire422;
  reg [(4'hf):(1'h0)] reg797 = (1'h0);
  reg [(3'h6):(1'h0)] reg796 = (1'h0);
  reg [(5'h12):(1'h0)] reg795 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg792 = (1'h0);
  reg [(4'hc):(1'h0)] reg791 = (1'h0);
  reg [(5'h12):(1'h0)] reg788 = (1'h0);
  reg [(4'ha):(1'h0)] reg786 = (1'h0);
  reg signed [(4'he):(1'h0)] reg785 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg784 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg783 = (1'h0);
  reg [(4'h8):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg779 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg776 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg775 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg774 = (1'h0);
  reg [(5'h12):(1'h0)] reg763 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg761 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg760 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg758 = (1'h0);
  reg [(3'h4):(1'h0)] reg755 = (1'h0);
  reg [(2'h3):(1'h0)] reg753 = (1'h0);
  reg signed [(4'he):(1'h0)] reg752 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg748 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg745 = (1'h0);
  reg [(3'h4):(1'h0)] reg740 = (1'h0);
  reg [(5'h18):(1'h0)] reg732 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg731 = (1'h0);
  reg [(4'hd):(1'h0)] reg730 = (1'h0);
  reg [(3'h7):(1'h0)] reg728 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg724 = (1'h0);
  reg [(5'h15):(1'h0)] reg721 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg718 = (1'h0);
  reg [(4'h9):(1'h0)] reg717 = (1'h0);
  reg [(5'h13):(1'h0)] reg711 = (1'h0);
  reg [(4'hb):(1'h0)] reg707 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg706 = (1'h0);
  reg [(4'hc):(1'h0)] reg698 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg694 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg693 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg689 = (1'h0);
  reg [(5'h16):(1'h0)] reg688 = (1'h0);
  reg [(4'he):(1'h0)] reg685 = (1'h0);
  reg [(5'h10):(1'h0)] reg683 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg682 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg681 = (1'h0);
  reg [(2'h3):(1'h0)] reg679 = (1'h0);
  reg [(3'h4):(1'h0)] reg677 = (1'h0);
  reg [(4'h8):(1'h0)] reg674 = (1'h0);
  reg [(3'h7):(1'h0)] reg672 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg666 = (1'h0);
  reg [(4'h9):(1'h0)] reg665 = (1'h0);
  reg signed [(4'he):(1'h0)] reg660 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg654 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg653 = (1'h0);
  reg [(4'hd):(1'h0)] reg645 = (1'h0);
  reg [(5'h16):(1'h0)] reg534 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg531 = (1'h0);
  reg [(5'h13):(1'h0)] reg530 = (1'h0);
  reg [(5'h13):(1'h0)] reg528 = (1'h0);
  reg [(4'hf):(1'h0)] reg523 = (1'h0);
  reg [(4'hb):(1'h0)] reg522 = (1'h0);
  reg [(4'h8):(1'h0)] reg521 = (1'h0);
  reg [(3'h5):(1'h0)] reg520 = (1'h0);
  reg [(3'h5):(1'h0)] reg506 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg512 = (1'h0);
  reg [(5'h14):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg505 = (1'h0);
  reg [(5'h16):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg500 = (1'h0);
  reg [(4'h9):(1'h0)] reg493 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg492 = (1'h0);
  reg [(5'h13):(1'h0)] reg490 = (1'h0);
  reg [(5'h11):(1'h0)] reg489 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg487 = (1'h0);
  reg [(4'ha):(1'h0)] reg486 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg485 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg484 = (1'h0);
  reg [(5'h16):(1'h0)] reg483 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg477 = (1'h0);
  reg [(4'h9):(1'h0)] reg475 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg472 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg466 = (1'h0);
  reg [(4'h8):(1'h0)] reg462 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg461 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg458 = (1'h0);
  reg [(5'h14):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg453 = (1'h0);
  reg [(5'h18):(1'h0)] reg452 = (1'h0);
  reg [(5'h16):(1'h0)] reg451 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg450 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg447 = (1'h0);
  reg [(4'ha):(1'h0)] reg445 = (1'h0);
  reg [(5'h18):(1'h0)] reg444 = (1'h0);
  reg [(4'h9):(1'h0)] reg438 = (1'h0);
  reg [(5'h17):(1'h0)] reg424 = (1'h0);
  reg [(4'hc):(1'h0)] reg427 = (1'h0);
  reg [(3'h5):(1'h0)] reg794 = (1'h0);
  reg [(5'h18):(1'h0)] reg793 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg790 = (1'h0);
  reg [(5'h11):(1'h0)] reg789 = (1'h0);
  reg [(4'h9):(1'h0)] reg787 = (1'h0);
  reg [(3'h7):(1'h0)] reg782 = (1'h0);
  reg [(3'h4):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg778 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar777 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar773 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar772 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg771 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg770 = (1'h0);
  reg [(5'h16):(1'h0)] forvar769 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar768 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg767 = (1'h0);
  reg [(4'hb):(1'h0)] reg766 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar765 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg762 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar757 = (1'h0);
  reg [(4'h9):(1'h0)] reg756 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg754 = (1'h0);
  reg [(3'h5):(1'h0)] reg751 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg750 = (1'h0);
  reg [(5'h12):(1'h0)] forvar749 = (1'h0);
  reg [(4'hf):(1'h0)] reg741 = (1'h0);
  reg [(4'h8):(1'h0)] reg747 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg746 = (1'h0);
  reg [(4'h9):(1'h0)] forvar744 = (1'h0);
  reg [(5'h15):(1'h0)] reg743 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg742 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar741 = (1'h0);
  reg [(3'h7):(1'h0)] reg739 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg738 = (1'h0);
  reg [(5'h10):(1'h0)] reg737 = (1'h0);
  reg [(3'h7):(1'h0)] reg736 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar735 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg734 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg733 = (1'h0);
  reg [(5'h14):(1'h0)] reg729 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg727 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg726 = (1'h0);
  reg [(3'h4):(1'h0)] reg725 = (1'h0);
  reg [(4'ha):(1'h0)] reg723 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg722 = (1'h0);
  reg [(3'h4):(1'h0)] forvar720 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg719 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg716 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar714 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar713 = (1'h0);
  reg [(4'he):(1'h0)] reg712 = (1'h0);
  reg [(2'h2):(1'h0)] reg710 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg709 = (1'h0);
  reg [(5'h18):(1'h0)] reg708 = (1'h0);
  reg [(4'h9):(1'h0)] forvar705 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg704 = (1'h0);
  reg [(4'he):(1'h0)] reg703 = (1'h0);
  reg [(5'h12):(1'h0)] forvar702 = (1'h0);
  reg [(5'h12):(1'h0)] reg701 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg700 = (1'h0);
  reg signed [(4'he):(1'h0)] reg699 = (1'h0);
  reg [(4'h8):(1'h0)] reg697 = (1'h0);
  reg [(3'h5):(1'h0)] reg696 = (1'h0);
  reg [(2'h2):(1'h0)] forvar695 = (1'h0);
  reg [(5'h11):(1'h0)] forvar692 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg692 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg691 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg690 = (1'h0);
  reg [(3'h4):(1'h0)] reg687 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg686 = (1'h0);
  reg [(5'h13):(1'h0)] reg684 = (1'h0);
  reg [(3'h4):(1'h0)] forvar680 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg678 = (1'h0);
  reg [(4'h9):(1'h0)] forvar672 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg676 = (1'h0);
  reg [(3'h5):(1'h0)] reg675 = (1'h0);
  reg [(3'h4):(1'h0)] reg673 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg671 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg669 = (1'h0);
  reg [(3'h6):(1'h0)] reg668 = (1'h0);
  reg [(4'ha):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg663 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar662 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg661 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar659 = (1'h0);
  reg [(5'h18):(1'h0)] reg658 = (1'h0);
  reg [(5'h14):(1'h0)] reg657 = (1'h0);
  reg [(3'h4):(1'h0)] reg656 = (1'h0);
  reg [(4'hd):(1'h0)] reg655 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg652 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg651 = (1'h0);
  reg [(3'h5):(1'h0)] reg650 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar649 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg648 = (1'h0);
  reg [(4'hf):(1'h0)] reg647 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg646 = (1'h0);
  reg [(5'h18):(1'h0)] reg644 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg533 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg532 = (1'h0);
  reg [(3'h5):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar527 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg526 = (1'h0);
  reg [(4'hf):(1'h0)] reg525 = (1'h0);
  reg [(2'h3):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg519 = (1'h0);
  reg [(2'h3):(1'h0)] forvar518 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg517 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg516 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar515 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar505 = (1'h0);
  reg [(2'h3):(1'h0)] reg514 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg511 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg509 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg508 = (1'h0);
  reg signed [(4'he):(1'h0)] reg507 = (1'h0);
  reg [(5'h12):(1'h0)] forvar506 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg503 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar502 = (1'h0);
  reg [(4'h8):(1'h0)] reg501 = (1'h0);
  reg signed [(4'he):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg498 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar497 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg497 = (1'h0);
  reg [(4'hb):(1'h0)] reg495 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg494 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg491 = (1'h0);
  reg [(3'h5):(1'h0)] reg488 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar482 = (1'h0);
  reg [(5'h14):(1'h0)] forvar481 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg476 = (1'h0);
  reg [(3'h5):(1'h0)] reg474 = (1'h0);
  reg [(3'h4):(1'h0)] forvar473 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg471 = (1'h0);
  reg [(3'h6):(1'h0)] reg470 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar469 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar468 = (1'h0);
  reg [(5'h12):(1'h0)] reg467 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg465 = (1'h0);
  reg [(5'h13):(1'h0)] forvar464 = (1'h0);
  reg [(4'ha):(1'h0)] reg463 = (1'h0);
  reg [(5'h17):(1'h0)] forvar459 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg455 = (1'h0);
  reg [(4'hc):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg460 = (1'h0);
  reg [(4'h8):(1'h0)] reg459 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg457 = (1'h0);
  reg [(3'h7):(1'h0)] forvar455 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg449 = (1'h0);
  reg [(4'he):(1'h0)] forvar448 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg446 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg443 = (1'h0);
  reg [(5'h15):(1'h0)] reg442 = (1'h0);
  reg [(5'h10):(1'h0)] forvar441 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg440 = (1'h0);
  reg [(5'h11):(1'h0)] reg439 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg436 = (1'h0);
  reg [(5'h11):(1'h0)] reg435 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar434 = (1'h0);
  reg [(2'h2):(1'h0)] forvar433 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg432 = (1'h0);
  reg [(4'ha):(1'h0)] reg431 = (1'h0);
  reg [(4'hd):(1'h0)] reg430 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg429 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar425 = (1'h0);
  reg [(5'h14):(1'h0)] reg426 = (1'h0);
  reg [(2'h3):(1'h0)] reg425 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar424 = (1'h0);
  assign y = {wire764,
                 wire642,
                 wire496,
                 wire480,
                 wire479,
                 wire422,
                 reg797,
                 reg796,
                 reg795,
                 reg792,
                 reg791,
                 reg788,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 reg781,
                 reg779,
                 reg776,
                 reg775,
                 reg774,
                 reg763,
                 reg761,
                 reg760,
                 reg758,
                 reg755,
                 reg753,
                 reg752,
                 reg748,
                 reg745,
                 reg740,
                 reg732,
                 reg731,
                 reg730,
                 reg728,
                 reg724,
                 reg721,
                 reg718,
                 reg717,
                 reg711,
                 reg707,
                 reg706,
                 reg698,
                 reg694,
                 reg693,
                 reg689,
                 reg688,
                 reg685,
                 reg683,
                 reg682,
                 reg681,
                 reg679,
                 reg677,
                 reg674,
                 reg672,
                 reg667,
                 reg666,
                 reg665,
                 reg660,
                 reg654,
                 reg653,
                 reg645,
                 reg534,
                 reg531,
                 reg530,
                 reg528,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 reg506,
                 reg513,
                 reg512,
                 reg510,
                 reg505,
                 reg504,
                 reg500,
                 reg493,
                 reg492,
                 reg490,
                 reg489,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg478,
                 reg477,
                 reg475,
                 reg472,
                 reg466,
                 reg462,
                 reg461,
                 reg458,
                 reg456,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg447,
                 reg445,
                 reg444,
                 reg438,
                 reg424,
                 reg427,
                 reg794,
                 reg793,
                 reg790,
                 reg789,
                 reg787,
                 reg782,
                 reg780,
                 reg778,
                 forvar777,
                 forvar773,
                 forvar772,
                 reg771,
                 reg770,
                 forvar769,
                 forvar768,
                 reg767,
                 reg766,
                 forvar765,
                 reg762,
                 reg759,
                 forvar757,
                 reg756,
                 reg754,
                 reg751,
                 reg750,
                 forvar749,
                 reg741,
                 reg747,
                 reg746,
                 forvar744,
                 reg743,
                 reg742,
                 forvar741,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 forvar735,
                 reg734,
                 reg733,
                 reg729,
                 reg727,
                 reg726,
                 reg725,
                 reg723,
                 reg722,
                 forvar720,
                 reg719,
                 reg716,
                 reg715,
                 forvar714,
                 forvar713,
                 reg712,
                 reg710,
                 reg709,
                 reg708,
                 forvar705,
                 reg704,
                 reg703,
                 forvar702,
                 reg701,
                 reg700,
                 reg699,
                 reg697,
                 reg696,
                 forvar695,
                 forvar692,
                 reg692,
                 reg691,
                 reg690,
                 reg687,
                 reg686,
                 reg684,
                 forvar680,
                 reg678,
                 forvar672,
                 reg676,
                 reg675,
                 reg673,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 reg664,
                 reg663,
                 forvar662,
                 reg661,
                 forvar659,
                 reg658,
                 reg657,
                 reg656,
                 reg655,
                 reg652,
                 reg651,
                 reg650,
                 forvar649,
                 reg648,
                 reg647,
                 reg646,
                 reg644,
                 reg535,
                 reg533,
                 reg532,
                 reg529,
                 forvar527,
                 reg526,
                 reg525,
                 reg524,
                 reg519,
                 forvar518,
                 reg517,
                 reg516,
                 forvar515,
                 forvar505,
                 reg514,
                 reg511,
                 reg509,
                 reg508,
                 reg507,
                 forvar506,
                 reg503,
                 forvar502,
                 reg501,
                 reg499,
                 reg498,
                 forvar497,
                 reg497,
                 reg495,
                 reg494,
                 reg491,
                 reg488,
                 forvar482,
                 forvar481,
                 reg476,
                 reg474,
                 forvar473,
                 reg471,
                 reg470,
                 forvar469,
                 forvar468,
                 reg467,
                 reg465,
                 forvar464,
                 reg463,
                 forvar459,
                 reg455,
                 reg448,
                 reg460,
                 reg459,
                 reg457,
                 forvar455,
                 reg449,
                 forvar448,
                 reg446,
                 reg443,
                 reg442,
                 forvar441,
                 reg440,
                 reg439,
                 reg437,
                 reg436,
                 reg435,
                 forvar434,
                 forvar433,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 forvar425,
                 reg426,
                 reg425,
                 forvar424,
                 (1'h0)};
  module108 #() modinst423 (wire422, clk, wire106, wire107, wire104, wire105, (8'h9e));
  always
    @(posedge clk) begin
      if ($signed($signed($signed(($unsigned((8'hb2)) * (wire422 ?
          wire105 : wire422))))))
        begin
          for (forvar424 = (1'h0); (forvar424 < (2'h2)); forvar424 = (forvar424 + (1'h1)))
            begin
              reg425 = wire104;
            end
          reg426 = ($signed(reg425[(1'h1):(1'h1)]) < {wire104[(5'h11):(3'h4)],
              $unsigned((7'h47))});
          reg427 <= (~(8'ha0));
        end
      else
        begin
          reg424 <= ((forvar424 * wire104) != (~&$unsigned((^reg427[(4'h9):(1'h1)]))));
          for (forvar425 = (1'h0); (forvar425 < (2'h3)); forvar425 = (forvar425 + (1'h1)))
            begin
              reg427 <= $unsigned((7'h45));
              reg428 = $signed($unsigned($unsigned(forvar424)));
              reg429 = {($unsigned($signed($signed(wire104))) | $signed({(wire104 ?
                          (8'hbc) : reg428),
                      wire105})),
                  (reg425 ^~ ((~^reg426) >>> (reg425 ?
                      (+reg424) : (!wire104))))};
              reg430 = ($unsigned($unsigned(($signed(forvar424) <<< $signed(reg425)))) < forvar425[(3'h7):(3'h5)]);
              reg431 = $unsigned($signed($unsigned(wire107)));
            end
        end
      reg432 = (~|reg424[(4'hd):(1'h0)]);
    end
  always
    @(posedge clk) begin
      for (forvar433 = (1'h0); (forvar433 < (1'h1)); forvar433 = (forvar433 + (1'h1)))
        begin
          for (forvar434 = (1'h0); (forvar434 < (3'h4)); forvar434 = (forvar434 + (1'h1)))
            begin
              reg435 = (+wire106[(4'h9):(3'h5)]);
            end
          if ($signed(({wire105, wire104[(4'hb):(3'h6)]} ?
              wire104[(5'h13):(3'h6)] : (~$signed({wire107})))))
            begin
              reg436 = ((-$unsigned((-(reg427 >= (8'hbf))))) ?
                  $signed(reg435) : (-{$unsigned((wire107 ?
                          forvar433 : reg424))}));
            end
          else
            begin
              reg436 = (reg427 ?
                  ($unsigned(((7'h44) > $unsigned((8'hb6)))) ?
                      reg427 : wire104[(3'h6):(2'h3)]) : $signed(($signed((wire104 ?
                      reg435 : reg435)) ~^ {$signed(wire422),
                      forvar433[(1'h1):(1'h0)]})));
              reg437 = wire107;
              reg438 <= (reg424 ^~ $unsigned((8'ha5)));
            end
          reg439 = ((+(~&reg438)) ?
              $unsigned($unsigned(((forvar434 ^ wire106) ?
                  (wire106 + reg427) : {wire105,
                      wire106}))) : (~|wire106[(2'h3):(1'h1)]));
          reg440 = $signed((({(forvar434 ?
                      reg437 : wire107)} ^ {reg439[(3'h5):(3'h4)]}) ?
              ($signed((forvar434 ? (7'h43) : wire105)) | ($unsigned(wire422) ?
                  forvar433 : reg439)) : ((&{reg435, reg424}) ?
                  wire105[(1'h1):(1'h1)] : $signed((wire107 && wire107)))));
        end
      for (forvar441 = (1'h0); (forvar441 < (1'h0)); forvar441 = (forvar441 + (1'h1)))
        begin
          if ($signed(reg435))
            begin
              reg442 = $signed(reg437[(3'h6):(2'h3)]);
              reg443 = {(reg439 ?
                      $unsigned(wire422) : ($signed((forvar441 | (7'h45))) ?
                          ({wire105} ?
                              reg439[(4'hd):(4'h8)] : (^forvar441)) : ($signed(reg440) && $unsigned(forvar433)))),
                  ($signed(reg438) ?
                      ({(wire104 >> (8'hbe))} <<< (~^$unsigned(forvar433))) : (((|(8'hac)) ?
                          $unsigned(reg436) : (8'ha9)) * reg442[(4'hf):(4'hd)]))};
            end
          else
            begin
              reg444 <= ((8'h9d) ? $unsigned((-(8'had))) : $signed(forvar441));
              reg445 <= {$unsigned(($unsigned($unsigned(reg440)) >= {$unsigned(reg437),
                      $signed(wire422)})),
                  (reg443 >> (wire106 || reg436[(4'hb):(1'h1)]))};
            end
          reg446 = forvar434;
        end
    end
  always
    @(posedge clk) begin
      if (wire107)
        begin
          reg447 <= ($signed(((|{reg444}) ?
                  ((reg427 << wire107) >>> (reg427 <= wire106)) : wire106[(4'hb):(1'h0)])) ?
              (!$unsigned(($unsigned(reg444) ?
                  (8'h9e) : (wire107 <= wire422)))) : (~^($signed({reg424,
                  reg445}) <= reg438)));
          for (forvar448 = (1'h0); (forvar448 < (2'h3)); forvar448 = (forvar448 + (1'h1)))
            begin
              reg449 = reg447[(1'h1):(1'h0)];
              reg450 <= (~reg427[(2'h3):(2'h3)]);
              reg451 <= {reg447};
              reg452 <= (({wire105[(4'h9):(2'h3)]} >>> (^(8'h9d))) ?
                  (^~(8'ha8)) : $unsigned($signed($unsigned(((8'hbd) >>> forvar448)))));
              reg453 <= ($unsigned($signed(wire105[(4'ha):(3'h4)])) ?
                  $signed($unsigned(reg450[(4'ha):(3'h4)])) : wire422[(2'h3):(1'h0)]);
            end
          reg454 <= (~|reg449);
          for (forvar455 = (1'h0); (forvar455 < (3'h4)); forvar455 = (forvar455 + (1'h1)))
            begin
              reg456 <= $unsigned(reg427[(1'h1):(1'h1)]);
              reg457 = (wire107 ?
                  ((wire107[(4'h9):(3'h5)] | (+reg445)) ^~ {{$unsigned(reg444)}}) : (reg456 ?
                      {((forvar448 ? reg452 : wire422) ?
                              $signed(wire107) : reg427),
                          {$unsigned((8'hb1))}} : ({$unsigned(reg447)} ?
                          reg424[(4'h9):(1'h0)] : $signed($signed(reg445)))));
              reg458 <= ($signed(reg451) ^ (^~{reg457[(1'h0):(1'h0)]}));
              reg459 = (|forvar448);
            end
          reg460 = $signed($signed(reg451[(4'hf):(4'h8)]));
        end
      else
        begin
          if ((~^(!{(reg460 | (8'ha1)), $signed({reg459, reg445})})))
            begin
              reg447 <= wire105;
              reg448 = reg456[(2'h3):(2'h3)];
              reg450 <= {(|(&((~&reg451) ?
                      $unsigned(reg459) : (wire105 ^~ forvar455)))),
                  $unsigned({$unsigned((reg451 ? reg452 : reg454))})};
            end
          else
            begin
              reg448 = (reg444 ?
                  ($signed({$unsigned((7'h4a))}) ?
                      wire422 : $signed(wire422)) : (wire105 ?
                      (&(forvar448 <<< reg457)) : reg459));
              reg449 = wire104[(4'h8):(1'h1)];
              reg455 = (($signed($signed($unsigned(reg454))) ?
                      ($unsigned($signed(forvar448)) ?
                          reg457 : $unsigned($unsigned(reg438))) : (~|$signed((~|wire106)))) ?
                  (($unsigned(reg447) == reg456[(1'h1):(1'h1)]) && ($signed(wire104[(4'h8):(4'h8)]) + (((7'h46) ~^ (8'hbb)) ?
                      (wire422 - forvar455) : $signed(reg448)))) : reg444[(5'h18):(5'h17)]);
              reg456 <= $unsigned($signed(reg456[(2'h3):(1'h0)]));
              reg458 <= (^~(^((^(reg456 ? reg456 : (8'haf))) || forvar455)));
            end
          for (forvar459 = (1'h0); (forvar459 < (2'h2)); forvar459 = (forvar459 + (1'h1)))
            begin
              reg461 <= forvar448[(4'hc):(3'h6)];
              reg462 <= (!(forvar459 != (reg457[(3'h5):(1'h1)] ?
                  $signed((reg456 ? reg438 : reg459)) : ({(8'hb0),
                      reg459} == reg450[(4'ha):(4'ha)]))));
            end
          reg463 = forvar459[(4'h9):(4'h8)];
          for (forvar464 = (1'h0); (forvar464 < (1'h0)); forvar464 = (forvar464 + (1'h1)))
            begin
              reg465 = $signed($signed((wire422 ?
                  reg445[(3'h5):(2'h2)] : $unsigned((reg453 ~^ reg452)))));
            end
        end
      reg466 <= reg451[(5'h12):(1'h1)];
      reg467 = reg427;
    end
  always
    @(posedge clk) begin
      for (forvar468 = (1'h0); (forvar468 < (2'h2)); forvar468 = (forvar468 + (1'h1)))
        begin
          for (forvar469 = (1'h0); (forvar469 < (2'h3)); forvar469 = (forvar469 + (1'h1)))
            begin
              reg470 = ({$unsigned(((reg445 | (8'hb7)) || $unsigned(reg452))),
                  $unsigned(reg466)} ~^ (reg450 ?
                  (8'hbc) : reg462[(2'h3):(2'h3)]));
              reg471 = $unsigned((reg450 & (!forvar469[(4'ha):(1'h0)])));
            end
          reg472 <= reg466;
          for (forvar473 = (1'h0); (forvar473 < (3'h4)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 = {((8'had) ?
                      (($signed(reg454) != (reg472 ?
                          reg456 : reg462)) && reg454[(5'h17):(2'h2)]) : wire422[(1'h0):(1'h0)]),
                  reg466[(3'h6):(1'h1)]};
              reg475 <= (forvar473 ?
                  (($unsigned((forvar468 ?
                      reg451 : reg424)) << $signed((reg470 ?
                      reg470 : reg466))) || $unsigned(($unsigned(reg444) ?
                      forvar469[(1'h1):(1'h1)] : $signed((8'hb0))))) : $unsigned(((~reg474) ?
                      ({forvar473, reg470} - $signed(reg451)) : ((reg447 ?
                          wire105 : reg458) ^ (+(8'hac))))));
              reg476 = $unsigned(reg453[(3'h5):(1'h0)]);
              reg477 <= $signed(((reg453 > reg450) ?
                  (^~reg451[(5'h16):(4'h8)]) : $signed((reg445 ?
                      wire105[(2'h2):(1'h1)] : (reg452 ? reg470 : reg447)))));
            end
        end
      reg478 <= $signed((!$unsigned(reg444)));
    end
  assign wire479 = $signed(((~^$signed((~^wire106))) == wire104[(4'h8):(3'h5)]));
  assign wire480 = $signed(reg447);
  always
    @(posedge clk) begin
      for (forvar481 = (1'h0); (forvar481 < (2'h2)); forvar481 = (forvar481 + (1'h1)))
        begin
          for (forvar482 = (1'h0); (forvar482 < (3'h4)); forvar482 = (forvar482 + (1'h1)))
            begin
              reg483 <= $unsigned($unsigned($signed(({reg451, wire422} ?
                  $signed((8'hbe)) : $signed(reg445)))));
              reg484 <= (wire107[(4'h8):(1'h1)] ?
                  (8'ha2) : $signed($unsigned((+(reg475 ? wire105 : reg475)))));
            end
          if (((^~(|(~^(wire480 ? wire479 : (8'hb0))))) ? wire480 : reg461))
            begin
              reg485 <= reg450[(4'ha):(4'ha)];
              reg486 <= $unsigned((($unsigned(reg484) ?
                  ((wire422 ? wire480 : wire106) ?
                      (reg472 ?
                          (8'hac) : wire106) : $unsigned(wire107)) : ($unsigned(reg444) & $unsigned((8'ha8)))) && (~&({wire422,
                  wire107} | $signed(wire104)))));
              reg487 <= wire422[(4'hd):(4'h9)];
              reg488 = ($signed(wire105[(4'h9):(3'h7)]) ?
                  (^reg438) : {$signed($signed((reg452 ? reg438 : reg458)))});
            end
          else
            begin
              reg485 <= (^~(({(&reg478)} ?
                  ((8'haa) ^ (~reg444)) : forvar482) != reg424[(4'hf):(4'hd)]));
              reg486 <= $unsigned((!($signed($unsigned(wire422)) ?
                  ((reg424 ? forvar481 : wire106) ?
                      $unsigned(forvar482) : (reg445 + reg487)) : $signed($unsigned(reg452)))));
            end
          reg489 <= {($signed($signed($signed(reg458))) ?
                  (^({wire422} ?
                      $unsigned(reg487) : reg462)) : $unsigned($unsigned((-wire422)))),
              $unsigned((^$unsigned($unsigned(reg462))))};
          if (($unsigned({(&(forvar482 >> reg450))}) >= ((|(reg475[(2'h2):(1'h0)] ?
              (wire422 <= forvar482) : $unsigned(reg484))) <<< reg452)))
            begin
              reg490 <= (+((^reg450) ?
                  wire107[(4'ha):(1'h1)] : $signed(($unsigned(forvar481) - reg489))));
              reg491 = reg475[(4'h8):(3'h5)];
            end
          else
            begin
              reg491 = ($signed($signed(reg483)) <<< ($unsigned(((reg450 ?
                      wire107 : reg462) >= (8'hbd))) ?
                  $signed($signed($signed(reg447))) : reg447[(3'h6):(3'h6)]));
              reg492 <= ((reg490 ?
                  forvar482 : $unsigned(((wire422 & reg489) ?
                      reg451 : $unsigned(reg475)))) ~^ $signed(wire422));
              reg493 <= (8'ha4);
              reg494 = $unsigned((wire480[(3'h4):(2'h3)] ?
                  reg488 : $signed({(reg466 ~^ wire106), (reg475 != reg453)})));
              reg495 = (({$signed(reg493[(3'h6):(3'h6)])} >>> ((&reg493[(1'h0):(1'h0)]) ?
                      $signed($unsigned(forvar481)) : ($signed(wire107) == $unsigned(reg490)))) ?
                  wire479 : (reg494 ?
                      reg488 : ($signed($signed(wire107)) ?
                          $signed((^~reg438)) : forvar482[(1'h0):(1'h0)])));
            end
        end
    end
  assign wire496 = (&reg438[(3'h6):(1'h0)]);
  always
    @(posedge clk) begin
      if (wire104)
        begin
          reg497 = ($unsigned(($signed({reg438, reg487}) ?
                  (8'h9f) : $signed((!(8'h9d))))) ?
              $signed((reg485[(4'h8):(1'h1)] - $unsigned((+reg427)))) : ((|{$unsigned(reg453)}) | $unsigned($unsigned(reg451))));
        end
      else
        begin
          for (forvar497 = (1'h0); (forvar497 < (2'h3)); forvar497 = (forvar497 + (1'h1)))
            begin
              reg498 = $unsigned($signed($unsigned((^reg489[(5'h10):(4'hc)]))));
              reg499 = {reg447[(4'ha):(4'ha)], (~reg452)};
              reg500 <= $unsigned($unsigned((~((wire106 && reg484) ?
                  reg483 : (+reg451)))));
              reg501 = reg490[(4'hc):(4'hb)];
            end
          for (forvar502 = (1'h0); (forvar502 < (3'h4)); forvar502 = (forvar502 + (1'h1)))
            begin
              reg503 = (reg477 ?
                  reg424 : {(!reg498[(4'h8):(1'h0)]),
                      $signed((~(reg450 * wire422)))});
            end
        end
      reg504 <= {(~|$unsigned((reg503 ?
              (reg438 ? reg489 : reg444) : reg503[(2'h3):(2'h2)]))),
          $unsigned($signed(($signed(wire479) ?
              (reg427 ? reg452 : reg503) : $unsigned(reg451))))};
    end
  always
    @(posedge clk) begin
      if ((($unsigned(wire479) * (reg487[(2'h3):(1'h0)] == reg466)) != reg466))
        begin
          reg505 <= wire105[(3'h6):(3'h6)];
          for (forvar506 = (1'h0); (forvar506 < (2'h3)); forvar506 = (forvar506 + (1'h1)))
            begin
              reg507 = {{((wire105 - (~|reg477)) >>> ((reg485 ?
                          wire479 : reg458) <= (7'h40)))}};
              reg508 = (reg452 >= (8'ha8));
              reg509 = (|(!$signed(((reg444 ^~ reg484) || reg462[(4'h8):(3'h6)]))));
            end
          reg510 <= ((reg486 ?
                  reg472 : ($unsigned(reg451[(4'hd):(4'hb)]) ?
                      {$signed((8'hb0)),
                          reg475[(4'h9):(3'h7)]} : {$signed(wire496)})) ?
              reg484 : reg445);
          if (((($unsigned(reg445[(3'h5):(1'h0)]) >>> reg427) <= $signed(((reg510 ?
              wire480 : reg445) >>> reg424[(3'h7):(2'h3)]))) - reg454))
            begin
              reg511 = reg485[(3'h7):(1'h1)];
            end
          else
            begin
              reg512 <= $signed(({((8'haf) <<< (reg451 + reg424))} ^~ {wire479}));
              reg513 <= ((~^(&$unsigned((7'h46)))) ?
                  $unsigned($unsigned((~|reg492[(2'h2):(2'h2)]))) : (-(-wire104)));
              reg514 = (~reg424);
            end
        end
      else
        begin
          for (forvar505 = (1'h0); (forvar505 < (1'h1)); forvar505 = (forvar505 + (1'h1)))
            begin
              reg506 <= (^~(($unsigned({(8'hb0)}) | ($signed((8'ha1)) ^ (wire479 ?
                      reg466 : (8'hb7)))) ?
                  (+reg489[(1'h1):(1'h0)]) : (reg510 - reg472)));
              reg507 = $signed({($unsigned(reg484) ?
                      ($signed(wire106) < wire480[(4'hc):(3'h7)]) : {(reg445 ^~ wire107),
                          ((8'hab) >> reg445)}),
                  (8'had)});
              reg510 <= $signed(reg453[(4'hf):(4'hb)]);
              reg511 = (wire496 ?
                  (reg454[(3'h5):(3'h4)] - reg424[(2'h2):(2'h2)]) : (((((8'h9e) ~^ reg444) ?
                              $signed(reg510) : {reg424, reg453}) ?
                          {$unsigned((8'haa))} : $unsigned($unsigned(reg475))) ?
                      $signed((-reg505)) : reg486[(4'h9):(3'h5)]));
            end
        end
      for (forvar515 = (1'h0); (forvar515 < (2'h3)); forvar515 = (forvar515 + (1'h1)))
        begin
          reg516 = $signed(wire105[(1'h1):(1'h0)]);
          reg517 = reg484[(4'hf):(4'h9)];
          for (forvar518 = (1'h0); (forvar518 < (2'h3)); forvar518 = (forvar518 + (1'h1)))
            begin
              reg519 = {$signed(reg462)};
              reg520 <= (reg509[(3'h5):(2'h2)] >> $unsigned($unsigned((|$unsigned(reg472)))));
              reg521 <= ({reg507[(3'h5):(3'h5)]} ?
                  (reg509 ^~ $unsigned((8'hb6))) : (((reg506[(1'h0):(1'h0)] + (wire107 > wire106)) ?
                          (reg486[(4'h8):(2'h3)] <<< (|(8'hac))) : {(reg513 + reg424),
                              (wire422 ? reg451 : reg511)}) ?
                      reg438[(2'h3):(1'h1)] : $signed({(^~reg512)})));
            end
          if ((+{(reg521 * ({reg514} == (^~forvar506))), (-{(~|reg506)})}))
            begin
              reg522 <= (reg445 ?
                  (wire422 ?
                      reg517[(2'h3):(2'h3)] : reg483[(5'h13):(5'h13)]) : (reg453[(5'h10):(4'h9)] ?
                      (^~reg486[(2'h2):(2'h2)]) : $signed({$unsigned(reg458),
                          reg487[(4'h8):(4'h8)]})));
              reg523 <= $unsigned((-reg504));
              reg524 = (~&$unsigned($unsigned($signed((reg486 ?
                  reg521 : reg509)))));
              reg525 = reg493[(3'h6):(2'h3)];
              reg526 = $unsigned(reg489);
            end
          else
            begin
              reg522 <= wire496;
            end
        end
      for (forvar527 = (1'h0); (forvar527 < (1'h1)); forvar527 = (forvar527 + (1'h1)))
        begin
          if (forvar515)
            begin
              reg528 <= wire105[(3'h4):(2'h3)];
              reg529 = {$unsigned(($signed($signed(reg517)) ?
                      $signed((reg477 && reg510)) : $signed((7'h4a))))};
              reg530 <= wire480[(5'h14):(3'h7)];
              reg531 <= reg451;
            end
          else
            begin
              reg528 <= reg477;
              reg530 <= reg472;
              reg532 = (8'hb0);
            end
          if (reg438[(4'h9):(2'h3)])
            begin
              reg533 = {$unsigned(((reg530[(1'h1):(1'h0)] != $signed(wire422)) ~^ reg532))};
            end
          else
            begin
              reg534 <= ((!wire480) ?
                  (reg525 ?
                      reg485[(1'h0):(1'h0)] : (~|(|reg526[(3'h7):(1'h1)]))) : (reg478 ?
                      $signed(((~|reg489) + (reg447 ?
                          reg513 : reg506))) : $unsigned(reg489)));
              reg535 = (reg453[(4'he):(3'h5)] >= $unsigned($signed((!(reg509 ?
                  reg506 : reg458)))));
            end
        end
    end
  module536 #() modinst643 (wire642, clk, reg500, reg534, reg456, reg512);
  always
    @(posedge clk) begin
      if (((7'h43) >= (reg472[(3'h7):(2'h2)] ?
          {$signed(reg484)} : reg513[(2'h2):(2'h2)])))
        begin
          reg644 = reg485[(2'h2):(1'h1)];
        end
      else
        begin
          if ((~(|reg444[(5'h11):(5'h10)])))
            begin
              reg645 <= reg534[(5'h12):(4'ha)];
            end
          else
            begin
              reg644 = (reg458[(1'h1):(1'h1)] < (7'h44));
              reg646 = reg453[(4'hf):(3'h6)];
            end
          reg647 = $unsigned(reg644[(1'h1):(1'h0)]);
        end
    end
  always
    @(posedge clk) begin
      reg648 = {{$signed($unsigned($signed(reg461)))},
          (~(~&(~$unsigned(wire422))))};
      for (forvar649 = (1'h0); (forvar649 < (3'h4)); forvar649 = (forvar649 + (1'h1)))
        begin
          reg650 = reg645[(4'h8):(1'h1)];
          reg651 = $signed(((reg530[(4'hc):(1'h1)] ?
              (8'hbf) : reg483) ^ $signed($unsigned(((8'hb9) ?
              reg477 : reg452)))));
          if ($unsigned((~reg445)))
            begin
              reg652 = $signed(($signed($unsigned(reg528[(4'hc):(3'h6)])) ~^ reg512));
              reg653 <= $signed($unsigned({reg648}));
              reg654 <= $unsigned(($signed($unsigned((|reg477))) ?
                  {$signed((~|wire480))} : {(~{reg653}),
                      ($signed(reg506) * reg520[(1'h1):(1'h0)])}));
            end
          else
            begin
              reg653 <= {(($unsigned($unsigned(reg522)) ?
                          reg454[(3'h7):(3'h4)] : reg475[(2'h3):(1'h0)]) ?
                      $unsigned((^~((8'hb7) >> wire479))) : reg453[(4'he):(3'h5)])};
              reg655 = $unsigned($signed((^reg648[(2'h2):(1'h0)])));
              reg656 = $signed({$signed(((&reg472) >>> $signed(reg489))),
                  $unsigned(reg530)});
              reg657 = reg447[(1'h0):(1'h0)];
            end
          reg658 = $signed(reg483);
          for (forvar659 = (1'h0); (forvar659 < (2'h3)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 <= wire479;
              reg661 = (^~(reg513[(2'h2):(1'h1)] ^~ reg452));
            end
        end
      for (forvar662 = (1'h0); (forvar662 < (1'h0)); forvar662 = (forvar662 + (1'h1)))
        begin
          if ((~|reg458[(1'h1):(1'h1)]))
            begin
              reg663 = $unsigned($unsigned($signed($signed((reg510 * reg451)))));
              reg664 = (8'hb1);
              reg665 <= reg658[(3'h7):(3'h5)];
              reg666 <= (reg478 * $signed($unsigned((reg523[(3'h4):(3'h4)] | (reg665 | wire642)))));
              reg667 <= (!((~|forvar659[(3'h4):(1'h0)]) ^~ (8'h9d)));
            end
          else
            begin
              reg665 <= ((reg651 << ($unsigned(reg504) <= $unsigned($unsigned((8'hb3))))) ?
                  ((!($unsigned(reg510) & $signed(reg534))) != (((!reg487) ?
                      $signed(reg475) : (reg461 ?
                          (8'ha6) : reg485)) < reg665[(2'h2):(2'h2)])) : reg500[(2'h2):(1'h0)]);
              reg668 = $unsigned((-(($unsigned((8'ha3)) ?
                      (reg492 ? reg490 : reg658) : ((8'h9d) < (7'h4a))) ?
                  ((reg485 ? wire106 : reg534) == (~&(8'ha7))) : ((reg650 ?
                      reg531 : reg512) & $unsigned(reg461)))));
              reg669 = $signed($signed($signed(((reg485 ? reg427 : reg506) ?
                  (+(8'hb7)) : $unsigned(reg451)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg670 = (&{reg472[(3'h5):(2'h3)], reg665[(1'h0):(1'h0)]});
      reg671 = {$unsigned((((wire422 ?
              reg447 : reg427) + $unsigned((7'h41))) << (reg666[(3'h7):(2'h3)] && (reg490 >> (8'hb0))))),
          ($signed((!(~|reg478))) ? reg505 : $signed(reg489[(4'ha):(2'h3)]))};
      if ({(~^(^($unsigned(reg452) ? (~&reg534) : $unsigned(wire106)))),
          reg667})
        begin
          if ($unsigned((~reg522)))
            begin
              reg672 <= $unsigned(({(8'hb9)} * (wire642 ?
                  ((~|(8'hbd)) >> $unsigned(reg458)) : reg528)));
              reg673 = ((^~($signed((reg654 ? reg454 : reg475)) ?
                      $unsigned((reg477 && (8'ha4))) : $unsigned(reg472[(1'h0):(1'h0)]))) ?
                  ($unsigned({$unsigned(reg660)}) & (^~(^~(reg478 ~^ reg667)))) : (reg504[(4'hd):(4'hb)] - {((wire105 ?
                          reg505 : (8'h9e)) | (7'h47))}));
            end
          else
            begin
              reg672 <= ((reg487 ?
                  (+((reg424 >> reg478) - ((8'h9d) | wire104))) : $signed((8'h9d))) >> (($signed($unsigned(wire107)) >= reg521) ?
                  $signed(((reg506 ? reg672 : reg510) ?
                      (reg672 || reg424) : $unsigned(reg512))) : reg534[(5'h13):(4'h8)]));
              reg674 <= reg424[(3'h5):(2'h3)];
              reg675 = $unsigned(($signed(wire480[(5'h13):(4'h8)]) != (~^({reg505} + $signed(reg472)))));
              reg676 = $signed($unsigned($unsigned(reg506)));
            end
        end
      else
        begin
          for (forvar672 = (1'h0); (forvar672 < (1'h0)); forvar672 = (forvar672 + (1'h1)))
            begin
              reg673 = $signed((+$unsigned((|reg513))));
              reg675 = reg453[(4'hd):(3'h6)];
              reg676 = reg489[(4'he):(2'h3)];
              reg677 <= ($unsigned({reg450[(2'h3):(2'h2)]}) ?
                  (~reg486) : reg493);
              reg678 = (~|(8'hac));
            end
        end
      reg679 <= reg674[(1'h1):(1'h1)];
      for (forvar680 = (1'h0); (forvar680 < (1'h1)); forvar680 = (forvar680 + (1'h1)))
        begin
          if ((($signed((((8'hae) ? reg513 : reg500) ?
                  (wire107 ? reg510 : reg674) : ((8'ha1) && (8'ha7)))) ?
              (((~|reg485) >> reg670) >>> reg672) : (-(~^reg513[(1'h0):(1'h0)]))) || reg427))
            begin
              reg681 <= ((reg472[(4'h9):(2'h2)] ?
                      forvar680[(2'h2):(2'h2)] : $unsigned(reg506)) ?
                  reg466[(4'ha):(3'h4)] : reg528);
              reg682 <= reg675;
              reg683 <= reg500[(5'h11):(4'hb)];
            end
          else
            begin
              reg681 <= $unsigned((+(-(~|reg681))));
              reg684 = (wire107[(3'h5):(2'h2)] ?
                  ((^reg427) ?
                      $signed((~^$signed(reg484))) : reg679[(1'h1):(1'h0)]) : (~|(reg485[(4'h9):(3'h6)] ?
                      (&$signed(reg452)) : reg472[(3'h7):(1'h1)])));
            end
          if (wire496)
            begin
              reg685 <= ((reg534[(4'hf):(4'hf)] ?
                  (($signed(reg475) | (wire480 >>> reg485)) != ((reg671 * reg490) ?
                      reg487[(2'h3):(2'h2)] : $signed(reg486))) : (!$unsigned($signed(reg490)))) ^ $signed(reg530));
              reg686 = $signed($unsigned((~|(^~(~|reg450)))));
            end
          else
            begin
              reg685 <= (~^wire107);
              reg686 = reg447;
              reg687 = $unsigned(wire480);
            end
          if ({(reg483[(4'hf):(4'h9)] - ($signed(reg483) ? reg485 : reg506)),
              (+(reg483 ~^ (8'hae)))})
            begin
              reg688 <= reg456;
              reg689 <= {reg523, (~&reg686)};
              reg690 = $unsigned($unsigned($signed(wire105[(3'h5):(2'h2)])));
              reg691 = (^~{reg653[(2'h2):(1'h1)]});
            end
          else
            begin
              reg690 = (forvar672 ?
                  (wire106[(1'h1):(1'h0)] ?
                      $unsigned({$signed(wire496),
                          reg504[(4'hb):(3'h4)]}) : reg453) : $signed($signed(((wire107 ?
                          reg445 : reg478) ?
                      $signed((8'hb3)) : reg444))));
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg447[(4'ha):(3'h5)])
        begin
          reg692 = ($signed(((((7'h43) + reg506) + (reg444 > (8'hb2))) ?
                  reg475[(3'h7):(2'h3)] : (reg492[(2'h3):(1'h1)] < reg683))) ?
              reg520 : $unsigned($signed(reg653[(1'h1):(1'h1)])));
        end
      else
        begin
          for (forvar692 = (1'h0); (forvar692 < (2'h3)); forvar692 = (forvar692 + (1'h1)))
            begin
              reg693 <= reg681;
            end
        end
      reg694 <= {wire480,
          (wire480[(3'h4):(2'h3)] ?
              reg466[(4'ha):(3'h6)] : $unsigned($unsigned((reg447 <<< reg454))))};
      for (forvar695 = (1'h0); (forvar695 < (1'h1)); forvar695 = (forvar695 + (1'h1)))
        begin
          if (reg453[(4'h9):(1'h1)])
            begin
              reg696 = (~^({reg454[(5'h10):(3'h4)], (7'h4a)} ?
                  (~&(8'hb7)) : reg493));
              reg697 = reg653;
            end
          else
            begin
              reg698 <= $signed(reg520);
              reg699 = wire480[(5'h10):(1'h0)];
              reg700 = $unsigned({(reg660[(1'h0):(1'h0)] ?
                      {$unsigned(reg451)} : reg531[(3'h7):(3'h4)])});
              reg701 = reg445[(3'h5):(2'h2)];
            end
          for (forvar702 = (1'h0); (forvar702 < (2'h3)); forvar702 = (forvar702 + (1'h1)))
            begin
              reg703 = ($signed($signed(reg451)) | $unsigned(wire480[(3'h7):(1'h0)]));
              reg704 = (wire104 ?
                  (reg477 ?
                      reg528 : ({(+reg493)} * ((reg483 ?
                          reg530 : reg454) <<< (^reg699)))) : $unsigned($unsigned($unsigned({reg667}))));
            end
          for (forvar705 = (1'h0); (forvar705 < (1'h0)); forvar705 = (forvar705 + (1'h1)))
            begin
              reg706 <= $unsigned($signed(((reg505[(4'h9):(1'h0)] ^ ((8'h9d) ?
                  reg681 : reg462)) < reg492)));
              reg707 <= $unsigned({reg438});
              reg708 = reg666;
              reg709 = reg703[(4'h8):(2'h2)];
              reg710 = reg424[(5'h14):(5'h11)];
            end
          reg711 <= ((^~{$signed((forvar692 * reg451)), {{reg444}}}) ?
              (~reg521) : $signed((^~{reg682})));
        end
      reg712 = (8'hb0);
      for (forvar713 = (1'h0); (forvar713 < (2'h2)); forvar713 = (forvar713 + (1'h1)))
        begin
          for (forvar714 = (1'h0); (forvar714 < (2'h3)); forvar714 = (forvar714 + (1'h1)))
            begin
              reg715 = reg665[(3'h4):(1'h0)];
              reg716 = $signed((~$unsigned((reg688[(4'hd):(4'hb)] | $unsigned(reg522)))));
              reg717 <= reg458;
              reg718 <= reg716;
            end
          reg719 = (reg444 == reg692);
          for (forvar720 = (1'h0); (forvar720 < (1'h1)); forvar720 = (forvar720 + (1'h1)))
            begin
              reg721 <= (reg486[(2'h3):(1'h1)] ?
                  $unsigned((-($signed(reg510) == $unsigned((8'ha5))))) : ($unsigned(({reg484,
                          reg450} ?
                      $unsigned(reg660) : (~reg475))) >> (((wire104 ~^ reg458) - (reg660 - (8'ha0))) ?
                      $unsigned((!forvar692)) : reg692)));
            end
          if ($signed(($unsigned({(|(8'ha1)),
              (reg717 >>> wire479)}) * (forvar720[(2'h2):(1'h0)] ?
              {(reg683 | reg654), {reg521}} : {$signed((8'h9e))}))))
            begin
              reg722 = (reg453 ?
                  (!reg447[(4'h9):(2'h3)]) : reg484[(4'hc):(4'h9)]);
            end
          else
            begin
              reg722 = reg534;
              reg723 = (-(reg453[(3'h5):(3'h4)] ^~ $signed($signed((8'ha9)))));
              reg724 <= reg698;
              reg725 = ((|wire480) - reg716[(2'h2):(1'h0)]);
              reg726 = reg709;
            end
        end
    end
  always
    @(posedge clk) begin
      if ((~|(8'ha8)))
        begin
          reg727 = {(reg424[(1'h0):(1'h0)] || (reg424 ?
                  reg451[(5'h14):(5'h10)] : ($unsigned(reg685) ?
                      reg493[(3'h7):(3'h4)] : (8'hb7))))};
        end
      else
        begin
          reg728 <= $signed(((^reg679[(2'h2):(2'h2)]) ?
              reg477[(4'hd):(4'h8)] : $signed(reg492[(3'h5):(2'h2)])));
          reg729 = (((^$unsigned($signed((8'hb9)))) >>> {((^wire106) != (reg512 - reg489)),
                  $signed(reg513)}) ?
              (-$unsigned(((reg693 ?
                  reg461 : reg505) || {reg505}))) : (~&reg707[(2'h3):(1'h0)]));
          if ($unsigned($signed($unsigned($unsigned((reg486 ?
              wire496 : reg522))))))
            begin
              reg730 <= $unsigned({wire106[(4'ha):(4'h8)]});
              reg731 <= (((~|((reg454 ? reg513 : reg456) ?
                  (~|wire496) : $signed(reg718))) ^ $signed((&wire479[(1'h0):(1'h0)]))) <<< (reg685 >>> $unsigned($signed({reg645}))));
              reg732 <= (($unsigned(((wire106 ?
                      reg505 : reg490) * reg731[(2'h2):(1'h1)])) | $unsigned((8'hab))) ?
                  $signed((^~(8'hba))) : (($signed((reg531 <= reg486)) != reg483) ?
                      (^~reg458[(3'h4):(1'h0)]) : reg681));
            end
          else
            begin
              reg730 <= ($unsigned(($signed($signed(reg504)) ^ ((reg510 ?
                      reg477 : reg523) || $signed(reg732)))) ?
                  $unsigned($signed({(reg677 == reg478)})) : $signed($unsigned(($unsigned((7'h47)) >= {(8'hb2),
                      reg466}))));
              reg731 <= $signed(reg688);
              reg732 <= (&(~^$signed($signed(reg730[(3'h6):(1'h0)]))));
              reg733 = (($signed((reg534 && reg486)) - reg685) ?
                  ($unsigned((+{reg504})) ~^ (reg645[(3'h4):(1'h0)] + (~^reg677))) : (reg484 - {reg450}));
              reg734 = (($signed($unsigned((reg730 ? reg505 : reg520))) ?
                  ((~(reg729 ?
                      reg462 : reg478)) > $unsigned(reg717)) : (|reg487)) <<< $signed($signed(reg504[(4'he):(3'h7)])));
            end
          for (forvar735 = (1'h0); (forvar735 < (2'h3)); forvar735 = (forvar735 + (1'h1)))
            begin
              reg736 = (~&((reg531[(4'hd):(4'h8)] < (+$signed((8'hbf)))) - $unsigned((reg711[(4'hb):(3'h4)] ?
                  reg484 : $unsigned(reg521)))));
              reg737 = $signed($unsigned($signed(reg727[(3'h6):(3'h5)])));
            end
        end
      reg738 = reg438[(3'h6):(1'h0)];
      reg739 = ($unsigned((wire107[(4'h8):(3'h6)] ? (!(~^reg472)) : reg683)) ?
          $signed((reg530[(4'hd):(4'hb)] <= $unsigned((+reg727)))) : ((~|(^~$unsigned(reg453))) ?
              (($unsigned(reg707) ?
                  (-(7'h49)) : {reg450}) - $signed(reg729[(5'h10):(4'h8)])) : ({{reg707,
                      reg500},
                  reg456[(3'h7):(2'h3)]} == $signed($unsigned(reg485)))));
      reg740 <= reg674[(4'h8):(1'h1)];
      if ((reg694[(1'h1):(1'h1)] ?
          ({($signed(reg707) ^~ (7'h4a))} ?
              $signed((~(8'hbd))) : (|reg740[(2'h2):(1'h0)])) : (^~((reg739[(3'h7):(1'h0)] ?
              (~^(8'ha9)) : (&(8'ha1))) >>> reg456))))
        begin
          for (forvar741 = (1'h0); (forvar741 < (1'h0)); forvar741 = (forvar741 + (1'h1)))
            begin
              reg742 = reg487;
              reg743 = (~|reg681[(5'h13):(4'hd)]);
            end
          for (forvar744 = (1'h0); (forvar744 < (2'h2)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 <= (((({reg666} ? reg522[(3'h5):(3'h5)] : (~|reg653)) ?
                      {$unsigned(reg530),
                          (reg492 ~^ reg711)} : $signed((|wire422))) ?
                  $signed(((reg706 ?
                      reg424 : reg737) > (~^(7'h47)))) : (~^$unsigned(reg711))) < (~|$unsigned((8'hb5))));
              reg746 = {((+(~(reg645 * (8'ha8)))) ?
                      (~^((-reg447) ?
                          (reg454 ?
                              reg718 : reg718) : $unsigned(reg462))) : $unsigned($signed($signed(reg653)))),
                  {$signed((reg682 != (~reg688))), reg689[(2'h2):(1'h1)]}};
            end
          reg747 = ($signed(reg427[(3'h7):(3'h6)]) - reg485[(4'h9):(1'h1)]);
          reg748 <= $unsigned(reg523[(2'h2):(1'h0)]);
        end
      else
        begin
          reg741 = $unsigned($signed(reg478));
          reg742 = (~|($signed(((reg484 && wire105) != $unsigned(reg451))) + $signed((~(reg674 * (8'h9d))))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar749 = (1'h0); (forvar749 < (3'h4)); forvar749 = (forvar749 + (1'h1)))
        begin
          reg750 = reg654;
          if (reg490[(4'hf):(3'h4)])
            begin
              reg751 = $signed((^~reg492));
              reg752 <= ((reg461 ?
                      $signed((~((8'ha9) & reg456))) : $unsigned($unsigned($signed(reg732)))) ?
                  (~&reg682[(2'h3):(1'h1)]) : (&$signed(((reg534 ?
                          reg523 : reg693) ?
                      (wire107 ? reg453 : reg427) : reg682))));
            end
          else
            begin
              reg752 <= $signed(($unsigned({{wire106, (8'h9d)}}) ?
                  {({(8'haa)} ? $unsigned(reg707) : $signed(reg520)),
                      reg478[(3'h4):(2'h3)]} : $unsigned(reg477[(5'h10):(5'h10)])));
              reg753 <= ((($signed((reg683 != reg645)) ?
                          reg653[(1'h0):(1'h0)] : $signed({(8'hb5)})) ?
                      $unsigned($unsigned((reg505 && reg528))) : ($signed(reg721) >> $unsigned((reg487 ?
                          reg534 : reg694)))) ?
                  (|$unsigned((|$signed(reg745)))) : (~|($unsigned($signed(reg500)) <<< (reg685[(4'hd):(3'h6)] ?
                      $unsigned(wire104) : (reg748 ? reg486 : reg522)))));
              reg754 = reg665[(3'h5):(1'h1)];
              reg755 <= $signed(({(~|(wire480 ? wire104 : reg732))} ?
                  reg530 : (8'hbd)));
            end
          reg756 = ({($signed((8'h9d)) ?
                  reg728 : $unsigned(((8'hab) ? reg493 : reg450))),
              ((reg456 ?
                  reg427 : (reg752 ^ reg732)) != reg513[(1'h0):(1'h0)])} <= reg492);
          for (forvar757 = (1'h0); (forvar757 < (1'h0)); forvar757 = (forvar757 + (1'h1)))
            begin
              reg758 <= $signed($unsigned($signed(reg721)));
              reg759 = (+reg456);
              reg760 <= $signed(reg694[(1'h1):(1'h1)]);
              reg761 <= (reg472[(4'h9):(2'h2)] - $unsigned(reg660));
            end
        end
      if ((~^{((reg462 ? (reg698 ? reg500 : reg753) : (reg534 ^~ forvar757)) ?
              ((|reg523) ? reg672[(1'h0):(1'h0)] : reg755) : reg665)}))
        begin
          reg762 = (|reg490);
        end
      else
        begin
          reg763 <= (reg461[(5'h11):(4'h8)] << ($signed({(8'hbe)}) ?
              $unsigned(reg718[(3'h5):(2'h3)]) : (^~reg759)));
        end
    end
  assign wire764 = (^~reg456);
  always
    @(posedge clk) begin
      for (forvar765 = (1'h0); (forvar765 < (3'h4)); forvar765 = (forvar765 + (1'h1)))
        begin
          reg766 = ((|$signed(reg451[(4'ha):(4'h9)])) || reg681);
          reg767 = $signed(reg672[(3'h4):(3'h4)]);
        end
      for (forvar768 = (1'h0); (forvar768 < (2'h3)); forvar768 = (forvar768 + (1'h1)))
        begin
          for (forvar769 = (1'h0); (forvar769 < (2'h2)); forvar769 = (forvar769 + (1'h1)))
            begin
              reg770 = reg685[(4'hc):(4'hc)];
            end
          reg771 = $signed($unsigned($unsigned($unsigned((reg485 ^ reg745)))));
        end
      for (forvar772 = (1'h0); (forvar772 < (1'h0)); forvar772 = (forvar772 + (1'h1)))
        begin
          for (forvar773 = (1'h0); (forvar773 < (1'h0)); forvar773 = (forvar773 + (1'h1)))
            begin
              reg774 <= ({(8'hb4),
                  reg477[(1'h0):(1'h0)]} | (($unsigned(reg732) ?
                  ({reg475,
                      reg645} != wire106[(2'h3):(1'h1)]) : $signed($unsigned(reg665))) || (8'ha8)));
            end
          reg775 <= (~|((reg438[(3'h4):(3'h4)] ^~ $signed(reg752[(2'h3):(2'h2)])) ?
              reg452 : ($signed((reg681 ? wire480 : reg732)) ?
                  $unsigned({reg683}) : reg760)));
          reg776 <= ({reg718} == (^~reg451));
          for (forvar777 = (1'h0); (forvar777 < (1'h0)); forvar777 = (forvar777 + (1'h1)))
            begin
              reg778 = reg760[(2'h2):(1'h1)];
              reg779 <= reg717;
              reg780 = reg438[(4'h9):(4'h8)];
              reg781 <= {{reg456[(1'h0):(1'h0)], ($unsigned((8'hba)) ^ reg654)},
                  ($unsigned($unsigned($unsigned(reg451))) ?
                      $signed({(8'hbc)}) : reg718)};
              reg782 = ($signed((((reg531 ? reg689 : reg745) >>> wire107) ?
                      $unsigned((reg452 ? reg484 : forvar777)) : ({reg478,
                          (7'h46)} - {reg456}))) ?
                  (+($unsigned((reg445 >>> reg654)) ?
                      $signed($unsigned(reg677)) : {reg717[(3'h7):(3'h4)]})) : {(reg711 * $signed((reg693 ^~ reg758)))});
            end
          reg783 <= (~&$unsigned($unsigned($unsigned((reg693 != reg740)))));
        end
      if (((reg522[(1'h1):(1'h1)] ?
              $unsigned($unsigned(reg688[(5'h16):(2'h2)])) : reg724) ?
          (((+reg774) ?
              $unsigned((~^reg776)) : ((+reg707) ?
                  $unsigned((8'hbf)) : (reg462 >= reg487))) ^~ reg522[(4'h8):(3'h4)]) : {(((forvar765 ?
                      reg512 : reg427) * reg693) ?
                  $unsigned(((8'hb1) ? wire480 : reg513)) : $signed({reg698,
                      (7'h42)}))}))
        begin
          reg784 <= (&{{(~|$unsigned(reg478))}});
          reg785 <= $unsigned(wire104[(3'h5):(2'h3)]);
          if ((&{reg775}))
            begin
              reg786 <= (($signed(reg665) ?
                  {((^~reg781) <<< reg505[(1'h1):(1'h1)])} : reg660[(3'h5):(1'h1)]) >>> (~&$unsigned((wire479[(2'h2):(2'h2)] >>> reg782[(1'h1):(1'h1)]))));
              reg787 = {$unsigned($signed((+$signed(reg778)))),
                  $unsigned($unsigned($signed((-(7'h46)))))};
              reg788 <= (-(reg707[(4'hb):(4'h8)] << $unsigned(((&reg688) && (forvar768 ?
                  reg484 : reg530)))));
            end
          else
            begin
              reg786 <= ($signed({forvar773[(4'hc):(1'h0)]}) ?
                  reg711[(4'hf):(2'h2)] : (^~$unsigned(reg753)));
              reg787 = ($unsigned(((~^reg660[(3'h5):(3'h4)]) ?
                  reg730 : {$signed((8'hb5))})) < ((forvar777 == $unsigned(((8'hac) ?
                      (8'hab) : wire106))) ?
                  ($unsigned(reg771[(3'h6):(2'h3)]) ?
                      $signed((^reg504)) : ((reg779 & reg447) - wire104)) : (($unsigned(reg534) ?
                      {reg487, reg452} : ((8'hb1) ?
                          reg521 : reg778)) != (+reg782[(2'h2):(1'h1)]))));
              reg789 = reg506;
              reg790 = $signed(reg475);
              reg791 <= wire764;
            end
          reg792 <= reg728[(2'h2):(1'h1)];
          if (reg758)
            begin
              reg793 = {(&(8'h9c))};
              reg794 = (8'ha7);
            end
          else
            begin
              reg793 = (&reg781[(1'h0):(1'h0)]);
              reg794 = $unsigned($unsigned($signed((~|(reg461 ?
                  reg793 : reg782)))));
              reg795 <= ($signed($unsigned(((reg444 != reg724) >>> $unsigned((8'hb0))))) ?
                  ($unsigned(($signed(reg766) - $unsigned(reg753))) >> $signed($unsigned({reg475}))) : ((~(|(~|reg444))) ?
                      $signed(reg654[(1'h1):(1'h1)]) : (+forvar772[(4'ha):(3'h4)])));
              reg796 <= $signed(($unsigned((~&$signed((8'hb9)))) ?
                  reg784 : $signed(reg458[(3'h4):(2'h2)])));
              reg797 <= $signed(wire479);
            end
        end
      else
        begin
          reg784 <= reg793[(4'hf):(3'h5)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module536  (y, clk, wire540, wire539, wire538, wire537);
  output wire [(32'h555):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h17):(1'h0)] wire540;
  input wire [(5'h16):(1'h0)] wire539;
  input wire signed [(5'h14):(1'h0)] wire538;
  input wire [(3'h7):(1'h0)] wire537;
  wire [(5'h13):(1'h0)] wire641;
  wire [(3'h6):(1'h0)] wire628;
  wire signed [(5'h10):(1'h0)] wire627;
  wire signed [(5'h11):(1'h0)] wire605;
  wire [(5'h18):(1'h0)] wire581;
  wire signed [(4'ha):(1'h0)] wire580;
  wire signed [(4'hf):(1'h0)] wire569;
  reg signed [(3'h6):(1'h0)] reg640 = (1'h0);
  reg [(5'h11):(1'h0)] reg639 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg636 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg635 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg633 = (1'h0);
  reg [(5'h18):(1'h0)] reg631 = (1'h0);
  reg [(4'hc):(1'h0)] reg630 = (1'h0);
  reg [(5'h15):(1'h0)] reg621 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg616 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg614 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg613 = (1'h0);
  reg [(4'ha):(1'h0)] reg612 = (1'h0);
  reg [(5'h10):(1'h0)] reg609 = (1'h0);
  reg [(5'h18):(1'h0)] reg607 = (1'h0);
  reg [(2'h3):(1'h0)] reg606 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg603 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg602 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg598 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg597 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg596 = (1'h0);
  reg [(5'h11):(1'h0)] reg595 = (1'h0);
  reg [(4'hb):(1'h0)] reg594 = (1'h0);
  reg [(4'ha):(1'h0)] reg590 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg588 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg586 = (1'h0);
  reg [(5'h12):(1'h0)] reg578 = (1'h0);
  reg [(2'h2):(1'h0)] reg575 = (1'h0);
  reg [(4'he):(1'h0)] reg573 = (1'h0);
  reg [(5'h16):(1'h0)] reg567 = (1'h0);
  reg [(3'h4):(1'h0)] reg566 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg561 = (1'h0);
  reg [(5'h18):(1'h0)] reg560 = (1'h0);
  reg [(4'hb):(1'h0)] reg555 = (1'h0);
  reg [(5'h13):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg553 = (1'h0);
  reg [(3'h7):(1'h0)] reg550 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg546 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg543 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg541 = (1'h0);
  reg [(5'h17):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg637 = (1'h0);
  reg [(2'h2):(1'h0)] reg634 = (1'h0);
  reg [(5'h13):(1'h0)] reg632 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg629 = (1'h0);
  reg [(4'h8):(1'h0)] reg626 = (1'h0);
  reg signed [(4'he):(1'h0)] reg625 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg624 = (1'h0);
  reg [(5'h12):(1'h0)] reg623 = (1'h0);
  reg [(5'h17):(1'h0)] reg622 = (1'h0);
  reg [(5'h10):(1'h0)] reg620 = (1'h0);
  reg [(4'h9):(1'h0)] reg619 = (1'h0);
  reg [(4'h8):(1'h0)] reg618 = (1'h0);
  reg [(4'hd):(1'h0)] reg617 = (1'h0);
  reg [(4'hd):(1'h0)] reg615 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg611 = (1'h0);
  reg [(5'h16):(1'h0)] reg610 = (1'h0);
  reg [(3'h5):(1'h0)] reg608 = (1'h0);
  reg [(3'h4):(1'h0)] reg604 = (1'h0);
  reg [(2'h2):(1'h0)] reg601 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg600 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg599 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg593 = (1'h0);
  reg [(5'h12):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg591 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg589 = (1'h0);
  reg [(5'h15):(1'h0)] reg587 = (1'h0);
  reg [(5'h16):(1'h0)] forvar585 = (1'h0);
  reg [(5'h18):(1'h0)] reg584 = (1'h0);
  reg [(5'h17):(1'h0)] forvar583 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg582 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg579 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg577 = (1'h0);
  reg [(5'h13):(1'h0)] forvar576 = (1'h0);
  reg [(5'h10):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg572 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg571 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar570 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg568 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg565 = (1'h0);
  reg [(5'h18):(1'h0)] reg563 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar562 = (1'h0);
  reg [(4'hd):(1'h0)] reg559 = (1'h0);
  reg [(5'h11):(1'h0)] reg558 = (1'h0);
  reg [(5'h11):(1'h0)] reg557 = (1'h0);
  reg [(5'h18):(1'h0)] reg556 = (1'h0);
  reg [(5'h13):(1'h0)] reg552 = (1'h0);
  reg [(4'ha):(1'h0)] reg551 = (1'h0);
  reg [(3'h4):(1'h0)] reg549 = (1'h0);
  reg [(2'h3):(1'h0)] reg548 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg547 = (1'h0);
  reg [(4'h8):(1'h0)] reg545 = (1'h0);
  reg [(5'h11):(1'h0)] forvar544 = (1'h0);
  reg [(3'h4):(1'h0)] reg542 = (1'h0);
  assign y = {wire641,
                 wire628,
                 wire627,
                 wire605,
                 wire581,
                 wire580,
                 wire569,
                 reg640,
                 reg639,
                 reg636,
                 reg635,
                 reg633,
                 reg631,
                 reg630,
                 reg621,
                 reg616,
                 reg614,
                 reg613,
                 reg612,
                 reg609,
                 reg607,
                 reg606,
                 reg603,
                 reg602,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 reg590,
                 reg588,
                 reg586,
                 reg578,
                 reg575,
                 reg573,
                 reg567,
                 reg566,
                 reg564,
                 reg561,
                 reg560,
                 reg555,
                 reg554,
                 reg553,
                 reg550,
                 reg546,
                 reg543,
                 reg541,
                 reg638,
                 reg637,
                 reg634,
                 reg632,
                 reg629,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 reg615,
                 reg611,
                 reg610,
                 reg608,
                 reg604,
                 reg601,
                 reg600,
                 reg599,
                 reg593,
                 reg592,
                 reg591,
                 reg589,
                 reg587,
                 forvar585,
                 reg584,
                 forvar583,
                 reg582,
                 reg579,
                 reg577,
                 forvar576,
                 reg574,
                 reg572,
                 reg571,
                 forvar570,
                 reg568,
                 reg565,
                 reg563,
                 forvar562,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 reg552,
                 reg551,
                 reg549,
                 reg548,
                 reg547,
                 reg545,
                 forvar544,
                 reg542,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg541 <= (($signed(wire537[(2'h2):(1'h1)]) <<< $unsigned((^wire540[(5'h10):(2'h3)]))) ?
          $unsigned((~|($signed(wire540) || $unsigned(wire538)))) : ($unsigned($signed($signed(wire537))) <<< $unsigned(((&wire538) ?
              $unsigned(wire540) : $unsigned(wire537)))));
      reg542 = $unsigned($unsigned(wire539[(5'h15):(3'h6)]));
      reg543 <= $unsigned((wire539 ? (8'haf) : (&{$signed(reg541)})));
      for (forvar544 = (1'h0); (forvar544 < (1'h0)); forvar544 = (forvar544 + (1'h1)))
        begin
          reg545 = forvar544;
          if ($unsigned($signed($signed(($signed(reg545) ?
              (-wire539) : forvar544)))))
            begin
              reg546 <= $unsigned($unsigned((~reg543[(4'h8):(1'h0)])));
            end
          else
            begin
              reg546 <= (|{($unsigned((!reg541)) ?
                      $unsigned((-reg543)) : {wire539,
                          reg542[(2'h2):(1'h1)]})});
              reg547 = $signed((wire538[(5'h14):(4'h8)] ?
                  (({reg541} ?
                          (wire538 ?
                              reg542 : wire538) : wire539[(4'hb):(2'h2)]) ?
                      (+(8'hb4)) : $signed((wire537 ?
                          reg541 : wire537))) : $unsigned({(reg545 ~^ reg542),
                      wire537})));
              reg548 = wire537[(1'h1):(1'h1)];
              reg549 = ((!((8'hbf) ?
                  $signed($signed((8'ha5))) : $signed((reg543 > reg542)))) <<< $signed({$signed((reg541 >= reg548))}));
            end
          reg550 <= ((-wire538[(3'h7):(3'h4)]) >>> (!(~&(~|reg543[(4'h8):(4'h8)]))));
          reg551 = $unsigned((7'h42));
          if (reg541[(1'h1):(1'h0)])
            begin
              reg552 = $unsigned(((^~$unsigned($unsigned(wire537))) ?
                  reg541[(2'h2):(1'h0)] : forvar544));
              reg553 <= ($signed((((reg546 - reg547) << (reg542 ?
                          wire539 : reg541)) ?
                      $unsigned(wire537) : reg543[(2'h3):(2'h2)])) ?
                  ($signed($unsigned($signed(reg542))) ?
                      $signed(((~reg542) ?
                          (reg542 * reg547) : $signed(reg545))) : ({reg546[(1'h1):(1'h0)]} ?
                          (!(|(8'ha2))) : (^~$signed(reg549)))) : ($unsigned((^reg541[(3'h4):(1'h1)])) ?
                      (wire537[(1'h0):(1'h0)] != (^~wire538[(4'h9):(4'h9)])) : {{reg551[(3'h4):(1'h0)]},
                          (~|{reg551})}));
              reg554 <= (reg545[(3'h4):(3'h4)] ^~ $signed(((forvar544 - (|reg548)) ?
                  $signed((reg553 ? reg551 : reg546)) : (~|(reg541 ?
                      forvar544 : reg549)))));
            end
          else
            begin
              reg552 = reg553[(3'h6):(3'h4)];
            end
        end
      if (reg554[(2'h2):(1'h1)])
        begin
          reg555 <= {forvar544[(5'h11):(4'h8)]};
        end
      else
        begin
          reg556 = ({(($unsigned(reg549) ? (&(8'ha7)) : (8'ha9)) ?
                      $signed($unsigned(reg542)) : ((forvar544 ?
                          (8'hae) : (8'hb9)) - $signed((8'hab)))),
                  (~|((reg550 ? wire537 : wire537) ?
                      (reg552 << reg547) : forvar544))} ?
              reg546 : (forvar544 >>> reg554));
          if (reg550[(2'h2):(1'h0)])
            begin
              reg557 = reg553;
              reg558 = (&$unsigned($signed($signed(wire537[(3'h5):(3'h4)]))));
              reg559 = {((reg557[(5'h11):(3'h6)] + {$unsigned((8'hbf))}) ?
                      reg542[(2'h2):(1'h1)] : $signed(reg547))};
            end
          else
            begin
              reg560 <= $unsigned($signed(wire540[(3'h6):(1'h1)]));
              reg561 <= wire537[(1'h1):(1'h0)];
            end
          for (forvar562 = (1'h0); (forvar562 < (2'h3)); forvar562 = (forvar562 + (1'h1)))
            begin
              reg563 = ((~&(~^(^wire539[(4'h9):(3'h4)]))) ?
                  {(($unsigned(wire540) != (reg557 & forvar562)) & reg551[(3'h4):(1'h0)])} : (reg555[(4'hb):(3'h6)] ?
                      reg542 : reg557));
              reg564 <= reg541[(2'h3):(1'h1)];
              reg565 = {$unsigned(($unsigned($signed(reg560)) ?
                      (((8'hbe) << reg543) == (reg563 != (8'hbb))) : {$unsigned(reg556),
                          $signed(wire540)})),
                  (reg550[(3'h4):(1'h1)] ? reg553 : reg554)};
              reg566 <= wire537[(2'h2):(1'h0)];
              reg567 <= (-$signed({(((8'had) ? reg564 : reg564) ?
                      reg565[(3'h5):(3'h4)] : $signed(reg546))}));
            end
          reg568 = ((!($signed(reg554[(5'h12):(5'h10)]) - (&reg551))) * (~$unsigned({(reg560 ^~ reg554)})));
        end
    end
  assign wire569 = (reg553[(4'ha):(3'h6)] ?
                       ((|{$unsigned(reg543), (reg550 ? reg541 : reg541)}) ?
                           ((reg561[(4'h9):(4'h8)] ?
                               (reg553 ?
                                   reg541 : reg567) : reg555) - ((~&reg553) == (reg550 ^ reg541))) : $unsigned(reg561)) : (+((-reg560) >> $unsigned((wire540 - reg546)))));
  always
    @(posedge clk) begin
      for (forvar570 = (1'h0); (forvar570 < (2'h3)); forvar570 = (forvar570 + (1'h1)))
        begin
          reg571 = ({$signed({{reg561}}),
                  $signed(($signed(reg541) ? $signed(wire540) : (8'ha5)))} ?
              {{$unsigned((~|reg567)),
                      (-(reg550 > wire540))}} : ($unsigned($unsigned((^~(8'hb5)))) ?
                  $unsigned($unsigned((reg541 ?
                      reg561 : wire537))) : $unsigned(((reg566 << reg541) && (wire540 ^~ reg555)))));
          if ((reg571[(1'h0):(1'h0)] ?
              $signed(reg543[(2'h3):(2'h2)]) : ($unsigned(wire569) ?
                  ((~^(reg554 ? reg555 : wire538)) ?
                      ((8'hb5) || (|reg543)) : $signed((8'ha2))) : $signed($unsigned((&wire538))))))
            begin
              reg572 = reg553[(4'hb):(1'h1)];
              reg573 <= $signed(wire538);
            end
          else
            begin
              reg572 = reg573[(4'hd):(4'hb)];
              reg573 <= ((((^~((7'h49) ? forvar570 : reg567)) ?
                      {{reg553,
                              reg543}} : (+$unsigned(wire537))) ^~ $unsigned(wire538[(2'h2):(1'h0)])) ?
                  $signed($unsigned($signed($unsigned(reg572)))) : ($signed((~(~|reg553))) >> wire569[(4'hf):(4'h9)]));
              reg574 = ($signed((!(~&reg561[(5'h15):(5'h11)]))) ?
                  forvar570[(5'h12):(3'h6)] : (($signed((reg567 >>> reg573)) && ($signed(reg541) ?
                      $signed(wire538) : (reg541 ?
                          reg555 : (8'hbc)))) ^ reg571[(3'h5):(1'h0)]));
            end
          reg575 <= reg546;
        end
      for (forvar576 = (1'h0); (forvar576 < (1'h0)); forvar576 = (forvar576 + (1'h1)))
        begin
          reg577 = (($signed((forvar576[(3'h7):(3'h4)] ?
                  $unsigned(reg550) : (7'h48))) ?
              {(-reg546[(4'h8):(3'h7)]),
                  reg573[(1'h1):(1'h1)]} : {($signed(reg543) ~^ reg573)}) * reg543);
          reg578 <= {reg555, wire538};
        end
      reg579 = ($signed($signed({{reg541}})) ?
          $signed($signed(wire537)) : reg564[(1'h1):(1'h0)]);
    end
  assign wire580 = reg575;
  assign wire581 = (wire537[(1'h0):(1'h0)] ?
                       ({($unsigned(wire538) ~^ ((8'hbf) >>> reg550))} ?
                           ($signed((^reg564)) >> $signed((reg541 ?
                               reg555 : wire540))) : (~&$unsigned(wire540))) : wire538[(5'h11):(4'hf)]);
  always
    @(posedge clk) begin
      reg582 = wire580[(4'h8):(3'h7)];
      for (forvar583 = (1'h0); (forvar583 < (1'h1)); forvar583 = (forvar583 + (1'h1)))
        begin
          reg584 = reg566;
          for (forvar585 = (1'h0); (forvar585 < (1'h1)); forvar585 = (forvar585 + (1'h1)))
            begin
              reg586 <= (~&(^~reg560[(4'hd):(4'hc)]));
              reg587 = $unsigned((reg573[(4'he):(4'h9)] ?
                  reg564[(3'h4):(2'h3)] : $signed($signed((reg554 != reg567)))));
              reg588 <= wire540[(1'h1):(1'h1)];
            end
        end
      reg589 = reg584[(3'h5):(3'h4)];
      if ((|(^$signed(((wire580 & (7'h43)) ?
          (wire580 ? reg561 : (8'hb0)) : wire539)))))
        begin
          reg590 <= ((({{reg543, reg550}} ?
              $signed((~|reg589)) : ((reg550 || reg573) ?
                  (reg543 > reg578) : $unsigned(wire537))) | reg582[(3'h6):(1'h0)]) & $signed($unsigned((~|wire581))));
        end
      else
        begin
          if ((~|$unsigned($signed($signed($signed(reg541))))))
            begin
              reg591 = (reg553 ?
                  (&$signed((~&reg553))) : $unsigned($signed($unsigned((forvar585 == reg588)))));
              reg592 = (~&((+reg587) ?
                  (reg566 ?
                      {$unsigned(reg561)} : (8'hb8)) : (reg588[(2'h2):(1'h1)] < reg587)));
              reg593 = (({{$unsigned(reg561), $signed(wire580)},
                          ($unsigned(reg591) - $signed(reg586))} ?
                      wire539 : $signed($signed((reg587 >= reg564)))) ?
                  (^~$unsigned(wire540)) : $unsigned(reg591));
              reg594 <= reg564[(3'h4):(1'h0)];
            end
          else
            begin
              reg590 <= reg575[(1'h0):(1'h0)];
              reg591 = (8'hb3);
            end
          if ({$unsigned((-reg587[(4'he):(2'h3)]))})
            begin
              reg595 <= $signed(($unsigned(wire538[(3'h7):(3'h4)]) ?
                  ($unsigned((wire539 | reg564)) ?
                      (~^{wire580,
                          reg584}) : reg593) : $signed($signed($unsigned(reg555)))));
            end
          else
            begin
              reg595 <= $signed(wire537);
              reg596 <= (8'hbb);
              reg597 <= (^~((7'h40) ?
                  ((~^(~|reg564)) ?
                      $signed((reg589 || reg594)) : (reg567[(4'hb):(4'h8)] - reg546)) : reg564[(3'h4):(2'h2)]));
              reg598 <= ($unsigned(reg592) * $signed({(~{wire581, wire540})}));
              reg599 = $unsigned($signed($unsigned(($unsigned(wire537) | (reg554 ?
                  reg567 : wire580)))));
            end
          if ($signed(($unsigned(((reg560 || reg573) ?
              $unsigned(wire538) : $signed(reg587))) << reg546)))
            begin
              reg600 = reg575;
              reg601 = ($unsigned((({wire538} ~^ {(8'hbd)}) > (^~$signed(reg543)))) ?
                  (reg575 ?
                      $unsigned($signed((reg575 <<< reg550))) : ($unsigned(reg599[(3'h7):(2'h2)]) ?
                          ($signed(reg590) ?
                              (+reg573) : $unsigned(reg573)) : $signed(reg553))) : $signed($signed($signed($unsigned(reg593)))));
              reg602 <= (^reg598);
            end
          else
            begin
              reg602 <= (8'h9f);
              reg603 <= $signed((reg578[(3'h5):(2'h2)] < (({reg597, wire538} ?
                      reg582 : {wire538}) ?
                  wire580[(4'ha):(2'h3)] : ($signed(reg601) ?
                      (reg543 + (7'h44)) : reg589[(2'h2):(2'h2)]))));
              reg604 = ($unsigned(reg541[(1'h1):(1'h0)]) >> ((+(((8'hb4) ?
                  reg564 : (8'h9f)) + reg598[(3'h6):(2'h3)])) == $unsigned(reg546[(3'h6):(3'h6)])));
            end
        end
    end
  assign wire605 = (reg555[(3'h6):(1'h1)] <= (&(8'ha8)));
  always
    @(posedge clk) begin
      reg606 <= reg560[(2'h2):(2'h2)];
      if ({wire605})
        begin
          if (((7'h44) | (~wire537)))
            begin
              reg607 <= wire537;
              reg608 = {(({$unsigned(wire605)} ?
                          (^~(wire605 & reg590)) : ($signed(reg550) ?
                              reg554[(3'h7):(2'h2)] : wire540)) ?
                      {((&reg560) ^ reg603[(3'h6):(3'h4)]),
                          reg588[(1'h1):(1'h0)]} : $signed(((7'h45) ^ (8'hbd))))};
              reg609 <= $unsigned(wire537[(3'h5):(3'h4)]);
              reg610 = $signed(reg573[(4'h9):(3'h5)]);
              reg611 = (wire580[(2'h3):(1'h1)] ?
                  reg575[(1'h0):(1'h0)] : (reg564 ?
                      $unsigned(((reg578 && reg567) + wire581[(5'h18):(4'hd)])) : $signed(reg575[(2'h2):(2'h2)])));
            end
          else
            begin
              reg608 = $signed(((($unsigned(wire581) == reg564[(2'h2):(1'h1)]) ?
                      $unsigned(reg573[(1'h0):(1'h0)]) : reg566) ?
                  wire580[(3'h6):(2'h3)] : $signed(wire539)));
              reg609 <= ((&(~|$unsigned({reg564, reg596}))) ?
                  wire581[(4'h8):(3'h6)] : reg610[(3'h7):(3'h6)]);
              reg612 <= ($unsigned($unsigned(reg595[(4'hc):(1'h1)])) ?
                  $signed($signed((reg609 || reg610[(5'h16):(4'h8)]))) : ((reg555 ?
                      wire537 : (reg588 & ((7'h44) ?
                          reg588 : reg598))) ^~ ($signed(reg595[(1'h1):(1'h0)]) ?
                      (^~reg602) : ((reg575 ? reg602 : reg553) ^ reg594))));
              reg613 <= (!$signed({$signed(reg541),
                  (reg602[(3'h4):(1'h0)] <<< (reg596 ? reg588 : reg588))}));
            end
          if (((-$signed((^~$unsigned((7'h44))))) <<< $unsigned(($signed({(7'h45)}) ?
              reg609[(3'h4):(2'h2)] : (^~(reg586 * reg603))))))
            begin
              reg614 <= reg567;
              reg615 = reg561;
              reg616 <= $unsigned({reg594,
                  (&$unsigned((reg564 ? reg615 : reg595)))});
            end
          else
            begin
              reg615 = ($unsigned((8'hbf)) ?
                  reg573[(1'h1):(1'h0)] : reg553[(3'h5):(1'h1)]);
              reg617 = {$signed((($unsigned(wire581) >> (~^reg596)) && $unsigned({wire540,
                      reg541}))),
                  (8'h9e)};
              reg618 = (((8'ha6) ?
                  reg602[(1'h0):(1'h0)] : $signed(($unsigned(reg594) ^ (reg612 ~^ reg543)))) >>> $unsigned($unsigned({((8'ha0) > reg586),
                  $signed(reg588)})));
              reg619 = ((((|wire539) ?
                  ($signed(reg575) ?
                      (wire540 ?
                          wire537 : reg618) : $signed(wire540)) : ((reg564 << reg554) ?
                      reg553 : $unsigned(reg553))) - ($unsigned($signed(reg546)) <= {reg618,
                  (reg554 ? reg602 : reg575)})) & {(+(wire539 ?
                      wire605 : reg555[(3'h6):(2'h3)]))});
              reg620 = $signed(reg603);
            end
        end
      else
        begin
          reg607 <= (($unsigned($unsigned((reg553 ?
                  (7'h49) : wire540))) != (((8'ha0) >> $unsigned(reg607)) * reg602[(1'h1):(1'h1)])) ?
              reg566[(1'h0):(1'h0)] : reg553);
          if ((~|$signed($signed(reg613))))
            begin
              reg609 <= {((reg554[(3'h7):(1'h0)] ?
                      reg606[(2'h3):(1'h0)] : (+(reg588 == wire569))) >>> reg609[(4'h9):(3'h5)])};
              reg612 <= (($unsigned(reg573[(4'h8):(3'h5)]) ?
                      (({reg620, reg612} + $unsigned((8'hb1))) ^~ ({reg553,
                              reg586} ?
                          wire569[(4'h8):(2'h2)] : reg620[(1'h0):(1'h0)])) : ((8'hae) <<< $signed(reg620))) ?
                  reg598 : (({{(8'ha3), reg608}, {reg541, reg543}} ?
                      (-$signed(reg610)) : reg597) <<< ($signed((reg555 ?
                      reg610 : reg617)) >>> (^$unsigned(reg608)))));
              reg613 <= (|($signed(reg607) ?
                  (reg618 ?
                      (reg603[(4'h8):(3'h5)] > ((7'h47) != reg614)) : {wire580}) : wire580[(4'h9):(3'h4)]));
              reg614 <= $unsigned($unsigned((!((reg597 ? reg611 : reg573) ?
                  {reg588} : (8'ha4)))));
            end
          else
            begin
              reg609 <= wire537;
              reg610 = (~&{$unsigned((~$unsigned((8'hb6))))});
            end
          reg616 <= $signed(reg616[(1'h0):(1'h0)]);
          if ({$unsigned((((~^reg586) & (reg546 ?
                  reg613 : reg617)) || reg596))})
            begin
              reg617 = reg550;
            end
          else
            begin
              reg621 <= $unsigned({$signed(((reg603 * (8'ha8)) * (reg614 ?
                      reg541 : reg603))),
                  $unsigned($unsigned((reg606 ? reg541 : (8'hb9))))});
              reg622 = (8'h9c);
              reg623 = {(wire539 && $signed((~&reg603))),
                  $signed({(reg541 << (|reg609)), (~^reg553[(4'h8):(3'h4)])})};
              reg624 = reg619;
              reg625 = $unsigned((({(reg543 - (8'hab)), (~&(8'hb1))} ?
                  (-((7'h44) || (8'hbc))) : reg550) & $unsigned(reg561)));
            end
          reg626 = (wire569[(4'he):(4'hb)] << reg603);
        end
    end
  assign wire627 = reg566[(2'h3):(1'h1)];
  assign wire628 = reg543[(3'h4):(2'h3)];
  always
    @(posedge clk) begin
      reg629 = reg612[(4'h9):(3'h4)];
    end
  always
    @(posedge clk) begin
      if (reg603)
        begin
          reg630 <= reg573[(4'hd):(3'h7)];
        end
      else
        begin
          reg630 <= (&$unsigned($signed({reg606, wire581})));
          reg631 <= reg607[(4'hb):(1'h1)];
          reg632 = wire569;
          reg633 <= (+(~|(&(~reg561[(3'h7):(3'h7)]))));
          if ((reg606[(2'h3):(1'h0)] ?
              reg546[(2'h2):(1'h1)] : $unsigned(reg588)))
            begin
              reg634 = (|wire628);
              reg635 <= (8'haf);
              reg636 <= (wire605 <= wire540[(4'h9):(3'h6)]);
              reg637 = $signed($signed(reg573[(3'h4):(1'h0)]));
            end
          else
            begin
              reg634 = $unsigned((|(-{{(8'hae)}})));
              reg637 = $unsigned(reg590[(2'h2):(2'h2)]);
              reg638 = $unsigned((reg541 - (8'ha7)));
              reg639 <= (8'ha9);
              reg640 <= (~^reg632);
            end
        end
    end
  assign wire641 = $unsigned(reg594);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module108
#(parameter param421 = (~(((((8'ha0) ? (8'h9f) : (8'h9d)) & ((8'hac) ? (8'h9e) : (8'hbb))) ? (((7'h46) ? (8'hba) : (7'h45)) <<< (+(8'hb3))) : (8'hba)) ? (|((~|(7'h49)) ? (~(8'ha3)) : (&(7'h4a)))) : ((!{(8'hb3), (7'h43)}) - (^(-(8'hb6)))))))
(y, clk, wire113, wire112, wire111, wire110, wire109);
  output wire [(32'h10c9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire113;
  input wire signed [(4'hb):(1'h0)] wire112;
  input wire [(3'h6):(1'h0)] wire111;
  input wire [(4'hb):(1'h0)] wire110;
  input wire [(2'h3):(1'h0)] wire109;
  wire [(4'ha):(1'h0)] wire334;
  wire [(5'h15):(1'h0)] wire333;
  wire [(3'h7):(1'h0)] wire306;
  wire signed [(4'hb):(1'h0)] wire265;
  wire signed [(5'h13):(1'h0)] wire115;
  wire signed [(4'hc):(1'h0)] wire114;
  reg signed [(3'h4):(1'h0)] reg418 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg417 = (1'h0);
  reg [(2'h2):(1'h0)] reg416 = (1'h0);
  reg [(4'he):(1'h0)] reg415 = (1'h0);
  reg [(3'h4):(1'h0)] reg414 = (1'h0);
  reg [(5'h11):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg409 = (1'h0);
  reg [(4'ha):(1'h0)] reg405 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg399 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg396 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg394 = (1'h0);
  reg [(5'h13):(1'h0)] reg389 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg388 = (1'h0);
  reg [(5'h14):(1'h0)] reg386 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg381 = (1'h0);
  reg [(5'h10):(1'h0)] reg379 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg375 = (1'h0);
  reg [(3'h5):(1'h0)] reg374 = (1'h0);
  reg [(4'hb):(1'h0)] reg373 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg370 = (1'h0);
  reg [(3'h6):(1'h0)] reg366 = (1'h0);
  reg [(4'hf):(1'h0)] reg363 = (1'h0);
  reg [(4'ha):(1'h0)] reg360 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg357 = (1'h0);
  reg [(5'h11):(1'h0)] reg355 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg353 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg352 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg349 = (1'h0);
  reg [(4'he):(1'h0)] reg348 = (1'h0);
  reg [(3'h6):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg340 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg336 = (1'h0);
  reg [(3'h6):(1'h0)] reg332 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg325 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg323 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg322 = (1'h0);
  reg [(4'hd):(1'h0)] reg321 = (1'h0);
  reg [(4'h9):(1'h0)] reg320 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg318 = (1'h0);
  reg [(2'h3):(1'h0)] reg317 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg314 = (1'h0);
  reg [(5'h18):(1'h0)] reg313 = (1'h0);
  reg [(4'hc):(1'h0)] reg312 = (1'h0);
  reg [(3'h4):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg310 = (1'h0);
  reg [(2'h2):(1'h0)] reg308 = (1'h0);
  reg [(3'h7):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg305 = (1'h0);
  reg [(4'h8):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg299 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg295 = (1'h0);
  reg [(5'h14):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg291 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg287 = (1'h0);
  reg [(4'hf):(1'h0)] reg286 = (1'h0);
  reg [(2'h2):(1'h0)] reg283 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg279 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg276 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg274 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg273 = (1'h0);
  reg [(4'hf):(1'h0)] reg271 = (1'h0);
  reg [(4'hd):(1'h0)] reg270 = (1'h0);
  reg [(4'hc):(1'h0)] reg267 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg263 = (1'h0);
  reg signed [(4'he):(1'h0)] reg256 = (1'h0);
  reg [(4'hf):(1'h0)] reg261 = (1'h0);
  reg [(5'h14):(1'h0)] reg260 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg259 = (1'h0);
  reg [(4'he):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg248 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg246 = (1'h0);
  reg [(3'h7):(1'h0)] reg245 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg243 = (1'h0);
  reg [(5'h13):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg240 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg239 = (1'h0);
  reg [(4'hb):(1'h0)] reg236 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg232 = (1'h0);
  reg [(5'h14):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg224 = (1'h0);
  reg [(4'hc):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg222 = (1'h0);
  reg [(2'h2):(1'h0)] reg219 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg218 = (1'h0);
  reg [(3'h5):(1'h0)] reg215 = (1'h0);
  reg [(5'h16):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg209 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg208 = (1'h0);
  reg [(5'h18):(1'h0)] reg206 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg205 = (1'h0);
  reg [(5'h15):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg197 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg193 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg189 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg188 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg186 = (1'h0);
  reg [(5'h11):(1'h0)] reg182 = (1'h0);
  reg [(4'he):(1'h0)] reg178 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg177 = (1'h0);
  reg [(5'h14):(1'h0)] reg176 = (1'h0);
  reg [(5'h18):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg172 = (1'h0);
  reg [(3'h5):(1'h0)] reg171 = (1'h0);
  reg [(4'he):(1'h0)] reg170 = (1'h0);
  reg [(3'h7):(1'h0)] reg163 = (1'h0);
  reg [(4'ha):(1'h0)] reg169 = (1'h0);
  reg [(4'ha):(1'h0)] reg168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg164 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg154 = (1'h0);
  reg [(2'h2):(1'h0)] reg153 = (1'h0);
  reg [(5'h14):(1'h0)] reg152 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg151 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg150 = (1'h0);
  reg [(5'h16):(1'h0)] reg148 = (1'h0);
  reg [(4'hc):(1'h0)] reg146 = (1'h0);
  reg [(3'h4):(1'h0)] reg138 = (1'h0);
  reg [(5'h18):(1'h0)] reg136 = (1'h0);
  reg [(5'h10):(1'h0)] reg135 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg125 = (1'h0);
  reg [(5'h13):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg420 = (1'h0);
  reg [(4'hb):(1'h0)] reg419 = (1'h0);
  reg [(4'hb):(1'h0)] reg413 = (1'h0);
  reg [(5'h18):(1'h0)] reg412 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg411 = (1'h0);
  reg [(4'hf):(1'h0)] forvar403 = (1'h0);
  reg [(4'he):(1'h0)] reg410 = (1'h0);
  reg [(5'h13):(1'h0)] reg408 = (1'h0);
  reg [(2'h3):(1'h0)] forvar407 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg406 = (1'h0);
  reg [(4'hf):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg400 = (1'h0);
  reg [(5'h16):(1'h0)] forvar397 = (1'h0);
  reg [(5'h14):(1'h0)] forvar395 = (1'h0);
  reg [(5'h16):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg392 = (1'h0);
  reg [(5'h13):(1'h0)] forvar391 = (1'h0);
  reg [(3'h4):(1'h0)] forvar390 = (1'h0);
  reg [(5'h12):(1'h0)] reg387 = (1'h0);
  reg [(3'h5):(1'h0)] reg385 = (1'h0);
  reg [(4'hc):(1'h0)] reg383 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg382 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg380 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg378 = (1'h0);
  reg [(4'hb):(1'h0)] forvar377 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg376 = (1'h0);
  reg [(3'h4):(1'h0)] forvar372 = (1'h0);
  reg [(2'h3):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg369 = (1'h0);
  reg [(4'ha):(1'h0)] reg368 = (1'h0);
  reg [(4'hb):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg365 = (1'h0);
  reg [(5'h17):(1'h0)] reg364 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg362 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg361 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar359 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg358 = (1'h0);
  reg [(5'h12):(1'h0)] reg356 = (1'h0);
  reg [(4'hf):(1'h0)] forvar354 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg351 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg350 = (1'h0);
  reg [(5'h17):(1'h0)] forvar347 = (1'h0);
  reg [(5'h17):(1'h0)] reg346 = (1'h0);
  reg [(5'h16):(1'h0)] reg345 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg342 = (1'h0);
  reg [(3'h7):(1'h0)] forvar341 = (1'h0);
  reg [(5'h13):(1'h0)] reg339 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg338 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar337 = (1'h0);
  reg [(4'hd):(1'h0)] reg335 = (1'h0);
  reg [(3'h7):(1'h0)] reg330 = (1'h0);
  reg [(3'h5):(1'h0)] reg329 = (1'h0);
  reg [(4'ha):(1'h0)] reg327 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar326 = (1'h0);
  reg [(3'h4):(1'h0)] forvar324 = (1'h0);
  reg [(5'h12):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg316 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg315 = (1'h0);
  reg [(4'h8):(1'h0)] forvar308 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg309 = (1'h0);
  reg [(3'h5):(1'h0)] reg304 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg301 = (1'h0);
  reg signed [(4'he):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar298 = (1'h0);
  reg [(5'h17):(1'h0)] reg297 = (1'h0);
  reg [(4'hf):(1'h0)] reg294 = (1'h0);
  reg [(3'h5):(1'h0)] forvar293 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar289 = (1'h0);
  reg [(5'h11):(1'h0)] forvar288 = (1'h0);
  reg [(5'h16):(1'h0)] reg285 = (1'h0);
  reg [(5'h18):(1'h0)] reg284 = (1'h0);
  reg [(5'h10):(1'h0)] forvar282 = (1'h0);
  reg [(5'h17):(1'h0)] reg281 = (1'h0);
  reg [(4'hc):(1'h0)] reg280 = (1'h0);
  reg [(4'hc):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg277 = (1'h0);
  reg [(4'he):(1'h0)] reg275 = (1'h0);
  reg [(3'h4):(1'h0)] forvar272 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg269 = (1'h0);
  reg [(5'h13):(1'h0)] forvar268 = (1'h0);
  reg [(4'h9):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg264 = (1'h0);
  reg [(5'h12):(1'h0)] reg262 = (1'h0);
  reg [(5'h18):(1'h0)] reg253 = (1'h0);
  reg [(5'h10):(1'h0)] reg258 = (1'h0);
  reg [(4'he):(1'h0)] reg257 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar256 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar253 = (1'h0);
  reg [(5'h11):(1'h0)] reg251 = (1'h0);
  reg [(3'h6):(1'h0)] reg244 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg241 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg238 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg237 = (1'h0);
  reg [(4'h8):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar233 = (1'h0);
  reg [(3'h6):(1'h0)] reg231 = (1'h0);
  reg [(2'h2):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar226 = (1'h0);
  reg [(5'h18):(1'h0)] reg230 = (1'h0);
  reg [(3'h6):(1'h0)] reg228 = (1'h0);
  reg [(4'hd):(1'h0)] forvar227 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg226 = (1'h0);
  reg [(5'h11):(1'h0)] reg216 = (1'h0);
  reg [(5'h18):(1'h0)] reg225 = (1'h0);
  reg [(3'h7):(1'h0)] reg221 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg220 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg217 = (1'h0);
  reg [(5'h13):(1'h0)] forvar216 = (1'h0);
  reg [(5'h11):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg212 = (1'h0);
  reg [(4'h9):(1'h0)] reg211 = (1'h0);
  reg [(4'hc):(1'h0)] reg210 = (1'h0);
  reg [(4'hc):(1'h0)] reg207 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar203 = (1'h0);
  reg [(4'hf):(1'h0)] reg202 = (1'h0);
  reg [(4'ha):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg198 = (1'h0);
  reg [(5'h17):(1'h0)] reg196 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg194 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg192 = (1'h0);
  reg [(5'h12):(1'h0)] reg191 = (1'h0);
  reg [(5'h15):(1'h0)] forvar190 = (1'h0);
  reg [(4'hc):(1'h0)] reg187 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg185 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg184 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg183 = (1'h0);
  reg [(5'h15):(1'h0)] reg181 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg180 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar179 = (1'h0);
  reg [(4'hd):(1'h0)] reg175 = (1'h0);
  reg [(5'h17):(1'h0)] reg173 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar167 = (1'h0);
  reg [(4'hb):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg167 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar166 = (1'h0);
  reg [(4'h9):(1'h0)] forvar163 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg162 = (1'h0);
  reg [(4'h9):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg160 = (1'h0);
  reg [(4'he):(1'h0)] reg159 = (1'h0);
  reg [(5'h13):(1'h0)] reg158 = (1'h0);
  reg [(5'h10):(1'h0)] reg157 = (1'h0);
  reg [(5'h18):(1'h0)] reg156 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar155 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg149 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg147 = (1'h0);
  reg [(5'h18):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar144 = (1'h0);
  reg [(5'h16):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg141 = (1'h0);
  reg [(5'h15):(1'h0)] forvar140 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg139 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg137 = (1'h0);
  reg [(3'h5):(1'h0)] forvar133 = (1'h0);
  reg [(4'hf):(1'h0)] forvar132 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg130 = (1'h0);
  reg [(5'h17):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg128 = (1'h0);
  reg [(4'ha):(1'h0)] reg127 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg124 = (1'h0);
  reg [(4'hb):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar122 = (1'h0);
  reg [(3'h6):(1'h0)] forvar116 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg122 = (1'h0);
  reg [(4'hc):(1'h0)] reg121 = (1'h0);
  reg [(5'h17):(1'h0)] reg120 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg116 = (1'h0);
  assign y = {wire334,
                 wire333,
                 wire306,
                 wire265,
                 wire115,
                 wire114,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg407,
                 reg409,
                 reg405,
                 reg403,
                 reg402,
                 reg401,
                 reg399,
                 reg398,
                 reg396,
                 reg394,
                 reg389,
                 reg388,
                 reg386,
                 reg384,
                 reg381,
                 reg379,
                 reg375,
                 reg374,
                 reg373,
                 reg370,
                 reg366,
                 reg363,
                 reg360,
                 reg357,
                 reg355,
                 reg353,
                 reg352,
                 reg349,
                 reg348,
                 reg343,
                 reg340,
                 reg336,
                 reg332,
                 reg331,
                 reg328,
                 reg325,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg318,
                 reg317,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg308,
                 reg307,
                 reg305,
                 reg303,
                 reg299,
                 reg296,
                 reg295,
                 reg292,
                 reg291,
                 reg287,
                 reg286,
                 reg283,
                 reg279,
                 reg276,
                 reg274,
                 reg273,
                 reg271,
                 reg270,
                 reg267,
                 reg263,
                 reg256,
                 reg261,
                 reg260,
                 reg259,
                 reg252,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg243,
                 reg242,
                 reg240,
                 reg239,
                 reg236,
                 reg232,
                 reg229,
                 reg224,
                 reg223,
                 reg222,
                 reg219,
                 reg218,
                 reg215,
                 reg214,
                 reg209,
                 reg208,
                 reg206,
                 reg205,
                 reg201,
                 reg199,
                 reg197,
                 reg195,
                 reg193,
                 reg189,
                 reg188,
                 reg186,
                 reg182,
                 reg178,
                 reg177,
                 reg176,
                 reg174,
                 reg172,
                 reg171,
                 reg170,
                 reg163,
                 reg169,
                 reg168,
                 reg165,
                 reg164,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg148,
                 reg146,
                 reg138,
                 reg136,
                 reg135,
                 reg134,
                 reg131,
                 reg126,
                 reg125,
                 reg119,
                 reg118,
                 reg117,
                 reg420,
                 reg419,
                 reg413,
                 reg412,
                 reg411,
                 forvar403,
                 reg410,
                 reg408,
                 forvar407,
                 reg406,
                 reg404,
                 reg400,
                 forvar397,
                 forvar395,
                 reg393,
                 reg392,
                 forvar391,
                 forvar390,
                 reg387,
                 reg385,
                 reg383,
                 reg382,
                 reg380,
                 reg378,
                 forvar377,
                 reg376,
                 forvar372,
                 reg371,
                 reg369,
                 reg368,
                 reg367,
                 reg365,
                 reg364,
                 reg362,
                 reg361,
                 forvar359,
                 reg358,
                 reg356,
                 forvar354,
                 reg351,
                 reg350,
                 forvar347,
                 reg346,
                 reg345,
                 reg344,
                 reg342,
                 forvar341,
                 reg339,
                 reg338,
                 forvar337,
                 reg335,
                 reg330,
                 reg329,
                 reg327,
                 forvar326,
                 forvar324,
                 reg319,
                 reg316,
                 reg315,
                 forvar308,
                 reg309,
                 reg304,
                 reg302,
                 reg301,
                 reg300,
                 forvar298,
                 reg297,
                 reg294,
                 forvar293,
                 reg290,
                 forvar289,
                 forvar288,
                 reg285,
                 reg284,
                 forvar282,
                 reg281,
                 reg280,
                 reg278,
                 reg277,
                 reg275,
                 forvar272,
                 reg269,
                 forvar268,
                 reg266,
                 reg264,
                 reg262,
                 reg253,
                 reg258,
                 reg257,
                 forvar256,
                 reg255,
                 reg254,
                 forvar253,
                 reg251,
                 reg244,
                 reg241,
                 reg238,
                 reg237,
                 reg235,
                 reg234,
                 forvar233,
                 reg231,
                 reg227,
                 forvar226,
                 reg230,
                 reg228,
                 forvar227,
                 reg226,
                 reg216,
                 reg225,
                 reg221,
                 reg220,
                 reg217,
                 forvar216,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg207,
                 reg204,
                 forvar203,
                 reg202,
                 reg200,
                 reg198,
                 reg196,
                 reg194,
                 reg192,
                 reg191,
                 forvar190,
                 reg187,
                 reg185,
                 reg184,
                 reg183,
                 reg181,
                 reg180,
                 forvar179,
                 reg175,
                 reg173,
                 forvar167,
                 reg166,
                 reg167,
                 forvar166,
                 forvar163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 forvar155,
                 reg149,
                 reg147,
                 reg145,
                 forvar144,
                 reg143,
                 reg142,
                 reg141,
                 forvar140,
                 reg139,
                 reg137,
                 forvar133,
                 forvar132,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg124,
                 reg123,
                 forvar122,
                 forvar116,
                 reg122,
                 reg121,
                 reg120,
                 reg116,
                 (1'h0)};
  assign wire114 = $unsigned($signed(((&$unsigned(wire112)) ?
                       ((^wire110) ?
                           (wire111 ? wire112 : wire111) : (wire113 ?
                               wire111 : wire113)) : wire111)));
  assign wire115 = ((7'h4a) ?
                       $unsigned((~|(~^(wire109 && wire110)))) : wire112[(2'h3):(1'h1)]);
  always
    @(posedge clk) begin
      if (($unsigned(((+(wire111 ? wire115 : wire109)) ?
              (wire113 ?
                  wire113[(1'h0):(1'h0)] : $signed(wire109)) : wire112[(3'h4):(1'h0)])) ?
          $signed(wire110[(3'h7):(2'h3)]) : $signed($unsigned($unsigned(wire114)))))
        begin
          reg116 = (($unsigned({wire111, {wire115}}) <= wire110) ?
              {(8'ha0)} : {$signed($signed(wire110)), $unsigned((7'h43))});
          if ({reg116[(3'h4):(1'h0)], wire115[(3'h5):(2'h2)]})
            begin
              reg117 <= $unsigned((!wire113[(1'h1):(1'h1)]));
              reg118 <= (reg116 || wire113);
              reg119 <= $signed($unsigned((reg116 <<< wire113)));
              reg120 = (!$unsigned(({(^reg116), wire114} ?
                  ((&wire109) ^ $signed(wire109)) : {wire112[(4'h9):(3'h4)],
                      (reg116 ? wire113 : reg119)})));
            end
          else
            begin
              reg117 <= (((reg117[(4'h9):(4'h8)] ?
                      $unsigned((!(7'h4a))) : wire109) & $unsigned($signed($signed((8'ha6))))) ?
                  wire111 : $unsigned((+reg117)));
              reg118 <= {$signed(reg117[(4'h8):(2'h2)])};
            end
          reg121 = (^~(wire111[(3'h6):(3'h5)] ^~ reg116[(1'h0):(1'h0)]));
          reg122 = ($unsigned($signed(({wire115, reg118} - (reg120 ?
              reg118 : wire114)))) ^~ (($unsigned((~wire112)) <= (8'hb0)) & ($unsigned($unsigned(reg119)) || $unsigned($signed(wire115)))));
        end
      else
        begin
          for (forvar116 = (1'h0); (forvar116 < (1'h1)); forvar116 = (forvar116 + (1'h1)))
            begin
              reg117 <= ((|{wire114[(2'h2):(1'h0)],
                  (^~$signed(wire109))}) & $signed({$unsigned(reg118[(1'h1):(1'h1)])}));
            end
          reg120 = (-{((!(7'h45)) ? wire115 : $signed($signed(wire115))),
              $signed((wire112[(1'h0):(1'h0)] ? {forvar116} : (^~(7'h44))))});
          reg121 = $unsigned((|$unsigned($unsigned((&reg119)))));
          for (forvar122 = (1'h0); (forvar122 < (1'h1)); forvar122 = (forvar122 + (1'h1)))
            begin
              reg123 = ((-({(!wire113),
                      $unsigned(wire114)} + (|((8'haf) ~^ reg116)))) ?
                  wire114[(4'h9):(3'h5)] : forvar116);
              reg124 = $unsigned((!$unsigned((+(+(8'hbe))))));
            end
          if (reg117[(4'hf):(3'h4)])
            begin
              reg125 <= (+wire114[(2'h2):(1'h0)]);
              reg126 <= (~wire112);
            end
          else
            begin
              reg127 = (8'ha2);
              reg128 = wire111;
              reg129 = (~&$signed(reg117[(3'h6):(3'h6)]));
              reg130 = (-(8'hac));
              reg131 <= reg129;
            end
        end
      for (forvar132 = (1'h0); (forvar132 < (2'h2)); forvar132 = (forvar132 + (1'h1)))
        begin
          for (forvar133 = (1'h0); (forvar133 < (1'h0)); forvar133 = (forvar133 + (1'h1)))
            begin
              reg134 <= $unsigned($signed((-((reg123 << wire112) >= $signed(reg120)))));
              reg135 <= reg128[(5'h13):(3'h6)];
              reg136 <= (7'h46);
              reg137 = ($signed(({reg125[(2'h2):(1'h0)],
                  $signed(reg129)} >>> wire115)) || wire109[(1'h1):(1'h1)]);
              reg138 <= $signed(reg116[(2'h2):(2'h2)]);
            end
          reg139 = ($signed(reg131[(3'h5):(2'h2)]) ?
              reg120[(5'h16):(5'h10)] : $unsigned($signed($signed((reg116 ?
                  reg138 : reg134)))));
        end
      for (forvar140 = (1'h0); (forvar140 < (3'h4)); forvar140 = (forvar140 + (1'h1)))
        begin
          reg141 = (($unsigned((reg134[(4'he):(4'h9)] || (wire114 <= wire109))) ?
                  (($signed(reg128) == (|(8'h9f))) ?
                      (!(reg127 || reg136)) : {$signed(reg118)}) : (+$unsigned(reg124[(2'h2):(2'h2)]))) ?
              wire109[(2'h2):(1'h1)] : (~reg122));
          if (reg135[(4'ha):(1'h0)])
            begin
              reg142 = $signed(reg139);
              reg143 = forvar122;
            end
          else
            begin
              reg142 = $unsigned(($unsigned((forvar116 ?
                  wire109[(2'h2):(2'h2)] : (reg128 ?
                      reg134 : reg138))) ~^ wire112));
              reg143 = wire115;
            end
          for (forvar144 = (1'h0); (forvar144 < (2'h3)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 = (^forvar133[(1'h1):(1'h0)]);
              reg146 <= (~&((reg126[(4'ha):(3'h4)] ?
                  $unsigned((|reg136)) : reg126[(3'h5):(3'h4)]) ^ $unsigned((^~(reg119 ?
                  reg131 : forvar140)))));
              reg147 = $unsigned((^~(~|(~(reg126 ? reg121 : (8'hb5))))));
              reg148 <= ((reg141 ~^ ($unsigned(wire110) ?
                  reg119 : ($unsigned(reg123) ?
                      (~|reg138) : forvar122[(3'h5):(2'h3)]))) <<< $unsigned(reg124[(2'h2):(2'h2)]));
              reg149 = reg125;
            end
        end
      if ($signed($signed((($signed(wire109) >> (8'had)) <<< (reg119 ?
          $signed(reg139) : (!reg148))))))
        begin
          if ((~|($unsigned((!reg142[(4'h8):(3'h4)])) ?
              $signed((8'hb2)) : wire112)))
            begin
              reg150 <= $unsigned((reg138 == $unsigned(((+forvar133) ?
                  {reg131, reg125} : $unsigned((8'hb1))))));
              reg151 <= ((|{(^~(~^wire113)), reg142[(3'h4):(1'h1)]}) ?
                  (~|($unsigned(reg128) > wire111[(3'h5):(2'h2)])) : $signed(((!$signed(reg134)) || forvar144)));
              reg152 <= ($unsigned(reg143) ^ (($unsigned((reg134 || forvar122)) & $signed({(8'hb5),
                      forvar116})) ?
                  $signed($signed($unsigned(reg150))) : ({reg134,
                          $unsigned(reg151)} ?
                      $unsigned((wire115 == (7'h44))) : reg131[(1'h0):(1'h0)])));
              reg153 <= {(reg139 ? $unsigned({{(8'ha6)}}) : {reg143}),
                  $signed(reg119[(3'h5):(1'h1)])};
              reg154 <= $unsigned(forvar132);
            end
          else
            begin
              reg150 <= wire110[(4'hb):(1'h1)];
              reg151 <= $unsigned($signed({(reg125 >= reg127[(4'ha):(2'h3)]),
                  $unsigned({forvar122})}));
            end
          for (forvar155 = (1'h0); (forvar155 < (3'h4)); forvar155 = (forvar155 + (1'h1)))
            begin
              reg156 = forvar144[(5'h12):(4'hb)];
              reg157 = reg119;
            end
          if (reg151[(2'h3):(2'h3)])
            begin
              reg158 = (8'ha8);
              reg159 = $unsigned({{((&reg151) == reg145[(5'h16):(5'h13)])}});
              reg160 = $unsigned(forvar140[(4'hc):(3'h4)]);
            end
          else
            begin
              reg158 = reg121;
              reg159 = reg153[(2'h2):(1'h1)];
            end
        end
      else
        begin
          reg150 <= reg145[(5'h15):(5'h11)];
        end
    end
  always
    @(posedge clk) begin
      if (reg146)
        begin
          reg161 = reg125;
          reg162 = reg148;
          for (forvar163 = (1'h0); (forvar163 < (1'h0)); forvar163 = (forvar163 + (1'h1)))
            begin
              reg164 <= reg161[(3'h4):(1'h1)];
              reg165 <= wire113[(2'h2):(1'h0)];
            end
          for (forvar166 = (1'h0); (forvar166 < (1'h0)); forvar166 = (forvar166 + (1'h1)))
            begin
              reg167 = ((^{(8'ha0)}) ^ (({$unsigned(wire111), reg165} ?
                      $signed(reg150) : reg136) ?
                  ($unsigned({wire109}) ?
                      reg164 : ((reg138 != reg126) ?
                          {reg117, forvar163} : (reg136 ?
                              reg165 : wire110))) : {(!(reg148 < reg162)),
                      ((~reg164) > reg135)}));
              reg168 <= reg138[(3'h4):(2'h2)];
              reg169 <= ($signed($unsigned(((~wire111) ?
                  $unsigned(reg167) : reg152))) & wire113[(1'h1):(1'h0)]);
            end
        end
      else
        begin
          if ((-reg136[(5'h12):(4'hf)]))
            begin
              reg163 <= (wire110 < ((((wire113 ? forvar163 : reg151) ?
                          (^~reg134) : reg136[(3'h7):(3'h6)]) ?
                      ({(7'h4a)} << ((8'haf) ?
                          (8'hb7) : reg154)) : (reg151[(1'h0):(1'h0)] < reg148[(4'he):(2'h3)])) ?
                  $unsigned(reg146[(3'h6):(1'h0)]) : $unsigned($unsigned(reg150[(3'h4):(1'h1)]))));
              reg164 <= {(|reg163[(3'h6):(2'h3)]), $unsigned(reg135)};
            end
          else
            begin
              reg163 <= reg161[(1'h1):(1'h0)];
              reg164 <= (({($unsigned(reg154) ?
                          $unsigned(reg165) : $signed(reg131)),
                      reg138[(1'h1):(1'h1)]} ?
                  ({$unsigned(reg161),
                      (wire113 * reg117)} << $signed($unsigned((8'ha5)))) : (reg135[(4'hc):(3'h5)] ?
                      wire111 : wire114[(3'h6):(2'h2)])) >= (reg154[(3'h4):(1'h0)] ?
                  wire110 : $signed($unsigned((reg154 ? (8'hb1) : wire111)))));
              reg165 <= ((8'hb3) ~^ ({(&reg136[(1'h1):(1'h0)])} ?
                  $signed(reg131) : reg119));
            end
          reg166 = ($unsigned($unsigned(reg126[(4'ha):(3'h7)])) ?
              $unsigned(reg117[(4'h8):(2'h2)]) : $signed((reg148[(4'hc):(1'h0)] ?
                  ((-reg167) - (reg148 ? reg150 : reg168)) : (|(~&reg153)))));
          for (forvar167 = (1'h0); (forvar167 < (2'h2)); forvar167 = (forvar167 + (1'h1)))
            begin
              reg168 <= reg167;
            end
        end
      if (($unsigned($signed((~^(&wire112)))) ?
          {reg135} : (reg117[(4'hf):(1'h0)] + {(8'hb1),
              $signed($signed(forvar167))})))
        begin
          reg170 <= {(($unsigned($unsigned(wire112)) ^~ ($signed(reg161) ?
                  reg161[(2'h2):(1'h1)] : {reg118})) & {(8'hba)}),
              (reg167 ? {reg118, (&((8'hbb) ? reg126 : reg125))} : wire110)};
          reg171 <= (&$unsigned(($unsigned(wire109) != reg150)));
          if ($signed(reg171[(2'h3):(2'h2)]))
            begin
              reg172 <= {(-wire110[(1'h0):(1'h0)])};
              reg173 = $unsigned(({reg118} * (8'h9f)));
              reg174 <= (^~$signed(reg165[(2'h2):(2'h2)]));
              reg175 = $unsigned(wire113);
            end
          else
            begin
              reg173 = reg118;
              reg174 <= $signed($signed($signed((~|$unsigned(reg118)))));
              reg176 <= $unsigned((-$signed(((~^reg166) | (~(8'hac))))));
              reg177 <= $unsigned($signed((~reg150)));
              reg178 <= $unsigned((-({reg170[(1'h0):(1'h0)],
                  reg152[(5'h11):(1'h1)]} ~^ $unsigned(reg170[(1'h1):(1'h1)]))));
            end
          for (forvar179 = (1'h0); (forvar179 < (1'h0)); forvar179 = (forvar179 + (1'h1)))
            begin
              reg180 = ((8'hbd) ?
                  (~^((reg166[(4'h9):(3'h5)] > (8'hae)) || $unsigned((+(8'h9d))))) : {reg135,
                      reg150});
              reg181 = $unsigned(reg170[(1'h1):(1'h0)]);
              reg182 <= $unsigned(wire113);
              reg183 = (^reg174[(3'h5):(1'h0)]);
              reg184 = $unsigned(forvar166[(3'h4):(3'h4)]);
            end
          if ({($signed((|(reg134 ?
                  reg150 : wire110))) >>> ({forvar179[(1'h1):(1'h0)],
                  $signed(wire115)} | (^$unsigned(reg184)))),
              reg117[(4'hc):(4'hb)]})
            begin
              reg185 = $signed($signed(forvar167[(1'h1):(1'h1)]));
              reg186 <= (&forvar166[(3'h5):(2'h3)]);
            end
          else
            begin
              reg185 = reg117;
              reg187 = $unsigned({($signed({wire115, reg117}) ?
                      $signed(reg180[(3'h4):(3'h4)]) : (+$unsigned(reg118))),
                  $unsigned((8'hb6))});
              reg188 <= $unsigned(wire114[(3'h4):(2'h2)]);
              reg189 <= ($signed({reg183[(4'h8):(3'h5)],
                      $unsigned(reg150[(4'h8):(3'h4)])}) ?
                  ((reg161[(1'h1):(1'h1)] >= (((8'h9e) ? wire112 : reg136) ?
                          $unsigned(reg153) : reg171[(2'h2):(1'h1)])) ?
                      {((reg151 ? (8'hb2) : wire113) ?
                              wire110[(3'h7):(1'h0)] : $signed(reg186))} : $unsigned(wire109[(2'h2):(1'h1)])) : $unsigned($signed($unsigned(reg176))));
            end
        end
      else
        begin
          reg173 = $unsigned((~(($signed(wire111) ~^ reg165[(3'h7):(3'h5)]) - {$unsigned(reg169)})));
        end
      for (forvar190 = (1'h0); (forvar190 < (2'h2)); forvar190 = (forvar190 + (1'h1)))
        begin
          reg191 = $signed($unsigned((((reg175 ? reg152 : reg126) ?
                  (reg175 << (8'hb2)) : reg170) ?
              $signed($unsigned(forvar166)) : ((reg180 - reg176) ?
                  $signed(wire115) : $unsigned((8'hba))))));
          if ((((reg131[(2'h2):(1'h1)] ?
              (|(reg136 ~^ reg126)) : reg186) & $signed(($unsigned(wire112) ?
              reg131 : (~|(8'ha9))))) * $unsigned($unsigned((~^(-reg170))))))
            begin
              reg192 = (reg175[(4'hc):(3'h6)] < $unsigned(reg167));
              reg193 <= (forvar163 ?
                  (reg117 ?
                      reg131[(2'h3):(1'h0)] : $signed($unsigned({wire112}))) : (reg184 ?
                      $unsigned(reg181[(3'h4):(2'h2)]) : reg178[(3'h5):(1'h0)]));
              reg194 = (8'haf);
            end
          else
            begin
              reg192 = $unsigned(reg178);
            end
          if ((reg166[(4'ha):(2'h2)] ? reg169 : $signed(reg136)))
            begin
              reg195 <= reg181;
              reg196 = $signed($signed(reg163));
              reg197 <= ((forvar179 ~^ $signed((8'h9d))) ?
                  reg195[(3'h5):(2'h3)] : $unsigned($signed($unsigned((reg161 ?
                      (8'hb4) : reg150)))));
              reg198 = $unsigned((8'hbf));
            end
          else
            begin
              reg195 <= reg152[(4'h8):(3'h4)];
            end
          reg199 <= reg175;
          if (wire113)
            begin
              reg200 = $signed($unsigned(((reg131 ?
                      (reg193 ^ reg162) : $signed(reg168)) ?
                  $unsigned(((8'h9e) ? reg196 : reg146)) : reg135)));
            end
          else
            begin
              reg201 <= $signed($signed(reg189[(4'h8):(3'h4)]));
              reg202 = (reg198 + ($signed($signed((~^(8'hb4)))) < $signed(reg181)));
            end
        end
      for (forvar203 = (1'h0); (forvar203 < (2'h2)); forvar203 = (forvar203 + (1'h1)))
        begin
          if ($unsigned({$signed(($unsigned(wire113) > $signed(forvar167)))}))
            begin
              reg204 = (+(8'ha5));
              reg205 <= $signed($unsigned(reg162));
              reg206 <= $unsigned((^reg178));
              reg207 = reg119;
            end
          else
            begin
              reg204 = reg172;
              reg205 <= reg187[(4'hc):(3'h7)];
              reg206 <= reg201;
              reg207 = forvar190[(4'h8):(4'h8)];
            end
          reg208 <= reg161;
          if ((~&wire111))
            begin
              reg209 <= (~$unsigned($signed(((~^reg193) ^~ $unsigned(reg184)))));
              reg210 = reg208[(1'h0):(1'h0)];
              reg211 = reg188;
              reg212 = reg148[(4'he):(4'he)];
            end
          else
            begin
              reg209 <= reg208[(2'h3):(2'h2)];
            end
          reg213 = ($signed((reg152[(3'h5):(3'h4)] ^~ ((reg154 + reg212) ?
                  reg186 : $unsigned(reg163)))) ?
              (reg135 - (~^(~$unsigned(reg131)))) : ($signed(reg125[(3'h4):(2'h3)]) * (+(reg135[(2'h3):(2'h2)] <<< reg172[(2'h3):(2'h3)]))));
          reg214 <= (((7'h40) ?
                  (($signed(reg197) ?
                      $signed(reg138) : $signed((8'hbe))) + $signed((~|reg154))) : (&($unsigned(reg171) ?
                      wire109[(2'h3):(2'h3)] : $signed(reg182)))) ?
              ($unsigned((^reg117[(3'h4):(1'h0)])) < {($unsigned(wire115) <= $signed(reg209)),
                  (((8'ha7) ? (8'ha9) : forvar203) ?
                      wire110 : $unsigned(reg186))}) : $signed(reg191[(1'h0):(1'h0)]));
        end
      reg215 <= $unsigned($unsigned($unsigned(reg178[(4'hc):(2'h3)])));
    end
  always
    @(posedge clk) begin
      if ((reg186[(1'h1):(1'h1)] ?
          reg201[(2'h2):(1'h1)] : reg152[(2'h3):(1'h0)]))
        begin
          for (forvar216 = (1'h0); (forvar216 < (1'h1)); forvar216 = (forvar216 + (1'h1)))
            begin
              reg217 = reg168;
              reg218 <= {reg117};
            end
          if ({($unsigned({$unsigned(reg150)}) >= ({reg215[(1'h1):(1'h1)],
                      (~^(8'ha0))} ?
                  (((8'hbd) ? reg214 : reg135) | wire113) : (reg218 ?
                      ((8'hb7) ? reg193 : reg163) : reg174))),
              {$unsigned($unsigned(reg176[(2'h3):(1'h0)])),
                  ((~^reg119) >> {$unsigned(wire110), $signed(reg205)})}})
            begin
              reg219 <= {(reg138 ?
                      reg150[(1'h0):(1'h0)] : $unsigned((~^(8'hbc)))),
                  (^(($unsigned(wire115) ?
                      (-reg153) : $unsigned((8'hbb))) & $signed(reg164[(4'hf):(3'h5)])))};
              reg220 = $unsigned(reg174[(4'hf):(3'h5)]);
              reg221 = {$signed($unsigned(wire115)),
                  ((^~(!(reg168 ? (8'hbb) : reg217))) & reg189)};
            end
          else
            begin
              reg219 <= $unsigned(({wire115, reg188} ?
                  ({reg146[(4'h9):(3'h5)], (reg176 ? reg218 : wire115)} ?
                      (~|(!reg164)) : reg117[(3'h7):(1'h0)]) : (8'hbc)));
              reg222 <= (^{($signed((reg206 >= reg146)) ~^ reg170)});
              reg223 <= wire113[(2'h3):(2'h2)];
              reg224 <= (~|{forvar216, $signed(reg186)});
              reg225 = reg170;
            end
        end
      else
        begin
          reg216 = $unsigned(reg218);
        end
      if (reg125)
        begin
          reg226 = $unsigned((reg206[(5'h15):(4'hf)] ?
              ((reg220 >> $signed(reg195)) ?
                  ({reg165} ?
                      (reg218 ?
                          reg199 : reg221) : reg214) : (reg193[(4'hc):(1'h0)] ?
                      (reg172 ?
                          (8'ha7) : wire114) : (~&(8'ha1)))) : reg215[(2'h3):(2'h3)]));
          for (forvar227 = (1'h0); (forvar227 < (2'h3)); forvar227 = (forvar227 + (1'h1)))
            begin
              reg228 = reg153;
              reg229 <= wire114[(4'hb):(4'h9)];
              reg230 = (reg186 * reg170[(3'h4):(3'h4)]);
            end
        end
      else
        begin
          for (forvar226 = (1'h0); (forvar226 < (3'h4)); forvar226 = (forvar226 + (1'h1)))
            begin
              reg227 = $signed(reg206[(4'hb):(3'h6)]);
              reg229 <= (~&(($unsigned((reg218 + reg177)) != ((reg152 == reg228) ?
                  (reg152 ?
                      forvar226 : reg168) : (wire115 <<< reg214))) != wire111[(3'h4):(3'h4)]));
              reg230 = reg220[(4'ha):(3'h4)];
              reg231 = ($signed((~&$signed(reg215))) >= ($signed(reg223[(4'h8):(2'h3)]) ?
                  $signed({$unsigned((8'h9e))}) : {wire112}));
            end
        end
      reg232 <= (|wire110[(4'h9):(3'h5)]);
      for (forvar233 = (1'h0); (forvar233 < (1'h1)); forvar233 = (forvar233 + (1'h1)))
        begin
          reg234 = ((|reg148) ?
              $unsigned(((^~{reg177, reg177}) ?
                  ((reg138 * wire111) ?
                      (reg125 ?
                          reg151 : reg219) : (wire109 < reg226)) : wire111)) : forvar233);
          reg235 = $signed((~(^(-(+wire111)))));
          if (((reg223 ?
                  (reg125 ^ wire109[(1'h1):(1'h1)]) : $signed(reg208[(3'h4):(1'h0)])) ?
              ((~^((reg151 | reg189) ?
                  {reg189} : $unsigned(reg214))) << $unsigned(($unsigned(reg170) ?
                  (7'h48) : reg163))) : (7'h42)))
            begin
              reg236 <= reg172[(3'h7):(3'h6)];
            end
          else
            begin
              reg237 = ($signed(($signed({reg150}) >= reg199[(3'h7):(3'h6)])) ?
                  ($unsigned($signed((^~reg236))) <= {((reg221 > wire114) ?
                          reg220 : $unsigned(reg163)),
                      $signed(reg151)}) : $unsigned(reg176));
              reg238 = (~|$unsigned((&reg228)));
              reg239 <= $unsigned(forvar233[(4'hd):(4'h9)]);
              reg240 <= reg220;
            end
          reg241 = (&(7'h45));
          reg242 <= reg146;
        end
      reg243 <= forvar227[(3'h6):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg244 = reg199[(1'h0):(1'h0)];
      if ((7'h48))
        begin
          reg245 <= reg125;
          if (((((&reg154) ?
                  ($unsigned(reg171) ?
                      wire112 : $unsigned(reg171)) : reg223[(3'h5):(1'h1)]) ?
              $signed($signed($signed((8'hbe)))) : $signed($unsigned($unsigned((8'hb8))))) > ($signed((~|((8'ha5) << reg153))) ?
              $unsigned($signed(reg176[(5'h14):(4'hd)])) : $unsigned(reg177[(3'h6):(3'h6)]))))
            begin
              reg246 <= (reg171 >= reg206[(5'h10):(4'hd)]);
              reg247 <= (+(~$unsigned(reg146)));
              reg248 <= $unsigned(((reg189[(3'h5):(2'h2)] ?
                      (~^(reg152 <= reg117)) : {(reg150 ? reg188 : reg182)}) ?
                  reg126[(4'ha):(4'h9)] : (((!reg119) < (7'h48)) ?
                      ($signed(reg218) ?
                          reg117[(1'h1):(1'h0)] : (reg188 ?
                              (8'hb1) : reg170)) : ($signed(reg244) < reg206))));
              reg249 <= (&(($signed((wire114 ^~ (8'ha1))) ?
                  reg229[(4'ha):(2'h2)] : (reg153[(2'h2):(2'h2)] ?
                      (reg222 ?
                          reg126 : reg182) : reg195[(1'h0):(1'h0)])) ~^ ((+reg193[(2'h2):(2'h2)]) && (~|reg195[(1'h1):(1'h1)]))));
              reg250 <= reg193[(4'h8):(3'h5)];
            end
          else
            begin
              reg246 <= reg209;
              reg247 <= reg215[(1'h0):(1'h0)];
              reg251 = $unsigned(reg205);
            end
          reg252 <= reg193[(4'ha):(1'h0)];
          for (forvar253 = (1'h0); (forvar253 < (1'h1)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 = $signed(reg197);
              reg255 = (|reg131);
            end
          for (forvar256 = (1'h0); (forvar256 < (2'h3)); forvar256 = (forvar256 + (1'h1)))
            begin
              reg257 = (^~reg205);
              reg258 = $unsigned(reg150);
              reg259 <= $signed(reg151[(2'h2):(1'h1)]);
              reg260 <= ($unsigned(($unsigned({reg131}) || $unsigned((reg119 ?
                  reg164 : reg182)))) <= $unsigned(($signed(reg199[(2'h2):(2'h2)]) ?
                  $signed((reg232 != (8'hbe))) : reg224)));
              reg261 <= ($unsigned(reg214) ?
                  $signed(reg134[(3'h5):(2'h2)]) : reg135[(3'h7):(1'h1)]);
            end
        end
      else
        begin
          reg245 <= $signed(($signed($unsigned((reg176 ?
              reg131 : reg249))) <= $unsigned(reg164[(2'h2):(2'h2)])));
          reg251 = (~reg250);
          if ($signed(($signed(($unsigned(forvar253) ?
                  reg172 : (reg126 ? reg146 : reg215))) ?
              (reg223 ? $signed({reg252}) : reg150) : reg154)))
            begin
              reg252 <= reg172;
              reg253 = (|$unsigned(reg138[(2'h2):(1'h0)]));
              reg256 <= ($signed(reg188) ?
                  ((8'h9c) <= $unsigned({reg259[(1'h0):(1'h0)]})) : (-((&(reg254 ?
                      reg254 : (8'hb9))) - ($signed(reg219) != (reg224 ?
                      reg146 : reg118)))));
              reg259 <= (($signed(($signed(reg195) ?
                          wire113[(1'h1):(1'h0)] : (reg243 ?
                              reg154 : reg205))) ?
                      (reg261[(4'he):(3'h7)] == $unsigned((^~reg209))) : $unsigned($unsigned((reg178 ~^ reg153)))) ?
                  {reg260[(4'h9):(2'h2)],
                      ((|$signed((7'h4a))) == {forvar253[(5'h16):(3'h7)]})} : (|$signed($unsigned($unsigned(forvar256)))));
            end
          else
            begin
              reg252 <= $signed(({reg135[(4'hf):(4'he)]} == {(wire115 > $unsigned(reg150)),
                  ((forvar253 >= (8'ha3)) - (8'hb5))}));
              reg256 <= ((((+(7'h43)) != $signed($signed(reg232))) ?
                      ($signed((~^(8'ha4))) <<< $unsigned($unsigned(reg253))) : (reg201[(3'h7):(2'h3)] * reg174)) ?
                  $unsigned((&reg154)) : reg171);
              reg259 <= $signed($signed($unsigned($signed(reg176))));
              reg262 = ((8'hae) + (((+(!wire115)) ?
                  (reg250 ^~ (&reg152)) : reg206) != reg257[(2'h3):(1'h1)]));
            end
          reg263 <= (^~(!reg186));
          reg264 = reg186[(2'h2):(2'h2)];
        end
    end
  assign wire265 = (~($signed(($unsigned(reg247) < {reg252, reg186})) ?
                       reg193[(4'hb):(3'h7)] : (^reg164[(4'h9):(4'h9)])));
  always
    @(posedge clk) begin
      reg266 = ((&$unsigned(reg125)) || $unsigned(($signed((wire115 || reg247)) ?
          {reg178} : ({reg178, reg152} ? {reg260, reg177} : (~&reg193)))));
      reg267 <= $unsigned({(^~(~&reg163[(3'h5):(2'h2)]))});
      for (forvar268 = (1'h0); (forvar268 < (3'h4)); forvar268 = (forvar268 + (1'h1)))
        begin
          reg269 = $signed({(forvar268[(5'h10):(4'hd)] - (reg117[(4'hc):(1'h1)] ?
                  $signed(reg174) : reg189)),
              {(reg118[(3'h5):(1'h0)] ?
                      $signed(reg209) : reg250[(4'hf):(3'h5)]),
                  reg214}});
          reg270 <= reg266[(3'h5):(3'h4)];
          reg271 <= ((-reg270) && ((($signed(reg178) ^ reg163[(3'h5):(3'h4)]) ^ $signed($signed(reg245))) ?
              ($signed(reg163) ?
                  {(8'ha8)} : {(wire111 ?
                          reg182 : reg195)}) : $signed(reg263)));
        end
      for (forvar272 = (1'h0); (forvar272 < (1'h1)); forvar272 = (forvar272 + (1'h1)))
        begin
          reg273 <= (~^(&reg214[(5'h14):(3'h6)]));
          reg274 <= {(|reg154)};
        end
    end
  always
    @(posedge clk) begin
      if ((!(($signed((~&reg245)) ? reg245 : $signed(wire111)) ?
          (~^(^$signed(reg146))) : $signed({{(7'h43)}, {reg240}}))))
        begin
          if ((8'ha7))
            begin
              reg275 = (7'h47);
              reg276 <= reg186[(3'h5):(3'h5)];
            end
          else
            begin
              reg276 <= reg246;
              reg277 = (wire115 ?
                  (~^($signed(reg188[(1'h1):(1'h0)]) ?
                      $unsigned(reg168[(3'h6):(3'h4)]) : reg164[(2'h2):(1'h1)])) : {(^~$unsigned((reg153 ?
                          reg165 : reg223)))});
              reg278 = (~reg205[(1'h0):(1'h0)]);
            end
          reg279 <= (reg199 ?
              $unsigned((reg171 + ((wire112 ^ wire115) >> reg215[(3'h5):(3'h4)]))) : reg193[(4'he):(4'hb)]);
          if ($signed(reg197[(3'h7):(1'h0)]))
            begin
              reg280 = (wire111[(3'h6):(1'h0)] ?
                  $unsigned($signed($signed(reg246))) : $unsigned(($unsigned(reg261[(4'h8):(2'h2)]) ?
                      $signed(reg214[(5'h16):(5'h10)]) : reg125)));
              reg281 = $unsigned($signed((reg278 | $unsigned(wire115))));
            end
          else
            begin
              reg280 = (((((^~reg164) ?
                      (~(8'ha8)) : {reg245, wire265}) >= $signed((+(7'h44)))) ?
                  $signed(($signed(reg197) ?
                      $signed(reg263) : (^~reg136))) : wire111[(1'h0):(1'h0)]) ^ $signed(({wire115} & $unsigned(reg172[(4'hb):(3'h7)]))));
            end
        end
      else
        begin
          reg275 = $unsigned($unsigned((reg261[(3'h6):(3'h5)] ?
              {(reg182 ? reg245 : (7'h40))} : reg281)));
        end
      for (forvar282 = (1'h0); (forvar282 < (2'h2)); forvar282 = (forvar282 + (1'h1)))
        begin
          reg283 <= $signed((7'h41));
          reg284 = ((^~reg193[(1'h1):(1'h1)]) & (reg152 ?
              {{$unsigned(reg273), $unsigned((8'hb2))},
                  (reg223[(1'h0):(1'h0)] - (reg252 ?
                      reg205 : reg277))} : ($signed((|reg138)) <= $unsigned((reg245 ?
                  (8'ha4) : reg136)))));
        end
      reg285 = (+($signed(($unsigned(reg138) ?
          reg260[(4'hb):(1'h1)] : reg172[(1'h1):(1'h0)])) != {$signed((reg152 <<< (8'hb1))),
          $signed((&wire114))}));
      reg286 <= ($signed((reg276[(3'h4):(2'h3)] - ((reg224 - reg186) ?
          (reg182 & reg199) : $signed(reg277)))) != {$signed((~^(reg135 ^~ reg256)))});
      reg287 <= $signed(reg242);
    end
  always
    @(posedge clk) begin
      for (forvar288 = (1'h0); (forvar288 < (2'h2)); forvar288 = (forvar288 + (1'h1)))
        begin
          for (forvar289 = (1'h0); (forvar289 < (3'h4)); forvar289 = (forvar289 + (1'h1)))
            begin
              reg290 = reg174;
              reg291 <= {({(reg197 ? reg232 : reg215[(3'h4):(1'h0)]),
                      $signed(reg252)} >>> $unsigned($signed((~&wire265)))),
                  (reg174 < $signed($signed($unsigned(reg229))))};
              reg292 <= reg279[(1'h1):(1'h1)];
            end
          for (forvar293 = (1'h0); (forvar293 < (3'h4)); forvar293 = (forvar293 + (1'h1)))
            begin
              reg294 = reg126;
              reg295 <= (($unsigned($unsigned(reg294[(3'h4):(2'h3)])) | (8'haf)) ?
                  reg259[(2'h2):(1'h1)] : $unsigned($signed(reg219)));
              reg296 <= $unsigned($signed($unsigned({(reg256 ? reg208 : reg273),
                  reg208})));
            end
          reg297 = {reg283,
              (wire265[(1'h0):(1'h0)] && $unsigned(({reg224,
                  (7'h49)} * (reg232 > reg186))))};
        end
      for (forvar298 = (1'h0); (forvar298 < (1'h1)); forvar298 = (forvar298 + (1'h1)))
        begin
          reg299 <= {reg243, (^$unsigned((~^reg199)))};
          reg300 = reg163;
          if ((((($signed(reg206) ? {reg290} : forvar289) ?
                  (^~$unsigned(reg138)) : ((reg119 ? (7'h43) : (7'h42)) ?
                      $unsigned(reg259) : $signed((7'h45)))) ?
              (((reg205 & reg283) <= reg208[(1'h0):(1'h0)]) < ($unsigned(reg239) ?
                  ((8'ha6) ? reg172 : reg182) : (wire110 ?
                      reg299 : reg267))) : (8'ha4)) > (~^$signed((reg154[(3'h4):(2'h3)] ?
              reg248[(3'h6):(3'h4)] : $unsigned(reg270))))))
            begin
              reg301 = (|(&reg215));
              reg302 = (((8'h9f) && reg188[(4'h9):(1'h0)]) ?
                  {$unsigned(wire111), {$signed(reg232)}} : reg249);
              reg303 <= $unsigned((8'hbc));
            end
          else
            begin
              reg301 = {$unsigned(reg297[(5'h11):(1'h0)])};
              reg303 <= (&reg242);
              reg304 = ((((&(reg236 + reg205)) >> (+(reg292 ?
                      reg223 : (8'ha9)))) ?
                  (reg239[(2'h2):(2'h2)] ?
                      ((7'h48) >= $unsigned(reg222)) : $signed(reg236)) : ($signed({reg153}) ?
                      ($unsigned((8'ha7)) ?
                          {(8'hb0),
                              reg279} : reg295[(5'h15):(2'h3)]) : $signed(reg247))) <= (+$signed($unsigned((reg188 ?
                  reg188 : reg201)))));
              reg305 <= (~&$signed($signed($unsigned($signed(reg267)))));
            end
        end
    end
  assign wire306 = (reg150 & {($signed(((8'hb8) && reg242)) & (&reg131))});
  always
    @(posedge clk) begin
      reg307 <= {{(reg118[(1'h0):(1'h0)] ?
                  ((reg150 ?
                      reg243 : reg118) >> reg182[(4'h8):(4'h8)]) : (reg138[(2'h2):(1'h1)] ?
                      reg267[(3'h5):(2'h2)] : {(8'ha1)})),
              (-wire114)},
          ((reg214 ?
              reg174 : ((8'had) ?
                  wire306[(1'h0):(1'h0)] : $signed(reg138))) ^ (reg276[(1'h0):(1'h0)] ?
              reg242[(4'hb):(2'h2)] : {(reg299 ? reg240 : (8'hac))}))};
      if ({(~|$signed((-reg240)))})
        begin
          reg308 <= $signed((reg243[(4'h8):(3'h5)] | (((reg291 ?
                  wire115 : (8'hb8)) ~^ (wire111 > reg214)) ?
              wire113 : ((reg186 ?
                  reg270 : reg274) != reg256[(1'h0):(1'h0)]))));
          reg309 = (!($signed({wire265[(2'h3):(1'h1)], (~^reg296)}) ?
              ($unsigned(((7'h41) ? reg215 : reg174)) ?
                  $signed(reg271) : ((8'hbd) ?
                      reg214 : (reg186 ?
                          reg206 : reg243))) : (+((reg165 <= wire109) > reg249[(3'h6):(2'h2)]))));
        end
      else
        begin
          for (forvar308 = (1'h0); (forvar308 < (1'h0)); forvar308 = (forvar308 + (1'h1)))
            begin
              reg310 <= (~&reg174);
              reg311 <= $signed(reg308[(2'h2):(2'h2)]);
              reg312 <= $signed({$unsigned(($signed(reg286) || {(8'hbf)}))});
              reg313 <= (reg260 ?
                  $signed($signed(((reg119 ? (8'ha8) : reg189) ?
                      (reg126 ?
                          reg214 : reg250) : reg205[(2'h2):(2'h2)]))) : (reg276 ?
                      ($unsigned(reg263) * {(~&reg150)}) : $signed($signed((8'ha6)))));
            end
          reg314 <= reg136[(3'h6):(1'h0)];
          reg315 = {{($signed((~|reg206)) ^ reg199)},
              {reg291[(4'h8):(4'h8)],
                  ($unsigned((reg271 ? (8'hb3) : (8'hab))) ?
                      (7'h49) : {$unsigned(reg205), (^~reg296)})}};
          if (({reg240[(5'h10):(4'ha)]} != (^{((~reg260) >= reg168)})))
            begin
              reg316 = ({((~reg195) == $unsigned(((7'h48) ? reg174 : reg247))),
                  {{(^~reg189)}}} && reg308);
              reg317 <= $signed($unsigned(reg193[(2'h3):(2'h2)]));
              reg318 <= reg151[(2'h3):(2'h2)];
              reg319 = reg310;
              reg320 <= reg248;
            end
          else
            begin
              reg316 = ($unsigned({{(reg172 ? reg273 : reg248)}}) ?
                  reg182[(4'h8):(2'h3)] : $signed(((+(8'ha8)) > (&$signed(forvar308)))));
              reg319 = ((8'ha1) ^~ $unsigned((wire306[(3'h5):(2'h2)] ?
                  $unsigned($signed(reg188)) : (reg248[(3'h4):(1'h0)] <<< $unsigned((8'hb8))))));
              reg320 <= (~^reg291[(3'h7):(2'h2)]);
              reg321 <= $signed($signed(({{reg136, (7'h43)},
                      $unsigned(reg292)} ?
                  (~&reg260[(4'h8):(1'h0)]) : (8'ha2))));
              reg322 <= reg319;
            end
          reg323 <= reg164;
        end
      for (forvar324 = (1'h0); (forvar324 < (1'h0)); forvar324 = (forvar324 + (1'h1)))
        begin
          reg325 <= ($signed((((forvar308 ? reg170 : reg240) ~^ (reg247 ?
                  reg308 : reg312)) ~^ ((~&reg152) ?
                  (wire265 == reg152) : $unsigned(reg118)))) ?
              $signed(wire113[(1'h1):(1'h1)]) : reg267[(4'hc):(1'h1)]);
          for (forvar326 = (1'h0); (forvar326 < (1'h0)); forvar326 = (forvar326 + (1'h1)))
            begin
              reg327 = {$signed($signed($unsigned((7'h4a)))),
                  ({((reg152 ? (8'hae) : reg245) ?
                              (~^(8'hb6)) : $signed((8'ha4))),
                          {(&reg152), reg165}} ?
                      ((((8'hba) ^~ (8'haa)) ?
                              (reg236 ?
                                  wire265 : reg168) : (reg229 <= wire115)) ?
                          reg261 : {reg151[(1'h1):(1'h1)],
                              $unsigned(reg267)}) : ({(reg163 != reg118),
                          forvar326[(4'hf):(4'hd)]} ^ (reg246 ?
                          (~^reg224) : (reg296 != reg276))))};
              reg328 <= forvar324[(1'h0):(1'h0)];
              reg329 = (-$unsigned((8'hb8)));
            end
        end
      reg330 = $signed((^(((reg323 <= forvar326) >>> {(8'hb8)}) ^ $signed($unsigned((8'hb4))))));
    end
  always
    @(posedge clk) begin
      reg331 <= $unsigned($unsigned(reg270[(1'h1):(1'h0)]));
      reg332 <= (^(~&(^reg243)));
    end
  assign wire333 = $unsigned((reg286 >> reg313[(5'h16):(5'h15)]));
  assign wire334 = ((($signed(reg176[(1'h0):(1'h0)]) ?
                       $signed(reg119[(4'h9):(4'h8)]) : (^reg134)) > wire113) == (7'h40));
  always
    @(posedge clk) begin
      reg335 = $unsigned(reg131[(1'h1):(1'h0)]);
      reg336 <= reg165[(3'h5):(3'h5)];
      for (forvar337 = (1'h0); (forvar337 < (2'h3)); forvar337 = (forvar337 + (1'h1)))
        begin
          reg338 = $unsigned((-(|((~&wire114) ? reg214 : reg250))));
          reg339 = reg215[(2'h3):(1'h0)];
          reg340 <= $signed(((8'ha8) ?
              $unsigned(((^reg339) ?
                  $unsigned(reg229) : (reg308 ?
                      reg328 : reg186))) : $signed($signed(reg188))));
          for (forvar341 = (1'h0); (forvar341 < (3'h4)); forvar341 = (forvar341 + (1'h1)))
            begin
              reg342 = {reg178};
              reg343 <= reg314;
              reg344 = reg229[(1'h0):(1'h0)];
              reg345 = $unsigned($unsigned((reg172 ?
                  (wire115 ?
                      $unsigned(reg308) : ((8'hab) & (8'h9c))) : ((8'h9e) > ((7'h49) ?
                      reg169 : wire265)))));
            end
          reg346 = $signed($signed($signed(reg172)));
        end
      for (forvar347 = (1'h0); (forvar347 < (3'h4)); forvar347 = (forvar347 + (1'h1)))
        begin
          if ((!reg178[(3'h4):(1'h1)]))
            begin
              reg348 <= $signed($unsigned($signed((reg170[(1'h1):(1'h1)] ?
                  (|reg276) : (reg274 >> reg208)))));
              reg349 <= $signed(reg296[(4'ha):(2'h3)]);
              reg350 = (~^(($unsigned(reg340[(5'h14):(2'h2)]) ?
                  reg252 : (&reg332[(3'h6):(3'h4)])) - $signed($unsigned(reg247[(4'hc):(3'h5)]))));
              reg351 = $unsigned({$signed(reg318), $unsigned(reg188)});
            end
          else
            begin
              reg350 = (($unsigned(((reg296 ? reg247 : (8'hb2)) ?
                      $unsigned(reg263) : $signed(reg154))) <= $unsigned(reg332[(3'h4):(3'h4)])) ?
                  $unsigned((((reg249 * reg176) ?
                          reg135[(4'ha):(2'h3)] : $unsigned(reg219)) ?
                      ((reg346 ^ (8'hb5)) ?
                          $unsigned(reg125) : $unsigned(reg138)) : reg186[(5'h11):(4'he)])) : reg219[(1'h1):(1'h1)]);
              reg352 <= reg134;
              reg353 <= reg239[(1'h0):(1'h0)];
            end
          for (forvar354 = (1'h0); (forvar354 < (1'h0)); forvar354 = (forvar354 + (1'h1)))
            begin
              reg355 <= (($signed(($signed(reg322) ?
                          reg346[(3'h7):(3'h5)] : $unsigned(reg299))) ?
                      {$unsigned((8'hbb))} : reg295) ?
                  (^reg186) : $signed({reg224[(5'h12):(4'he)],
                      {(~&(8'hb3)), (forvar354 ? reg246 : (7'h48))}}));
              reg356 = reg174[(3'h6):(3'h4)];
              reg357 <= $signed((!(-(reg292 ? (|reg246) : $signed(reg177)))));
              reg358 = reg188;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar359 = (1'h0); (forvar359 < (3'h4)); forvar359 = (forvar359 + (1'h1)))
        begin
          if (reg193[(2'h3):(2'h3)])
            begin
              reg360 <= ($signed($unsigned(reg219[(1'h0):(1'h0)])) ?
                  (reg343 >> reg308) : $unsigned(reg340[(5'h17):(3'h6)]));
              reg361 = (($unsigned((&$unsigned(reg229))) ?
                      $signed(({reg134} << (reg243 || (8'hbd)))) : reg126[(4'ha):(2'h3)]) ?
                  (({{reg349, reg186}, reg224[(5'h10):(4'hd)]} ?
                      ($unsigned(reg271) == $signed(reg138)) : (|{reg360,
                          reg360})) <<< reg229[(4'hd):(3'h4)]) : reg171);
            end
          else
            begin
              reg361 = {reg270[(3'h4):(1'h1)], wire109};
              reg362 = reg246[(5'h12):(4'ha)];
              reg363 <= $signed((&(!reg320[(3'h6):(1'h0)])));
              reg364 = ((~{$signed($signed(reg295)),
                      ($unsigned(reg312) < $signed(reg348))}) ?
                  reg299 : reg246);
              reg365 = ($signed(((~^(reg151 ?
                  reg172 : reg348)) + (~$unsigned((8'h9d))))) ^ $signed(({(+reg224)} & (reg286 != $signed(reg247)))));
            end
          if (({reg250[(3'h6):(2'h2)],
              ((~^(reg240 << reg303)) ~^ $signed((!reg283)))} || (!reg165[(1'h0):(1'h0)])))
            begin
              reg366 <= reg363;
              reg367 = (+(&$unsigned({$unsigned((8'hb6))})));
              reg368 = reg349[(4'ha):(3'h4)];
            end
          else
            begin
              reg366 <= {$signed(reg172)};
              reg367 = (~|(-(&reg357)));
              reg368 = reg368;
            end
          if (reg125)
            begin
              reg369 = ((reg332[(2'h2):(1'h0)] ?
                      $unsigned($unsigned($signed(reg363))) : reg135[(4'hf):(4'ha)]) ?
                  ({$unsigned($signed(reg150)), reg299} ?
                      $signed(reg224[(3'h4):(3'h4)]) : $unsigned($signed((~|reg151)))) : $unsigned(({(|(8'hb8))} << $signed((8'hbb)))));
              reg370 <= ($signed(((~$signed(reg369)) ^ (((8'hbb) - reg332) ~^ ((7'h41) == reg343)))) ?
                  $signed((8'h9c)) : reg310[(3'h4):(1'h0)]);
            end
          else
            begin
              reg369 = $signed($signed(({reg349} != $signed(reg310))));
            end
          reg371 = $unsigned((|(+reg154[(2'h3):(2'h3)])));
        end
      for (forvar372 = (1'h0); (forvar372 < (2'h2)); forvar372 = (forvar372 + (1'h1)))
        begin
          reg373 <= reg219[(2'h2):(1'h0)];
          if ($signed(wire333))
            begin
              reg374 <= ((!((+(-reg308)) >= reg328[(1'h1):(1'h1)])) ^~ reg363);
              reg375 <= reg299;
              reg376 = (|wire333[(3'h6):(1'h0)]);
            end
          else
            begin
              reg376 = reg366;
            end
          for (forvar377 = (1'h0); (forvar377 < (2'h3)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg378 = (|(~&reg171));
              reg379 <= $signed($unsigned($signed((+$signed((7'h48))))));
            end
          reg380 = {reg271};
        end
    end
  always
    @(posedge clk) begin
      reg381 <= (-((($signed((7'h49)) ?
              reg243[(4'hc):(2'h2)] : ((8'hb7) + reg366)) | $unsigned((|reg146))) ?
          reg260[(4'h9):(4'h8)] : reg209));
      reg382 = (~&$unsigned(((reg321 ? reg320 : (reg249 ? reg370 : (8'ha7))) ?
          $unsigned(((8'hb2) != reg270)) : ((^~reg119) ?
              {reg307} : $unsigned((8'hb8))))));
      if ((^~$signed((!((wire111 ~^ reg381) ?
          ((8'h9e) || reg287) : (reg151 ? reg321 : reg154))))))
        begin
          reg383 = reg229;
        end
      else
        begin
          if (reg125[(4'hc):(1'h1)])
            begin
              reg384 <= ($unsigned(reg219) - $signed($signed(reg283)));
              reg385 = ((7'h44) || ($signed(reg222[(3'h6):(3'h6)]) ?
                  ($signed((reg256 ?
                      reg370 : reg174)) ^ $unsigned($signed(reg349))) : $signed(({reg274,
                          reg313} ?
                      (reg134 ? reg171 : (8'hac)) : reg375[(2'h3):(1'h0)]))));
            end
          else
            begin
              reg384 <= (|reg154);
              reg386 <= $unsigned(reg118);
            end
          reg387 = $signed(((-$unsigned((~reg296))) * $unsigned((~(reg353 ?
              reg311 : wire333)))));
          reg388 <= ((-reg263[(5'h16):(4'ha)]) << (reg224 ? (7'h42) : reg323));
        end
      reg389 <= ($unsigned(reg340) <<< $unsigned(reg311));
      for (forvar390 = (1'h0); (forvar390 < (1'h1)); forvar390 = (forvar390 + (1'h1)))
        begin
          for (forvar391 = (1'h0); (forvar391 < (1'h0)); forvar391 = (forvar391 + (1'h1)))
            begin
              reg392 = (({((reg321 ? reg214 : reg165) ?
                          reg259[(4'h8):(1'h1)] : wire115[(5'h10):(4'he)])} < $unsigned(reg296[(4'hc):(2'h3)])) ?
                  (|$signed(((reg305 ? reg307 : wire334) ~^ {(8'ha4),
                      (7'h42)}))) : $signed($unsigned((reg325 ?
                      reg317 : (reg312 ? reg169 : reg215)))));
              reg393 = (-(&(reg206[(3'h5):(3'h4)] > (8'h9f))));
              reg394 <= ((($unsigned((8'ha3)) >= $unsigned((reg271 ?
                  reg182 : reg186))) - $unsigned($signed((^~reg118)))) >>> $unsigned(reg248[(1'h1):(1'h1)]));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar395 = (1'h0); (forvar395 < (2'h3)); forvar395 = (forvar395 + (1'h1)))
        begin
          reg396 <= $signed((-(((!reg322) > (reg343 ? reg186 : (7'h42))) ?
              reg239 : {$unsigned(reg195)})));
          for (forvar397 = (1'h0); (forvar397 < (3'h4)); forvar397 = (forvar397 + (1'h1)))
            begin
              reg398 <= reg119[(4'hc):(4'h9)];
              reg399 <= (reg169 ?
                  {$signed(reg239)} : {reg189[(3'h4):(2'h2)],
                      (reg261[(4'hf):(4'ha)] ?
                          (!(reg224 == reg224)) : reg215)});
            end
          reg400 = {reg152, $unsigned($signed($signed((&reg247))))};
          reg401 <= reg153[(1'h0):(1'h0)];
          reg402 <= $unsigned(reg379);
        end
      if ((~|$signed(reg232[(1'h1):(1'h1)])))
        begin
          if ((reg150[(3'h5):(1'h1)] == reg176))
            begin
              reg403 <= $unsigned($unsigned(({wire112,
                      ((8'ha0) ? reg239 : reg214)} ?
                  $unsigned(reg401[(4'h9):(4'h9)]) : reg153)));
              reg404 = (8'h9d);
              reg405 <= $signed(reg125);
            end
          else
            begin
              reg404 = reg214[(3'h4):(3'h4)];
            end
          reg406 = {{(reg310[(4'hc):(3'h7)] ?
                      {(reg163 * reg164)} : reg222[(4'hf):(1'h1)])}};
          for (forvar407 = (1'h0); (forvar407 < (2'h2)); forvar407 = (forvar407 + (1'h1)))
            begin
              reg408 = ({(8'ha4)} * (($unsigned(reg276[(1'h1):(1'h1)]) ?
                      ((reg215 ?
                          reg188 : reg138) ~^ $unsigned(reg245)) : $signed(wire265[(3'h7):(1'h0)])) ?
                  ($unsigned(forvar395) ?
                      reg177 : reg152[(5'h14):(4'hf)]) : (~|$unsigned((^wire333)))));
              reg409 <= $signed(wire333);
              reg410 = (~^({$unsigned($signed(reg355))} ?
                  (~|(8'hab)) : {$unsigned((reg399 ? reg343 : reg178))}));
            end
        end
      else
        begin
          for (forvar403 = (1'h0); (forvar403 < (3'h4)); forvar403 = (forvar403 + (1'h1)))
            begin
              reg405 <= (7'h45);
              reg407 <= $unsigned($signed($signed(({reg197} ?
                  reg243[(3'h5):(3'h5)] : $unsigned(reg177)))));
              reg408 = (^reg153[(1'h0):(1'h0)]);
              reg409 <= $unsigned(reg307[(3'h4):(1'h1)]);
              reg410 = (reg125[(1'h1):(1'h0)] ?
                  (^wire265[(3'h4):(3'h4)]) : $signed((^({(8'hb4)} ?
                      {(7'h49)} : ((7'h49) ? (7'h49) : reg195)))));
            end
          if ((~|reg388[(3'h4):(1'h0)]))
            begin
              reg411 = $unsigned({reg394[(1'h0):(1'h0)]});
            end
          else
            begin
              reg411 = ((&(((8'ha4) >>> {reg307}) != $signed((+wire109)))) ?
                  (reg134[(4'hf):(4'ha)] ?
                      (!reg232) : ($unsigned($signed(reg239)) * reg252)) : {reg208[(1'h0):(1'h0)],
                      $unsigned({reg401})});
              reg412 = $unsigned(reg177);
              reg413 = reg168[(2'h2):(2'h2)];
              reg414 <= $unsigned(reg352[(4'hf):(4'ha)]);
            end
          if ($signed(((&$signed($signed(reg295))) ?
              {({reg229, (8'ha0)} ?
                      (reg313 ? (8'hbe) : reg171) : (reg209 ? reg165 : reg399)),
                  (|$unsigned(reg402))} : $unsigned(((reg394 > reg349) < (-reg394))))))
            begin
              reg415 <= ($signed((~^((wire109 * (8'hbd)) || (reg295 ?
                      (8'haa) : reg406)))) ?
                  (~&$unsigned((((8'ha1) ? reg170 : reg263) ?
                      reg404[(3'h7):(2'h3)] : ((8'ha5) >>> reg178)))) : reg409);
              reg416 <= (reg396 ?
                  (!((8'hb8) ?
                      $signed($unsigned(wire115)) : $unsigned(reg224[(4'hb):(4'h8)]))) : reg374[(3'h5):(2'h2)]);
              reg417 <= (!(8'hb2));
              reg418 <= reg386;
              reg419 = ((7'h4a) ?
                  (reg125 >> ((~|(reg352 ? reg328 : forvar403)) ?
                      reg310 : $unsigned(reg296))) : (^~$signed({wire114[(3'h5):(1'h0)]})));
            end
          else
            begin
              reg415 <= (^(reg307[(3'h6):(1'h1)] ?
                  (^$signed($signed(reg154))) : (((reg401 >> reg270) && $signed(reg413)) ?
                      reg274[(3'h7):(2'h2)] : (~&(8'hac)))));
              reg419 = (+reg218[(2'h2):(2'h2)]);
            end
          reg420 = wire111[(1'h1):(1'h1)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1527  (y, clk, wire1531, wire1530, wire1529, wire1528);
  output wire [(32'h47e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire1531;
  input wire [(3'h6):(1'h0)] wire1530;
  input wire signed [(4'h9):(1'h0)] wire1529;
  input wire signed [(5'h12):(1'h0)] wire1528;
  wire [(5'h17):(1'h0)] wire1616;
  wire signed [(2'h3):(1'h0)] wire1601;
  wire signed [(2'h2):(1'h0)] wire1600;
  wire [(5'h13):(1'h0)] wire1532;
  reg signed [(3'h6):(1'h0)] reg1615 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1612 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1611 = (1'h0);
  reg [(2'h3):(1'h0)] reg1610 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1608 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1606 = (1'h0);
  reg [(4'h8):(1'h0)] reg1604 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1598 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1594 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1591 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1588 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1587 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1585 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1578 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1582 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1581 = (1'h0);
  reg [(3'h7):(1'h0)] reg1577 = (1'h0);
  reg [(5'h12):(1'h0)] reg1575 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1574 = (1'h0);
  reg [(5'h14):(1'h0)] reg1573 = (1'h0);
  reg [(4'hc):(1'h0)] reg1571 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1569 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1568 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1567 = (1'h0);
  reg [(2'h3):(1'h0)] reg1566 = (1'h0);
  reg [(5'h12):(1'h0)] reg1563 = (1'h0);
  reg [(3'h6):(1'h0)] reg1562 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1559 = (1'h0);
  reg [(3'h5):(1'h0)] reg1557 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1555 = (1'h0);
  reg [(3'h4):(1'h0)] reg1554 = (1'h0);
  reg [(3'h4):(1'h0)] reg1553 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1552 = (1'h0);
  reg [(4'hf):(1'h0)] reg1549 = (1'h0);
  reg [(4'hb):(1'h0)] reg1548 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1546 = (1'h0);
  reg [(4'h9):(1'h0)] reg1545 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1543 = (1'h0);
  reg [(3'h5):(1'h0)] reg1540 = (1'h0);
  reg [(2'h3):(1'h0)] reg1539 = (1'h0);
  reg [(5'h10):(1'h0)] reg1538 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1537 = (1'h0);
  reg [(5'h17):(1'h0)] reg1534 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1609 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1614 = (1'h0);
  reg [(5'h14):(1'h0)] reg1613 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1609 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1607 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1605 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1603 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1602 = (1'h0);
  reg [(4'hc):(1'h0)] reg1599 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1597 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1596 = (1'h0);
  reg [(5'h16):(1'h0)] reg1595 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1593 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1590 = (1'h0);
  reg [(5'h17):(1'h0)] reg1589 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1586 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1584 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1583 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1577 = (1'h0);
  reg [(4'ha):(1'h0)] reg1580 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1579 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1578 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1576 = (1'h0);
  reg [(4'h9):(1'h0)] reg1572 = (1'h0);
  reg [(3'h4):(1'h0)] reg1570 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1569 = (1'h0);
  reg [(4'hf):(1'h0)] reg1565 = (1'h0);
  reg [(4'hc):(1'h0)] reg1564 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1561 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1560 = (1'h0);
  reg [(2'h2):(1'h0)] reg1556 = (1'h0);
  reg [(5'h12):(1'h0)] reg1558 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1556 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1551 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1550 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1541 = (1'h0);
  reg [(5'h14):(1'h0)] reg1535 = (1'h0);
  reg [(3'h6):(1'h0)] reg1533 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1547 = (1'h0);
  reg [(4'hf):(1'h0)] reg1544 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1542 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1541 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1536 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1535 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1533 = (1'h0);
  assign y = {wire1616,
                 wire1601,
                 wire1600,
                 wire1532,
                 reg1615,
                 reg1612,
                 reg1611,
                 reg1610,
                 reg1608,
                 reg1606,
                 reg1604,
                 reg1598,
                 reg1594,
                 reg1591,
                 reg1588,
                 reg1587,
                 reg1585,
                 reg1578,
                 reg1582,
                 reg1581,
                 reg1577,
                 reg1575,
                 reg1574,
                 reg1573,
                 reg1571,
                 reg1569,
                 reg1568,
                 reg1567,
                 reg1566,
                 reg1563,
                 reg1562,
                 reg1559,
                 reg1557,
                 reg1555,
                 reg1554,
                 reg1553,
                 reg1552,
                 reg1549,
                 reg1548,
                 reg1546,
                 reg1545,
                 reg1543,
                 reg1540,
                 reg1539,
                 reg1538,
                 reg1537,
                 reg1534,
                 reg1609,
                 reg1614,
                 reg1613,
                 forvar1609,
                 reg1607,
                 reg1605,
                 reg1603,
                 reg1602,
                 reg1599,
                 reg1597,
                 forvar1596,
                 reg1595,
                 reg1593,
                 reg1592,
                 forvar1590,
                 reg1589,
                 reg1586,
                 reg1584,
                 reg1583,
                 forvar1577,
                 reg1580,
                 reg1579,
                 forvar1578,
                 reg1576,
                 reg1572,
                 reg1570,
                 forvar1569,
                 reg1565,
                 reg1564,
                 forvar1561,
                 reg1560,
                 reg1556,
                 reg1558,
                 forvar1556,
                 forvar1551,
                 reg1550,
                 reg1541,
                 reg1535,
                 reg1533,
                 reg1547,
                 reg1544,
                 reg1542,
                 forvar1541,
                 reg1536,
                 forvar1535,
                 forvar1533,
                 (1'h0)};
  assign wire1532 = (wire1529[(1'h0):(1'h0)] ?
                        (({(wire1530 ?
                                wire1528 : wire1528)} | {(wire1528 - wire1531)}) - $unsigned(((^(8'hb3)) ?
                            wire1530 : (wire1531 << wire1530)))) : ({(&wire1531[(5'h12):(4'ha)]),
                                $signed(wire1531[(5'h10):(4'h8)])} ?
                            (~(8'hb8)) : (&((!wire1529) << (7'h46)))));
  always
    @(posedge clk) begin
      if ((-wire1530))
        begin
          for (forvar1533 = (1'h0); (forvar1533 < (2'h3)); forvar1533 = (forvar1533 + (1'h1)))
            begin
              reg1534 <= $unsigned($unsigned(wire1528[(4'ha):(4'h9)]));
            end
          for (forvar1535 = (1'h0); (forvar1535 < (2'h2)); forvar1535 = (forvar1535 + (1'h1)))
            begin
              reg1536 = $unsigned(wire1531[(4'he):(4'hd)]);
              reg1537 <= ($signed($unsigned(({wire1531,
                  wire1532} ~^ (&forvar1535)))) >> $signed(wire1528));
              reg1538 <= (+(&$unsigned({reg1537})));
              reg1539 <= reg1536;
              reg1540 <= $unsigned(($signed($unsigned(reg1537[(2'h3):(2'h2)])) ~^ $signed(wire1531)));
            end
          for (forvar1541 = (1'h0); (forvar1541 < (1'h0)); forvar1541 = (forvar1541 + (1'h1)))
            begin
              reg1542 = $signed($signed(wire1530[(3'h5):(2'h3)]));
              reg1543 <= wire1530[(3'h5):(3'h4)];
              reg1544 = $unsigned($signed((^~(((7'h41) >>> forvar1535) - (reg1543 >>> wire1528)))));
              reg1545 <= (reg1539[(2'h3):(2'h3)] + (($unsigned((reg1542 << reg1539)) ?
                      ((~|reg1534) > reg1536[(3'h7):(3'h5)]) : wire1531[(4'hf):(3'h4)]) ?
                  reg1544[(2'h3):(2'h3)] : $signed(((7'h46) ?
                      {reg1539} : (wire1529 <= reg1538)))));
            end
          if ($unsigned($unsigned((-((wire1530 >= reg1542) ^ $signed(reg1544))))))
            begin
              reg1546 <= (reg1543[(2'h2):(1'h0)] & (7'h49));
              reg1547 = (^(~^((+$signed(reg1534)) ?
                  $signed(reg1542) : (~^$unsigned(reg1538)))));
              reg1548 <= $signed((reg1537 ^ $unsigned((&reg1536[(1'h0):(1'h0)]))));
              reg1549 <= reg1543;
            end
          else
            begin
              reg1546 <= wire1530[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg1533 = $signed(wire1530);
          if (($unsigned($unsigned(wire1532)) ~^ reg1544[(4'h9):(1'h0)]))
            begin
              reg1535 = wire1530;
              reg1536 = {((reg1540 && wire1530[(1'h1):(1'h0)]) ?
                      (~^(^(&reg1542))) : $unsigned({reg1537}))};
              reg1537 <= ($unsigned((-reg1539[(1'h1):(1'h1)])) >> (!(reg1548[(4'h9):(2'h3)] ?
                  ((~reg1548) || ((7'h46) > wire1531)) : ($signed(reg1536) ?
                      reg1535[(5'h12):(2'h2)] : $unsigned(reg1533)))));
              reg1538 <= $unsigned((($signed($signed(reg1548)) ?
                      $signed(reg1533[(1'h0):(1'h0)]) : ($unsigned(wire1532) & $unsigned(reg1543))) ?
                  (~^reg1539[(1'h0):(1'h0)]) : $signed(wire1531[(1'h0):(1'h0)])));
              reg1539 <= $signed((~^(((reg1533 <<< forvar1533) ?
                      (7'h45) : (wire1528 ~^ wire1528)) ?
                  $signed({reg1537, reg1539}) : $unsigned(reg1549))));
            end
          else
            begin
              reg1535 = (^wire1528);
              reg1536 = {({$signed(reg1543[(1'h1):(1'h0)])} == $unsigned((^{reg1543,
                      reg1534}))),
                  $signed({(^$unsigned((8'hbc))), reg1547})};
              reg1541 = {(wire1531 <<< (8'hb4))};
            end
        end
      if (($unsigned($signed(reg1538[(2'h3):(1'h1)])) && $unsigned($unsigned(((~reg1534) ?
          $unsigned(reg1536) : forvar1535)))))
        begin
          reg1550 = (~|reg1547[(4'ha):(1'h1)]);
          for (forvar1551 = (1'h0); (forvar1551 < (2'h3)); forvar1551 = (forvar1551 + (1'h1)))
            begin
              reg1552 <= reg1533[(1'h1):(1'h0)];
              reg1553 <= reg1544[(4'he):(4'h9)];
              reg1554 <= $unsigned($signed((forvar1533 >> (reg1541[(3'h6):(2'h3)] ?
                  $signed(reg1546) : $signed((7'h45))))));
              reg1555 <= ((((&(wire1531 ? reg1543 : forvar1541)) ?
                      reg1545 : (8'ha6)) ?
                  forvar1551 : (!reg1545[(1'h1):(1'h0)])) - reg1549);
            end
          for (forvar1556 = (1'h0); (forvar1556 < (2'h2)); forvar1556 = (forvar1556 + (1'h1)))
            begin
              reg1557 <= $signed(reg1533[(2'h3):(1'h0)]);
              reg1558 = (&reg1545[(1'h1):(1'h1)]);
              reg1559 <= $unsigned(reg1533[(3'h4):(1'h1)]);
            end
        end
      else
        begin
          reg1550 = forvar1535;
          for (forvar1551 = (1'h0); (forvar1551 < (3'h4)); forvar1551 = (forvar1551 + (1'h1)))
            begin
              reg1556 = (~|$signed((^$signed({reg1552}))));
              reg1558 = ($unsigned(($unsigned($signed(reg1539)) ?
                      {(reg1548 != forvar1551)} : (~^reg1536))) ?
                  $unsigned(($unsigned($unsigned(forvar1556)) >> ((!reg1547) == ((8'h9e) * (7'h43))))) : $unsigned($signed(reg1538[(3'h7):(3'h7)])));
            end
          reg1560 = ({(|$signed(reg1554)),
                  ($signed((8'hba)) ?
                      reg1549 : ((wire1528 != reg1550) & reg1539[(1'h0):(1'h0)]))} ?
              reg1537 : $unsigned(($unsigned($signed(forvar1541)) ?
                  forvar1556[(2'h2):(1'h1)] : reg1544[(1'h1):(1'h1)])));
          for (forvar1561 = (1'h0); (forvar1561 < (1'h1)); forvar1561 = (forvar1561 + (1'h1)))
            begin
              reg1562 <= {(reg1560[(3'h7):(2'h3)] >>> (+{(^(7'h46)),
                      (reg1536 ? (8'hbd) : (8'h9d))}))};
              reg1563 <= (reg1549 | (reg1542 >>> (~|{(wire1530 ?
                      reg1562 : forvar1556),
                  {forvar1535}})));
              reg1564 = $unsigned((reg1535[(4'hf):(3'h6)] ?
                  (~|($signed(reg1546) < $unsigned(wire1528))) : (~|(~|{reg1563}))));
              reg1565 = reg1550;
            end
        end
      reg1566 <= reg1554;
      reg1567 <= ((~|reg1537) ?
          (reg1555[(4'h8):(1'h0)] ?
              (7'h40) : wire1532[(3'h7):(2'h2)]) : ($unsigned(reg1555) | $unsigned((forvar1556[(2'h2):(2'h2)] < $signed(reg1543)))));
      reg1568 <= reg1560[(3'h6):(3'h6)];
    end
  always
    @(posedge clk) begin
      if ((^{(($signed(wire1532) && $unsigned(reg1539)) ^ $signed(wire1531[(3'h7):(2'h3)])),
          reg1566}))
        begin
          reg1569 <= reg1546[(4'hf):(4'hc)];
        end
      else
        begin
          for (forvar1569 = (1'h0); (forvar1569 < (3'h4)); forvar1569 = (forvar1569 + (1'h1)))
            begin
              reg1570 = $signed(($unsigned((reg1559 && reg1548)) ?
                  reg1537 : ({(forvar1569 ? reg1557 : reg1568),
                      reg1545[(4'h9):(2'h2)]} <= {(reg1552 ~^ reg1569)})));
              reg1571 <= (reg1562 ?
                  $unsigned(({(~&forvar1569), {reg1548}} ?
                      (-$signed((8'hb7))) : (-((8'hbd) >= reg1567)))) : ({$signed((!reg1568))} ?
                      (8'hb2) : ($signed(reg1570[(3'h4):(1'h1)]) ^ $signed((reg1562 ?
                          wire1530 : reg1549)))));
              reg1572 = $signed($signed(reg1570[(1'h0):(1'h0)]));
              reg1573 <= forvar1569[(2'h2):(2'h2)];
              reg1574 <= $signed((reg1570[(1'h0):(1'h0)] ?
                  (reg1552 || ((reg1538 | wire1531) ?
                      (wire1529 & reg1534) : (8'hb2))) : ({(reg1539 == wire1529)} == $unsigned((~reg1555)))));
            end
          reg1575 <= reg1574;
          reg1576 = $unsigned(($unsigned($unsigned(reg1573)) == (((~(8'hb1)) ?
              $unsigned(reg1559) : reg1563[(4'ha):(1'h1)]) <= $unsigned($signed(reg1554)))));
        end
      if ((~&$unsigned($unsigned($signed({forvar1569})))))
        begin
          reg1577 <= (wire1532 ?
              reg1559[(3'h4):(1'h1)] : (&((reg1546 ? (~reg1540) : {reg1563}) ?
                  ((reg1573 >>> reg1554) ?
                      $signed(wire1528) : $signed(reg1569)) : $unsigned(reg1563[(4'h8):(2'h3)]))));
          for (forvar1578 = (1'h0); (forvar1578 < (1'h0)); forvar1578 = (forvar1578 + (1'h1)))
            begin
              reg1579 = ($signed($unsigned($unsigned(reg1567))) ?
                  (reg1562 <= reg1555[(2'h2):(2'h2)]) : $unsigned(reg1567));
              reg1580 = {$signed($unsigned((reg1579[(4'h9):(3'h4)] ?
                      (+(8'hb2)) : (8'ha2))))};
              reg1581 <= (!reg1537[(1'h1):(1'h0)]);
              reg1582 <= $signed($signed($signed((^~(forvar1578 ?
                  forvar1569 : reg1553)))));
            end
        end
      else
        begin
          for (forvar1577 = (1'h0); (forvar1577 < (3'h4)); forvar1577 = (forvar1577 + (1'h1)))
            begin
              reg1578 <= reg1581[(5'h11):(4'hf)];
              reg1579 = (reg1580 ?
                  $signed(((reg1559[(2'h3):(2'h3)] ?
                      (+reg1576) : $unsigned(reg1549)) | {{reg1571,
                          reg1563}})) : reg1575[(3'h7):(2'h3)]);
            end
          reg1580 = reg1580;
          reg1581 <= ($unsigned(reg1575[(1'h0):(1'h0)]) || $signed(reg1578));
        end
      if ($unsigned(({({reg1570} && reg1538)} ?
          wire1531[(5'h12):(2'h3)] : (8'ha1))))
        begin
          reg1583 = (reg1570[(2'h3):(2'h2)] != (^reg1562));
          if ({(-($unsigned(((7'h41) && (7'h40))) ?
                  (8'hae) : reg1545[(1'h1):(1'h0)])),
              reg1540[(3'h4):(2'h3)]})
            begin
              reg1584 = forvar1578;
              reg1585 <= $signed(($unsigned(reg1552[(5'h11):(2'h2)]) >= ($unsigned(((7'h46) ?
                  reg1572 : reg1582)) ^ ((reg1584 ? reg1557 : reg1543) ?
                  reg1538[(1'h1):(1'h0)] : (reg1569 != reg1555)))));
            end
          else
            begin
              reg1584 = (($unsigned((~^(reg1570 ?
                  wire1532 : reg1574))) + $unsigned($unsigned({reg1571}))) >= (^$signed(reg1546[(4'hf):(1'h1)])));
              reg1586 = (!$unsigned(forvar1577[(5'h15):(1'h0)]));
              reg1587 <= reg1562;
              reg1588 <= $signed($signed(reg1579));
              reg1589 = $unsigned(reg1586[(4'hd):(4'hc)]);
            end
          for (forvar1590 = (1'h0); (forvar1590 < (2'h2)); forvar1590 = (forvar1590 + (1'h1)))
            begin
              reg1591 <= reg1562[(3'h6):(2'h2)];
              reg1592 = reg1534[(5'h12):(3'h5)];
              reg1593 = ($unsigned(wire1529[(3'h4):(2'h3)]) ?
                  $signed(($unsigned((reg1591 >>> (8'h9f))) ?
                      (wire1531 ?
                          reg1570 : (reg1571 ^~ reg1549)) : $signed((reg1557 ?
                          reg1571 : reg1576)))) : (reg1569[(4'h8):(1'h0)] >> $unsigned(({reg1582} << $signed(reg1557)))));
              reg1594 <= {((reg1554 || $unsigned($unsigned(reg1592))) > ((&reg1555[(3'h5):(2'h2)]) ?
                      {$unsigned(wire1528),
                          $signed(reg1578)} : (reg1539[(1'h0):(1'h0)] ?
                          $unsigned((7'h49)) : (reg1568 <= reg1585))))};
            end
          reg1595 = $unsigned(reg1586);
          for (forvar1596 = (1'h0); (forvar1596 < (1'h0)); forvar1596 = (forvar1596 + (1'h1)))
            begin
              reg1597 = (^(^(forvar1577 + ({reg1534, reg1534} ?
                  $unsigned((8'hbe)) : reg1576))));
            end
        end
      else
        begin
          if ($unsigned((((~$unsigned((8'had))) ?
              ((reg1593 ? (8'ha5) : reg1582) != ((8'hab) ?
                  reg1588 : forvar1578)) : reg1588[(4'h9):(1'h1)]) >> (-(-{reg1585,
              reg1540})))))
            begin
              reg1583 = {(~^reg1539[(2'h2):(1'h0)])};
              reg1584 = $unsigned($signed(reg1549[(4'hb):(3'h4)]));
              reg1585 <= $unsigned(reg1538[(1'h0):(1'h0)]);
              reg1586 = reg1589;
              reg1587 <= (-(reg1557 ?
                  reg1597[(2'h3):(2'h2)] : ((reg1588 ?
                      reg1591 : {reg1553,
                          reg1585}) || $signed($signed(reg1563)))));
            end
          else
            begin
              reg1583 = $unsigned($unsigned($signed($unsigned(forvar1577[(2'h2):(1'h1)]))));
              reg1584 = $signed($unsigned(wire1529[(3'h5):(1'h0)]));
              reg1586 = (+$unsigned(reg1582));
              reg1587 <= ({((~|(wire1532 ? reg1567 : reg1553)) ?
                          reg1588 : (~reg1545[(3'h7):(2'h3)])),
                      $signed(((|reg1548) ? $signed(reg1591) : wire1531))} ?
                  ($unsigned($signed((reg1580 ? reg1585 : (8'hbf)))) ?
                      $signed(((reg1570 ? reg1539 : reg1578) ?
                          reg1587[(2'h3):(2'h2)] : $unsigned(reg1538))) : (reg1568 == ($unsigned(reg1553) ?
                          forvar1596 : {reg1594,
                              (7'h49)}))) : reg1554[(2'h3):(1'h0)]);
              reg1588 <= ((8'ha6) << (^~reg1577[(3'h6):(3'h4)]));
            end
        end
      reg1598 <= {$unsigned($unsigned($unsigned(reg1552))),
          {(^~(~^(~(8'h9d)))), reg1573[(3'h4):(1'h0)]}};
      reg1599 = (|((-(~reg1539[(1'h0):(1'h0)])) <<< {(~|$unsigned(reg1549)),
          (~|{reg1593, (8'hb0)})}));
    end
  assign wire1600 = (($signed($unsigned(reg1585[(4'hf):(4'hf)])) >>> reg1537[(1'h1):(1'h1)]) || (-(~&reg1568[(5'h17):(4'hc)])));
  assign wire1601 = reg1566;
  always
    @(posedge clk) begin
      reg1602 = (+$signed(reg1566));
      if (reg1540)
        begin
          if ((($signed($signed((^~reg1540))) > {reg1539[(1'h1):(1'h0)],
              $signed((reg1553 ? wire1531 : reg1552))}) - $unsigned((reg1554 ?
              (wire1532[(2'h2):(1'h0)] ?
                  $signed(reg1598) : (^wire1601)) : reg1540))))
            begin
              reg1603 = ($signed(reg1552[(1'h1):(1'h0)]) ?
                  $unsigned(reg1587[(1'h1):(1'h1)]) : (((+$unsigned(wire1529)) ^ $unsigned(wire1601[(1'h1):(1'h1)])) >> (!wire1529[(4'h8):(3'h6)])));
              reg1604 <= (~&(~^$unsigned((-$signed(reg1552)))));
              reg1605 = ((+$unsigned(((^reg1581) ^ $signed(reg1538)))) ?
                  (reg1571[(4'ha):(3'h6)] + (~|$signed((+reg1581)))) : ($unsigned({(wire1531 - reg1554)}) ?
                      reg1548 : ($signed((reg1540 > reg1582)) <<< ($signed((8'hbe)) | {reg1540,
                          wire1532}))));
              reg1606 <= $unsigned($signed((|$unsigned(reg1578[(2'h2):(1'h0)]))));
              reg1607 = $unsigned($signed((8'hbb)));
            end
          else
            begin
              reg1604 <= ((~^reg1548[(2'h2):(1'h0)]) > $unsigned((~|(reg1569 ?
                  (~reg1594) : reg1554[(1'h0):(1'h0)]))));
              reg1605 = wire1600[(1'h0):(1'h0)];
              reg1606 <= reg1594;
              reg1608 <= $unsigned(reg1545[(3'h4):(2'h2)]);
            end
          for (forvar1609 = (1'h0); (forvar1609 < (1'h0)); forvar1609 = (forvar1609 + (1'h1)))
            begin
              reg1610 <= reg1555[(2'h3):(1'h1)];
              reg1611 <= (+reg1574[(5'h17):(2'h2)]);
              reg1612 <= reg1539;
              reg1613 = (~({$unsigned((reg1608 + reg1546)),
                      $unsigned($signed(wire1529))} ?
                  reg1603 : ((^~{reg1540, reg1534}) ?
                      {$signed(reg1575),
                          reg1607[(3'h4):(1'h0)]} : ((reg1594 <= reg1587) ?
                          $signed(reg1575) : (-(8'hbb))))));
              reg1614 = (+($signed((^~$unsigned(reg1549))) == reg1553[(3'h4):(1'h1)]));
            end
        end
      else
        begin
          reg1603 = (~((&($signed(wire1531) ?
              reg1545[(1'h1):(1'h0)] : (wire1528 ?
                  reg1573 : reg1613))) - (|({(8'hb9),
              reg1549} <= $signed(wire1529)))));
          reg1604 <= ($signed((+(~(reg1548 ?
              reg1611 : wire1530)))) < ((((reg1602 && reg1614) ?
                  (reg1548 <<< reg1582) : reg1591[(4'h8):(3'h6)]) && (^~(^wire1532))) ?
              $unsigned(wire1530[(2'h2):(1'h0)]) : $unsigned({$unsigned(reg1613),
                  $signed(reg1613)})));
          reg1605 = reg1538;
          if (reg1552[(5'h13):(4'ha)])
            begin
              reg1607 = $signed($unsigned($signed($unsigned(wire1601[(1'h0):(1'h0)]))));
              reg1609 = ((($signed($unsigned(reg1559)) <= $signed((!reg1546))) ?
                  wire1532 : $signed((^~(reg1577 != reg1571)))) && $unsigned(reg1608[(3'h7):(2'h2)]));
              reg1610 <= $unsigned((reg1594[(2'h3):(1'h1)] & (($signed((7'h41)) ?
                  (reg1539 | forvar1609) : reg1594) >> $signed((-reg1582)))));
              reg1613 = (reg1562[(3'h6):(1'h0)] ?
                  $unsigned(((|reg1611) & reg1587[(3'h7):(3'h6)])) : (+reg1563));
              reg1615 <= $unsigned(((({reg1534, reg1562} ?
                  (reg1534 ? reg1611 : wire1530) : (8'hbc)) == ((reg1546 ?
                      reg1548 : reg1545) ?
                  $signed((8'hbc)) : reg1577[(1'h0):(1'h0)])) ^~ (8'hb1)));
            end
          else
            begin
              reg1607 = (~|reg1606);
              reg1609 = {$unsigned($unsigned($unsigned((reg1545 >> (7'h42))))),
                  (reg1585[(1'h1):(1'h1)] >>> ((!(~|(8'hb3))) >= $signed($signed(reg1540))))};
            end
        end
    end
  assign wire1616 = wire1528;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1227
#(parameter param1452 = (!((^~(((8'ha8) - (8'hb6)) ? {(8'hbb), (8'h9d)} : {(8'ha7)})) ? ((((8'hb6) & (8'hb9)) > {(7'h45)}) ~^ ((7'h49) ~^ (-(8'hbf)))) : ({((7'h41) <<< (8'hba))} ? (((8'ha8) ? (8'hab) : (8'ha4)) ? (-(8'ha6)) : ((8'hb7) | (7'h43))) : ({(8'h9e), (8'hae)} ? {(8'h9f), (8'hb8)} : {(8'hbb)})))))
(y, clk, wire1232, wire1231, wire1230, wire1229, wire1228);
  output wire [(32'hb4f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire1232;
  input wire [(5'h16):(1'h0)] wire1231;
  input wire signed [(2'h2):(1'h0)] wire1230;
  input wire [(2'h2):(1'h0)] wire1229;
  input wire [(5'h12):(1'h0)] wire1228;
  wire [(3'h6):(1'h0)] wire1425;
  wire [(5'h11):(1'h0)] wire1423;
  wire signed [(4'h8):(1'h0)] wire1422;
  wire signed [(5'h16):(1'h0)] wire1421;
  wire [(4'h8):(1'h0)] wire1326;
  wire signed [(5'h17):(1'h0)] wire1296;
  wire [(2'h2):(1'h0)] wire1244;
  reg signed [(2'h2):(1'h0)] reg1450 = (1'h0);
  reg [(4'h8):(1'h0)] reg1447 = (1'h0);
  reg [(5'h16):(1'h0)] reg1442 = (1'h0);
  reg [(4'h8):(1'h0)] reg1441 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1440 = (1'h0);
  reg [(5'h18):(1'h0)] reg1438 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1437 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1436 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1430 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1426 = (1'h0);
  reg [(5'h18):(1'h0)] reg1420 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1419 = (1'h0);
  reg [(3'h6):(1'h0)] reg1418 = (1'h0);
  reg [(4'ha):(1'h0)] reg1415 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1414 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1413 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1410 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1408 = (1'h0);
  reg [(3'h4):(1'h0)] reg1407 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1405 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1401 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1397 = (1'h0);
  reg [(5'h18):(1'h0)] reg1396 = (1'h0);
  reg [(4'hb):(1'h0)] reg1393 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1392 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1391 = (1'h0);
  reg [(2'h2):(1'h0)] reg1387 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1386 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1385 = (1'h0);
  reg [(4'hf):(1'h0)] reg1382 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1379 = (1'h0);
  reg [(5'h13):(1'h0)] reg1377 = (1'h0);
  reg [(2'h3):(1'h0)] reg1376 = (1'h0);
  reg [(4'hb):(1'h0)] reg1375 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1369 = (1'h0);
  reg [(4'h9):(1'h0)] reg1364 = (1'h0);
  reg [(3'h5):(1'h0)] reg1362 = (1'h0);
  reg [(4'ha):(1'h0)] reg1357 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1356 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1353 = (1'h0);
  reg [(4'h8):(1'h0)] reg1351 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1347 = (1'h0);
  reg [(4'he):(1'h0)] reg1346 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1341 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1340 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1339 = (1'h0);
  reg [(4'ha):(1'h0)] reg1330 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1337 = (1'h0);
  reg [(2'h2):(1'h0)] reg1335 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1334 = (1'h0);
  reg [(3'h7):(1'h0)] reg1320 = (1'h0);
  reg [(3'h5):(1'h0)] reg1317 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1315 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1314 = (1'h0);
  reg [(3'h4):(1'h0)] reg1312 = (1'h0);
  reg [(5'h13):(1'h0)] reg1311 = (1'h0);
  reg [(4'h8):(1'h0)] reg1310 = (1'h0);
  reg [(5'h16):(1'h0)] reg1309 = (1'h0);
  reg [(3'h6):(1'h0)] reg1308 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1305 = (1'h0);
  reg [(3'h4):(1'h0)] reg1304 = (1'h0);
  reg [(5'h10):(1'h0)] reg1302 = (1'h0);
  reg [(3'h7):(1'h0)] reg1300 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1297 = (1'h0);
  reg [(5'h14):(1'h0)] reg1294 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1293 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1291 = (1'h0);
  reg [(4'he):(1'h0)] reg1289 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1282 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1280 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1279 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1276 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1274 = (1'h0);
  reg [(3'h4):(1'h0)] reg1270 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1269 = (1'h0);
  reg [(5'h11):(1'h0)] reg1267 = (1'h0);
  reg [(5'h10):(1'h0)] reg1264 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1261 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1258 = (1'h0);
  reg [(5'h11):(1'h0)] reg1256 = (1'h0);
  reg [(4'he):(1'h0)] reg1254 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1253 = (1'h0);
  reg [(4'he):(1'h0)] reg1251 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1249 = (1'h0);
  reg [(5'h14):(1'h0)] reg1246 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1242 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1241 = (1'h0);
  reg [(4'hd):(1'h0)] reg1240 = (1'h0);
  reg [(4'hb):(1'h0)] reg1238 = (1'h0);
  reg [(4'hf):(1'h0)] reg1234 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1237 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1451 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1449 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1448 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1446 = (1'h0);
  reg [(5'h14):(1'h0)] reg1445 = (1'h0);
  reg [(4'ha):(1'h0)] reg1444 = (1'h0);
  reg [(5'h10):(1'h0)] reg1443 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1439 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1435 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1434 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1433 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1432 = (1'h0);
  reg [(5'h14):(1'h0)] reg1431 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1429 = (1'h0);
  reg [(4'h8):(1'h0)] reg1428 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1427 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1424 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1417 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1416 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1412 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1411 = (1'h0);
  reg [(4'hd):(1'h0)] reg1409 = (1'h0);
  reg [(3'h7):(1'h0)] reg1406 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1404 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1403 = (1'h0);
  reg [(4'ha):(1'h0)] reg1402 = (1'h0);
  reg [(4'he):(1'h0)] forvar1400 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1399 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1398 = (1'h0);
  reg [(5'h13):(1'h0)] reg1395 = (1'h0);
  reg [(4'he):(1'h0)] forvar1394 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1390 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1389 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1388 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1384 = (1'h0);
  reg [(5'h18):(1'h0)] reg1383 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1381 = (1'h0);
  reg [(5'h18):(1'h0)] reg1380 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1378 = (1'h0);
  reg [(3'h4):(1'h0)] reg1374 = (1'h0);
  reg [(4'h8):(1'h0)] reg1373 = (1'h0);
  reg [(5'h12):(1'h0)] reg1372 = (1'h0);
  reg [(3'h5):(1'h0)] reg1371 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1370 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1368 = (1'h0);
  reg [(4'h8):(1'h0)] reg1367 = (1'h0);
  reg [(3'h5):(1'h0)] reg1366 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1365 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1363 = (1'h0);
  reg [(4'he):(1'h0)] reg1361 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1360 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1359 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1358 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1355 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1354 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1352 = (1'h0);
  reg [(3'h7):(1'h0)] reg1350 = (1'h0);
  reg [(4'hc):(1'h0)] reg1349 = (1'h0);
  reg [(2'h2):(1'h0)] reg1348 = (1'h0);
  reg [(5'h17):(1'h0)] reg1345 = (1'h0);
  reg [(5'h17):(1'h0)] reg1344 = (1'h0);
  reg [(4'hc):(1'h0)] reg1343 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1342 = (1'h0);
  reg [(4'he):(1'h0)] reg1338 = (1'h0);
  reg [(4'hb):(1'h0)] reg1336 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1333 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1332 = (1'h0);
  reg [(5'h15):(1'h0)] reg1331 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1330 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1329 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1328 = (1'h0);
  reg [(4'he):(1'h0)] reg1327 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1316 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1325 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1324 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1323 = (1'h0);
  reg [(4'h9):(1'h0)] reg1322 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1321 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1319 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1318 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1316 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1313 = (1'h0);
  reg [(5'h16):(1'h0)] reg1307 = (1'h0);
  reg [(5'h18):(1'h0)] reg1306 = (1'h0);
  reg [(4'hd):(1'h0)] reg1303 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1301 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1299 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1298 = (1'h0);
  reg [(5'h12):(1'h0)] reg1295 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1292 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1290 = (1'h0);
  reg [(3'h5):(1'h0)] reg1288 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1287 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1286 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1285 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1284 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1277 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1273 = (1'h0);
  reg [(3'h4):(1'h0)] reg1283 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1281 = (1'h0);
  reg [(5'h16):(1'h0)] reg1278 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1277 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1275 = (1'h0);
  reg [(3'h7):(1'h0)] reg1273 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1272 = (1'h0);
  reg [(3'h5):(1'h0)] reg1271 = (1'h0);
  reg [(5'h18):(1'h0)] reg1268 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1266 = (1'h0);
  reg [(4'he):(1'h0)] forvar1265 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1263 = (1'h0);
  reg [(5'h16):(1'h0)] reg1262 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1260 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1259 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1257 = (1'h0);
  reg [(3'h5):(1'h0)] reg1255 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1252 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1250 = (1'h0);
  reg [(4'h9):(1'h0)] reg1248 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1247 = (1'h0);
  reg [(5'h14):(1'h0)] reg1245 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1243 = (1'h0);
  reg [(4'h9):(1'h0)] reg1239 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1236 = (1'h0);
  reg [(4'hf):(1'h0)] reg1235 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1234 = (1'h0);
  reg [(5'h18):(1'h0)] reg1233 = (1'h0);
  assign y = {wire1425,
                 wire1423,
                 wire1422,
                 wire1421,
                 wire1326,
                 wire1296,
                 wire1244,
                 reg1450,
                 reg1447,
                 reg1442,
                 reg1441,
                 reg1440,
                 reg1438,
                 reg1437,
                 reg1436,
                 reg1430,
                 reg1426,
                 reg1420,
                 reg1419,
                 reg1418,
                 reg1415,
                 reg1414,
                 reg1413,
                 reg1410,
                 reg1408,
                 reg1407,
                 reg1405,
                 reg1401,
                 reg1397,
                 reg1396,
                 reg1393,
                 reg1392,
                 reg1391,
                 reg1387,
                 reg1386,
                 reg1385,
                 reg1382,
                 reg1379,
                 reg1377,
                 reg1376,
                 reg1375,
                 reg1369,
                 reg1364,
                 reg1362,
                 reg1357,
                 reg1356,
                 reg1353,
                 reg1351,
                 reg1347,
                 reg1346,
                 reg1341,
                 reg1340,
                 reg1339,
                 reg1330,
                 reg1337,
                 reg1335,
                 reg1334,
                 reg1320,
                 reg1317,
                 reg1315,
                 reg1314,
                 reg1312,
                 reg1311,
                 reg1310,
                 reg1309,
                 reg1308,
                 reg1305,
                 reg1304,
                 reg1302,
                 reg1300,
                 reg1297,
                 reg1294,
                 reg1293,
                 reg1291,
                 reg1289,
                 reg1282,
                 reg1280,
                 reg1279,
                 reg1276,
                 reg1274,
                 reg1270,
                 reg1269,
                 reg1267,
                 reg1264,
                 reg1261,
                 reg1258,
                 reg1256,
                 reg1254,
                 reg1253,
                 reg1251,
                 reg1249,
                 reg1246,
                 reg1242,
                 reg1241,
                 reg1240,
                 reg1238,
                 reg1234,
                 reg1237,
                 reg1451,
                 reg1449,
                 reg1448,
                 forvar1446,
                 reg1445,
                 reg1444,
                 reg1443,
                 reg1439,
                 forvar1435,
                 reg1434,
                 forvar1433,
                 reg1432,
                 reg1431,
                 reg1429,
                 reg1428,
                 forvar1427,
                 reg1424,
                 forvar1417,
                 reg1416,
                 forvar1412,
                 forvar1411,
                 reg1409,
                 reg1406,
                 reg1404,
                 reg1403,
                 reg1402,
                 forvar1400,
                 reg1399,
                 reg1398,
                 reg1395,
                 forvar1394,
                 forvar1390,
                 reg1389,
                 reg1388,
                 forvar1384,
                 reg1383,
                 reg1381,
                 reg1380,
                 reg1378,
                 reg1374,
                 reg1373,
                 reg1372,
                 reg1371,
                 forvar1370,
                 reg1368,
                 reg1367,
                 reg1366,
                 reg1365,
                 reg1363,
                 reg1361,
                 reg1360,
                 forvar1359,
                 reg1358,
                 reg1355,
                 reg1354,
                 forvar1352,
                 reg1350,
                 reg1349,
                 reg1348,
                 reg1345,
                 reg1344,
                 reg1343,
                 reg1342,
                 reg1338,
                 reg1336,
                 reg1333,
                 reg1332,
                 reg1331,
                 forvar1330,
                 reg1329,
                 forvar1328,
                 reg1327,
                 forvar1316,
                 reg1325,
                 reg1324,
                 forvar1323,
                 reg1322,
                 forvar1321,
                 reg1319,
                 reg1318,
                 reg1316,
                 reg1313,
                 reg1307,
                 reg1306,
                 reg1303,
                 reg1301,
                 reg1299,
                 forvar1298,
                 reg1295,
                 reg1292,
                 forvar1290,
                 reg1288,
                 reg1287,
                 reg1286,
                 forvar1285,
                 forvar1284,
                 reg1277,
                 forvar1273,
                 reg1283,
                 forvar1281,
                 reg1278,
                 forvar1277,
                 reg1275,
                 reg1273,
                 reg1272,
                 reg1271,
                 reg1268,
                 forvar1266,
                 forvar1265,
                 reg1263,
                 reg1262,
                 reg1260,
                 reg1259,
                 reg1257,
                 reg1255,
                 forvar1252,
                 reg1250,
                 reg1248,
                 forvar1247,
                 reg1245,
                 reg1243,
                 reg1239,
                 reg1236,
                 reg1235,
                 forvar1234,
                 reg1233,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned({wire1228[(5'h10):(5'h10)]}))
        begin
          reg1233 = wire1232;
          for (forvar1234 = (1'h0); (forvar1234 < (1'h0)); forvar1234 = (forvar1234 + (1'h1)))
            begin
              reg1235 = (wire1228[(3'h7):(3'h7)] & ({({forvar1234, reg1233} ?
                      {wire1229} : $unsigned(wire1228))} <= ($unsigned((~&wire1231)) ?
                  (((8'h9c) ? wire1228 : forvar1234) ?
                      (^~wire1232) : (wire1228 >> (8'hb4))) : $unsigned(((8'hbb) <<< wire1228)))));
              reg1236 = (8'had);
              reg1237 <= wire1232;
            end
        end
      else
        begin
          reg1234 <= (forvar1234 ? wire1229 : $unsigned(wire1228));
          reg1237 <= ($signed((wire1228[(2'h3):(1'h0)] & ((&reg1237) ?
              wire1232[(1'h1):(1'h1)] : wire1229))) || ((~^($signed(reg1233) ?
              $unsigned(forvar1234) : $unsigned(wire1228))) & $unsigned(((reg1237 && wire1229) ?
              ((8'hb1) ? wire1228 : reg1236) : {reg1236}))));
        end
      if (wire1230[(1'h1):(1'h0)])
        begin
          reg1238 <= {$unsigned((^~((reg1236 ?
                  reg1236 : reg1237) <<< reg1235[(4'hc):(2'h2)])))};
          reg1239 = {$unsigned($signed((!$signed(wire1232))))};
        end
      else
        begin
          reg1239 = $signed((~wire1229));
          reg1240 <= (!$signed(($unsigned(wire1231) ?
              (~|reg1238[(3'h4):(1'h1)]) : $signed(forvar1234[(3'h4):(2'h2)]))));
          reg1241 <= {reg1240};
          reg1242 <= reg1237;
          reg1243 = (wire1228[(4'hd):(4'hd)] && reg1238);
        end
    end
  assign wire1244 = reg1234;
  always
    @(posedge clk) begin
      reg1245 = $unsigned($signed(((((8'hbc) || reg1240) ?
              (wire1228 + wire1229) : $signed(wire1232)) ?
          $unsigned(((8'ha5) != wire1244)) : ($signed(reg1242) & (wire1244 ?
              wire1229 : reg1237)))));
      reg1246 <= ($unsigned((reg1241[(4'he):(4'hd)] < $signed((wire1228 > (8'hb0))))) >= ($signed((!(wire1231 <= wire1231))) != (($signed(wire1228) ?
          (reg1238 ? reg1245 : reg1245) : (reg1238 ?
              reg1234 : (7'h40))) * $signed($signed(reg1245)))));
      for (forvar1247 = (1'h0); (forvar1247 < (1'h0)); forvar1247 = (forvar1247 + (1'h1)))
        begin
          if ((-$unsigned((($signed((8'hb0)) ?
              wire1244 : (forvar1247 ?
                  (7'h43) : wire1231)) != ((reg1246 ~^ wire1230) & (-forvar1247))))))
            begin
              reg1248 = ((~({(reg1241 && wire1230)} ?
                      ((wire1244 < (7'h42)) != reg1234[(1'h1):(1'h0)]) : (((7'h46) ?
                          reg1246 : wire1229) ~^ (wire1228 || wire1229)))) ?
                  (wire1232 - {reg1238[(4'h9):(2'h2)]}) : forvar1247[(1'h0):(1'h0)]);
              reg1249 <= (~&wire1230[(2'h2):(1'h1)]);
              reg1250 = reg1241;
              reg1251 <= ((wire1228 ^~ (!((reg1234 ?
                      reg1240 : forvar1247) - $unsigned((8'hb3))))) ?
                  {$unsigned((+(reg1246 ? reg1240 : reg1238))),
                      {(reg1234 ?
                              (reg1234 ?
                                  reg1248 : wire1244) : $signed(reg1241))}} : $signed(($signed((wire1232 ?
                          reg1250 : wire1229)) ?
                      ({reg1238, reg1245} ?
                          wire1228 : $signed(forvar1247)) : $unsigned(wire1229[(1'h1):(1'h0)]))));
            end
          else
            begin
              reg1248 = (((-((|reg1240) ?
                      ((8'hb7) - wire1244) : reg1251[(3'h4):(3'h4)])) ?
                  reg1240 : ((&(!reg1249)) > (8'hab))) || (!($signed(wire1232[(4'h8):(4'h8)]) > reg1240)));
              reg1250 = $signed(((-reg1234[(1'h1):(1'h0)]) ?
                  $unsigned(reg1240) : $signed((wire1230[(1'h1):(1'h0)] & (reg1242 ?
                      reg1248 : reg1246)))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1252 = (1'h0); (forvar1252 < (3'h4)); forvar1252 = (forvar1252 + (1'h1)))
        begin
          if (reg1242[(2'h3):(1'h1)])
            begin
              reg1253 <= $unsigned((($unsigned(((8'ha1) ?
                      (8'hb3) : (8'h9d))) < ($unsigned(reg1251) ^~ (forvar1252 ?
                      wire1228 : reg1237))) ?
                  (~|(reg1249[(2'h2):(2'h2)] ?
                      (~^wire1229) : forvar1252)) : (8'haf)));
              reg1254 <= {$signed(wire1228)};
              reg1255 = $unsigned(reg1242[(3'h4):(1'h0)]);
              reg1256 <= $unsigned({reg1234[(1'h0):(1'h0)]});
              reg1257 = ($unsigned(wire1232) <= (~|$signed($unsigned(reg1242[(5'h10):(3'h5)]))));
            end
          else
            begin
              reg1255 = (reg1240[(4'hd):(4'h9)] ?
                  wire1244[(2'h2):(2'h2)] : (^~forvar1252[(1'h0):(1'h0)]));
              reg1257 = $signed($signed(($unsigned($unsigned(reg1241)) + reg1237[(5'h12):(5'h12)])));
              reg1258 <= $signed($unsigned((({wire1229} ?
                      $unsigned((8'ha1)) : wire1231) ?
                  ($signed(reg1246) ?
                      (&(8'hbc)) : $unsigned(wire1231)) : reg1238)));
            end
          reg1259 = (~|forvar1252);
          if (((^wire1231[(3'h5):(1'h1)]) * $unsigned($unsigned(wire1228[(3'h5):(3'h4)]))))
            begin
              reg1260 = wire1229[(1'h1):(1'h0)];
              reg1261 <= (8'hac);
              reg1262 = ((((reg1246[(5'h10):(3'h5)] ?
                              {(8'hb5), (8'hb9)} : (^~wire1231)) ?
                          reg1240 : $signed($unsigned(reg1260))) ?
                      $signed((+(wire1229 + reg1260))) : $signed((|$signed(wire1231)))) ?
                  ($unsigned((~&reg1242)) == (({wire1244, reg1234} ?
                      {reg1256,
                          reg1259} : reg1261) << $unsigned($signed(wire1229)))) : reg1249);
              reg1263 = $signed((|$signed((wire1244 ?
                  (~|(8'ha7)) : $signed(wire1232)))));
            end
          else
            begin
              reg1261 <= $unsigned((((|reg1258) ?
                      $unsigned($signed(reg1251)) : (|wire1231[(2'h3):(1'h0)])) ?
                  {{$signed(reg1258), $signed(wire1228)}} : {(wire1244 ?
                          {(7'h49)} : reg1238)}));
            end
          reg1264 <= reg1251[(2'h2):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar1265 = (1'h0); (forvar1265 < (1'h1)); forvar1265 = (forvar1265 + (1'h1)))
        begin
          for (forvar1266 = (1'h0); (forvar1266 < (3'h4)); forvar1266 = (forvar1266 + (1'h1)))
            begin
              reg1267 <= wire1228[(4'ha):(2'h2)];
              reg1268 = $signed({((reg1261[(1'h0):(1'h0)] ?
                      $signed(reg1254) : {reg1253}) & reg1261[(4'hc):(2'h3)])});
            end
          reg1269 <= reg1261[(4'hb):(3'h7)];
          reg1270 <= ((reg1251 << (!reg1246)) >>> (forvar1265[(4'hd):(1'h1)] ?
              wire1231 : $signed(reg1261)));
        end
      reg1271 = (reg1258[(4'h9):(3'h5)] != ((wire1244[(1'h0):(1'h0)] + ((reg1242 ^ reg1234) ?
          (forvar1266 <<< reg1254) : (wire1231 <= wire1228))) == $signed(wire1229[(1'h1):(1'h0)])));
      if ((8'hb2))
        begin
          if ((~(reg1246 ? forvar1266 : (7'h41))))
            begin
              reg1272 = $unsigned((&(!(|((8'hb2) ? reg1254 : reg1242)))));
            end
          else
            begin
              reg1272 = wire1231;
              reg1273 = $signed(wire1244[(1'h1):(1'h1)]);
              reg1274 <= (^~wire1231[(4'ha):(2'h3)]);
              reg1275 = $signed($unsigned((&(8'h9c))));
              reg1276 <= $signed(({(^(|(7'h4a)))} ?
                  reg1242 : $signed($signed(reg1246))));
            end
          for (forvar1277 = (1'h0); (forvar1277 < (2'h2)); forvar1277 = (forvar1277 + (1'h1)))
            begin
              reg1278 = wire1230[(2'h2):(1'h1)];
              reg1279 <= $signed({(($signed(reg1246) ?
                      ((8'ha4) ?
                          reg1240 : reg1241) : wire1228[(3'h6):(2'h3)]) >= (reg1268[(3'h6):(2'h3)] >= (8'ha6)))});
              reg1280 <= reg1271[(2'h2):(1'h0)];
            end
          for (forvar1281 = (1'h0); (forvar1281 < (1'h1)); forvar1281 = (forvar1281 + (1'h1)))
            begin
              reg1282 <= $signed($unsigned((^reg1251)));
            end
          reg1283 = ((^{((7'h41) ? reg1258 : forvar1281),
              wire1232[(3'h5):(2'h3)]}) ^ ($signed({(reg1237 ?
                      wire1231 : reg1271)}) ?
              reg1280[(4'h8):(4'h8)] : reg1270));
        end
      else
        begin
          reg1272 = $unsigned((7'h43));
          for (forvar1273 = (1'h0); (forvar1273 < (2'h3)); forvar1273 = (forvar1273 + (1'h1)))
            begin
              reg1275 = (((reg1264[(2'h3):(2'h2)] >> reg1249) << $unsigned(((~reg1249) ?
                      {reg1275} : {reg1234}))) ?
                  $unsigned($unsigned($signed({(7'h42), reg1238}))) : wire1230);
              reg1276 <= ((^~forvar1281) - $unsigned($signed((reg1282[(2'h3):(1'h1)] ?
                  ((8'hb9) ? wire1232 : reg1240) : ((7'h43) ?
                      reg1240 : forvar1273)))));
              reg1277 = (((^~(~|forvar1265[(4'he):(1'h0)])) <= $signed((!reg1251))) + $signed((({reg1275,
                      reg1251} ?
                  (reg1246 ? reg1268 : reg1274) : (reg1267 ?
                      reg1276 : reg1282)) == {{(8'hbf)}, forvar1265})));
              reg1278 = ((($signed((!wire1232)) ?
                      reg1271 : (reg1242 ? $unsigned(reg1249) : reg1268)) ?
                  {((reg1234 <= (7'h48)) <= reg1278),
                      ($signed((8'ha5)) ?
                          $unsigned(reg1277) : (~&(8'h9d)))} : reg1241) && {(((+reg1261) ?
                          forvar1277[(3'h5):(1'h0)] : {(8'haa), wire1229}) ?
                      ($unsigned(wire1232) | reg1280) : ($signed(reg1238) ?
                          $unsigned(reg1278) : (^(8'hab))))});
              reg1279 <= reg1280;
            end
          reg1280 <= {reg1268[(4'hc):(4'h9)],
              ($unsigned((|(reg1280 + reg1256))) | {((|(8'ha9)) ?
                      $unsigned(reg1264) : (reg1283 == reg1234)),
                  reg1283[(2'h2):(1'h1)]})};
        end
      for (forvar1284 = (1'h0); (forvar1284 < (1'h1)); forvar1284 = (forvar1284 + (1'h1)))
        begin
          for (forvar1285 = (1'h0); (forvar1285 < (2'h2)); forvar1285 = (forvar1285 + (1'h1)))
            begin
              reg1286 = ($signed(reg1267[(5'h11):(4'he)]) ?
                  reg1280 : $signed(reg1241[(4'he):(4'hb)]));
              reg1287 = ((($signed(((8'ha2) ? wire1229 : reg1237)) ?
                      ((reg1274 ? wire1230 : reg1274) ?
                          $unsigned(reg1269) : reg1279) : {$signed(wire1229)}) ?
                  reg1269[(2'h2):(1'h1)] : (($signed(reg1242) ?
                          $unsigned(reg1234) : (~|reg1269)) ?
                      $unsigned({reg1270, reg1254}) : ({reg1274,
                          reg1267} >> (forvar1281 ?
                          reg1253 : reg1280)))) << $unsigned((7'h49)));
              reg1288 = ((~^reg1282[(1'h0):(1'h0)]) >> $signed(($unsigned((reg1276 != (7'h48))) ?
                  reg1286 : (reg1273[(3'h5):(2'h3)] ?
                      (~reg1268) : (~|reg1280)))));
              reg1289 <= reg1254;
            end
          for (forvar1290 = (1'h0); (forvar1290 < (1'h0)); forvar1290 = (forvar1290 + (1'h1)))
            begin
              reg1291 <= (^~((reg1238 ^ $signed((reg1242 ?
                      reg1287 : forvar1277))) ?
                  {(reg1242 ^~ (|reg1246))} : $signed((forvar1284 - reg1256))));
              reg1292 = ((~&$signed({(!reg1275)})) + (!(reg1253 ?
                  (~&$unsigned(reg1240)) : (~reg1273[(1'h0):(1'h0)]))));
              reg1293 <= (^~reg1272);
              reg1294 <= (&(forvar1285[(5'h14):(4'hb)] ?
                  $unsigned(reg1279[(1'h0):(1'h0)]) : ($signed($signed(reg1234)) ?
                      wire1228[(2'h3):(2'h2)] : $unsigned(wire1232[(2'h3):(2'h2)]))));
              reg1295 = {{$signed($signed($unsigned((8'hb7)))),
                      forvar1290[(3'h6):(1'h1)]}};
            end
        end
    end
  assign wire1296 = $unsigned((reg1234[(3'h5):(2'h3)] ?
                        $signed((reg1246 || ((8'hb0) ?
                            reg1291 : reg1294))) : (^($unsigned(reg1264) ^ $unsigned(reg1237)))));
  always
    @(posedge clk) begin
      reg1297 <= $unsigned($signed($signed(($signed(reg1282) ?
          reg1251 : (reg1267 != reg1249)))));
      for (forvar1298 = (1'h0); (forvar1298 < (3'h4)); forvar1298 = (forvar1298 + (1'h1)))
        begin
          reg1299 = $signed(reg1264);
          if (reg1249[(4'h9):(1'h0)])
            begin
              reg1300 <= ($unsigned($signed($signed((wire1231 ?
                      reg1240 : reg1297)))) ?
                  ({{reg1299[(3'h6):(2'h2)]},
                      ((^wire1228) + $signed(reg1267))} == wire1229) : (8'h9f));
              reg1301 = reg1241;
              reg1302 <= reg1249;
              reg1303 = reg1254[(4'h9):(3'h4)];
              reg1304 <= (^reg1261);
            end
          else
            begin
              reg1301 = {reg1249[(4'hc):(4'h8)], reg1241};
              reg1302 <= ($signed(reg1276[(3'h5):(1'h0)]) - reg1253[(2'h3):(1'h0)]);
              reg1304 <= reg1253;
              reg1305 <= ($unsigned($unsigned(reg1261[(1'h1):(1'h1)])) ?
                  ((^({reg1258, wire1232} || (wire1244 < reg1264))) ?
                      reg1304[(3'h4):(1'h1)] : reg1302) : ((($signed((7'h41)) ?
                          (reg1291 ?
                              wire1231 : reg1267) : (reg1258 == reg1269)) ?
                      reg1302 : reg1256[(4'hb):(1'h0)]) || ((reg1258[(4'he):(4'hd)] ?
                      reg1303 : (reg1289 << reg1251)) <= (8'hb8))));
              reg1306 = reg1253;
            end
          reg1307 = $signed(reg1297);
        end
      reg1308 <= {({(~|(reg1242 | (8'hb9)))} >>> {((reg1291 ?
                  wire1229 : wire1244) || $unsigned(wire1296)),
              $signed($unsigned(reg1301))})};
      reg1309 <= (reg1242 <= reg1240[(4'hb):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg1310 <= (wire1230 ?
          (~&(^~(reg1294[(3'h7):(1'h1)] >>> (reg1251 ?
              reg1270 : reg1300)))) : reg1269);
      reg1311 <= reg1304[(1'h0):(1'h0)];
      reg1312 <= {(reg1241 << reg1310)};
      if (($unsigned(((wire1244[(2'h2):(2'h2)] ?
          {(8'ha0)} : (~wire1231)) + $unsigned($unsigned(reg1274)))) == {(|reg1291[(1'h1):(1'h0)])}))
        begin
          reg1313 = (((^(!(reg1269 ? reg1249 : reg1249))) ?
              reg1280 : (({reg1276} ?
                      ((8'hb0) ?
                          wire1228 : reg1280) : wire1228[(4'h8):(3'h6)]) ?
                  $signed((reg1261 - (8'hb3))) : (((8'hae) >= wire1229) ?
                      $unsigned(reg1293) : $signed(wire1296)))) ^~ $signed(reg1270[(1'h1):(1'h0)]));
        end
      else
        begin
          reg1314 <= reg1297[(2'h3):(1'h1)];
        end
      if (($signed($unsigned($unsigned(((7'h46) ?
          reg1305 : wire1231)))) || ((8'ha4) ?
          reg1280 : reg1279[(2'h3):(2'h3)])))
        begin
          reg1315 <= ((~|$signed(((reg1237 ^ wire1296) ?
                  $unsigned(reg1279) : $unsigned(reg1282)))) ?
              $signed(reg1241) : {$signed(($signed(reg1267) - $signed(reg1314)))});
          reg1316 = $signed((~^$unsigned($signed(reg1279))));
          if ($unsigned((+$signed(wire1229))))
            begin
              reg1317 <= $signed({(^wire1229[(1'h0):(1'h0)]),
                  reg1304[(2'h3):(1'h0)]});
              reg1318 = reg1289[(4'hd):(4'hb)];
              reg1319 = ((reg1313 | $unsigned((~reg1242))) ?
                  $unsigned($signed($unsigned((reg1237 ?
                      reg1254 : reg1293)))) : reg1261[(3'h5):(2'h3)]);
              reg1320 <= $unsigned($signed($signed(((+reg1317) ?
                  $signed(wire1244) : reg1293))));
            end
          else
            begin
              reg1318 = ($unsigned(reg1256) ?
                  ((&(-(&reg1270))) ?
                      reg1276 : (^~{wire1229[(2'h2):(2'h2)]})) : $signed(reg1267));
            end
          for (forvar1321 = (1'h0); (forvar1321 < (1'h0)); forvar1321 = (forvar1321 + (1'h1)))
            begin
              reg1322 = (($unsigned(reg1311) ? reg1258 : (^reg1238)) & reg1258);
            end
          for (forvar1323 = (1'h0); (forvar1323 < (2'h3)); forvar1323 = (forvar1323 + (1'h1)))
            begin
              reg1324 = wire1230;
              reg1325 = (~(|reg1311));
            end
        end
      else
        begin
          reg1315 <= reg1320[(1'h1):(1'h0)];
          for (forvar1316 = (1'h0); (forvar1316 < (2'h3)); forvar1316 = (forvar1316 + (1'h1)))
            begin
              reg1318 = $unsigned((~(forvar1316[(2'h2):(1'h1)] ?
                  $signed($signed(reg1237)) : (-reg1311[(4'he):(4'ha)]))));
            end
          reg1320 <= reg1258[(1'h1):(1'h1)];
          for (forvar1321 = (1'h0); (forvar1321 < (2'h3)); forvar1321 = (forvar1321 + (1'h1)))
            begin
              reg1322 = forvar1321[(5'h14):(3'h6)];
            end
        end
    end
  assign wire1326 = $signed(((reg1280 * $signed((~reg1314))) ?
                        (&{{(8'hb0), (8'hb8)},
                            (reg1308 <= wire1229)}) : (|($signed(reg1256) ?
                            (reg1256 <<< reg1304) : (~&reg1304)))));
  always
    @(posedge clk) begin
      reg1327 = reg1253[(3'h7):(2'h2)];
      if ({$signed(reg1320), reg1305})
        begin
          for (forvar1328 = (1'h0); (forvar1328 < (2'h2)); forvar1328 = (forvar1328 + (1'h1)))
            begin
              reg1329 = $signed((-reg1289[(3'h4):(3'h4)]));
            end
          for (forvar1330 = (1'h0); (forvar1330 < (3'h4)); forvar1330 = (forvar1330 + (1'h1)))
            begin
              reg1331 = reg1246;
              reg1332 = (reg1256 ^~ (reg1308[(1'h1):(1'h0)] ^ $signed(wire1296[(5'h15):(5'h12)])));
              reg1333 = $signed($signed($signed({forvar1328})));
              reg1334 <= ((&((8'ha9) ?
                  (reg1264[(4'hd):(1'h1)] ?
                      $unsigned(reg1238) : reg1254) : wire1231)) >>> (($unsigned(wire1231) ?
                      ((^reg1297) || $unsigned(reg1315)) : reg1256[(5'h11):(2'h2)]) ?
                  $unsigned(reg1309) : $unsigned(($signed(reg1302) - (8'hac)))));
            end
          if (reg1334)
            begin
              reg1335 <= ((reg1309 ?
                      ($signed((reg1251 ^~ reg1276)) * ($signed(reg1315) ?
                          (reg1305 * reg1264) : (|(8'hb8)))) : $signed(((reg1300 && (7'h44)) ?
                          {reg1317, reg1251} : reg1274))) ?
                  ($signed((^~$signed(reg1269))) < (&wire1230[(1'h0):(1'h0)])) : (|reg1291));
            end
          else
            begin
              reg1336 = $signed(({(8'hb8)} ?
                  ($signed($unsigned(wire1231)) < ((^~reg1320) == (~reg1329))) : $signed(wire1232[(3'h7):(1'h0)])));
              reg1337 <= reg1312;
            end
        end
      else
        begin
          for (forvar1328 = (1'h0); (forvar1328 < (2'h2)); forvar1328 = (forvar1328 + (1'h1)))
            begin
              reg1330 <= {wire1232, forvar1330};
              reg1334 <= $unsigned(($signed($signed($unsigned(reg1269))) ?
                  (^~$signed(reg1308[(3'h4):(1'h1)])) : ($signed(reg1304[(1'h0):(1'h0)]) || (^~reg1329[(5'h10):(4'h9)]))));
              reg1336 = (-($signed(($unsigned((8'hbf)) ?
                  {(8'hb1)} : $signed(reg1291))) * wire1232[(2'h2):(1'h1)]));
            end
          if (reg1276[(5'h15):(1'h0)])
            begin
              reg1337 <= (7'h41);
              reg1338 = ($signed((+(reg1291[(1'h0):(1'h0)] ?
                      $signed(reg1320) : reg1241[(3'h7):(2'h3)]))) ?
                  reg1305[(3'h6):(2'h3)] : (~^(reg1282[(2'h2):(1'h1)] ?
                      reg1234[(1'h1):(1'h1)] : ((|reg1311) > $unsigned(wire1229)))));
              reg1339 <= ($unsigned(reg1334[(1'h0):(1'h0)]) >= $signed(reg1258));
              reg1340 <= reg1334;
            end
          else
            begin
              reg1337 <= ($unsigned($unsigned(reg1330)) << $signed((^~(reg1256 ?
                  $signed((8'ha2)) : reg1297))));
              reg1339 <= reg1314;
              reg1340 <= {(&reg1331),
                  (reg1338 <<< (&{reg1312[(1'h0):(1'h0)]}))};
              reg1341 <= ($unsigned((|(reg1258[(4'he):(3'h7)] ?
                  reg1339 : (+reg1340)))) + reg1282[(2'h3):(2'h3)]);
              reg1342 = $unsigned({(+reg1276)});
            end
          if ($unsigned($unsigned(((8'h9e) ^ (~^(~&reg1270))))))
            begin
              reg1343 = $unsigned({($signed(reg1261) ?
                      (reg1339 ?
                          reg1312 : (8'haf)) : $signed(reg1294[(4'hf):(4'h9)]))});
              reg1344 = (+reg1331);
              reg1345 = (((reg1311[(5'h10):(4'h8)] ^ reg1338[(2'h2):(2'h2)]) <= $unsigned((!reg1341))) >>> ({(-((8'ha1) + reg1294)),
                      (~|wire1229[(1'h0):(1'h0)])} ?
                  (~|($signed(reg1291) << (reg1294 <<< wire1228))) : (reg1270[(2'h2):(1'h1)] ?
                      (&$signed(reg1317)) : ({wire1228} ^ {reg1274}))));
              reg1346 <= (|reg1267[(5'h11):(4'h9)]);
            end
          else
            begin
              reg1343 = reg1258[(5'h11):(4'h9)];
              reg1346 <= $unsigned(reg1289[(1'h0):(1'h0)]);
              reg1347 <= (~$signed((($unsigned(reg1270) ?
                  $unsigned(wire1231) : (reg1300 ?
                      reg1302 : forvar1328)) ^ $signed((~^reg1246)))));
            end
          if ($unsigned($unsigned((reg1336[(4'ha):(4'h9)] <<< ({wire1229} ^ ((7'h46) ?
              reg1346 : reg1258))))))
            begin
              reg1348 = wire1228;
              reg1349 = (-reg1249);
              reg1350 = $signed($signed($signed(reg1291[(3'h4):(2'h3)])));
            end
          else
            begin
              reg1351 <= reg1334[(1'h1):(1'h1)];
            end
          for (forvar1352 = (1'h0); (forvar1352 < (2'h2)); forvar1352 = (forvar1352 + (1'h1)))
            begin
              reg1353 <= $signed($unsigned((~^reg1302)));
              reg1354 = reg1334;
              reg1355 = reg1340[(3'h7):(2'h3)];
              reg1356 <= (^~reg1338[(4'h8):(3'h7)]);
            end
        end
      reg1357 <= wire1230;
      reg1358 = reg1294;
    end
  always
    @(posedge clk) begin
      for (forvar1359 = (1'h0); (forvar1359 < (1'h0)); forvar1359 = (forvar1359 + (1'h1)))
        begin
          reg1360 = {reg1300[(3'h5):(3'h4)]};
        end
      if ((&reg1256))
        begin
          if ($signed($unsigned({(reg1309 + (~&wire1326)),
              $signed(((8'haf) || reg1314))})))
            begin
              reg1361 = ({$unsigned($signed((-reg1346)))} < (~|$signed($unsigned((reg1315 > reg1308)))));
              reg1362 <= $signed(reg1237[(1'h0):(1'h0)]);
              reg1363 = $unsigned(reg1356);
              reg1364 <= {reg1256[(1'h0):(1'h0)],
                  $unsigned(reg1237[(5'h10):(4'hf)])};
              reg1365 = reg1267[(4'ha):(1'h1)];
            end
          else
            begin
              reg1361 = $unsigned(reg1254[(2'h3):(1'h0)]);
              reg1362 <= reg1340[(4'hb):(4'h9)];
              reg1363 = $signed($unsigned((((reg1317 ?
                      (8'hb5) : reg1251) <= $signed(reg1300)) ?
                  (-$signed(reg1241)) : (reg1365 ?
                      (reg1353 ? reg1320 : reg1315) : $unsigned(reg1304)))));
            end
        end
      else
        begin
          reg1361 = $signed(reg1249[(3'h7):(3'h4)]);
          reg1363 = $signed((wire1229[(2'h2):(2'h2)] ?
              {reg1351} : (-((wire1244 != reg1317) <= (reg1347 ?
                  reg1337 : reg1294)))));
        end
      reg1366 = $unsigned(reg1311[(4'hb):(1'h0)]);
      if ($unsigned($unsigned($unsigned($signed((-reg1341))))))
        begin
          reg1367 = (~^reg1337[(1'h1):(1'h0)]);
          reg1368 = reg1240[(3'h6):(3'h4)];
        end
      else
        begin
          if ((!{$signed($signed((~|reg1364))),
              ($signed($signed(reg1270)) > (^(reg1340 <<< (8'hac))))}))
            begin
              reg1369 <= ((({reg1320[(3'h7):(1'h1)]} - $signed((reg1261 || reg1242))) >= (-$unsigned((reg1335 + reg1361)))) && $signed(((reg1267 ?
                      reg1310[(4'h8):(3'h5)] : $signed(reg1294)) ?
                  ($signed(reg1347) ? reg1251 : reg1249) : reg1367)));
            end
          else
            begin
              reg1367 = (-(^~($signed({reg1330}) ?
                  (^~(~reg1368)) : $signed(reg1309))));
              reg1369 <= (~|($unsigned(reg1274[(2'h2):(1'h1)]) > (~&reg1267)));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1370 = (1'h0); (forvar1370 < (1'h1)); forvar1370 = (forvar1370 + (1'h1)))
        begin
          if (reg1364[(4'h8):(3'h7)])
            begin
              reg1371 = $unsigned(reg1276);
              reg1372 = reg1314;
              reg1373 = $unsigned({(-(&(!(7'h49))))});
              reg1374 = (~|reg1373[(4'h8):(4'h8)]);
              reg1375 <= {$signed(((8'ha6) ?
                      {$unsigned(forvar1370),
                          reg1261[(4'h9):(3'h6)]} : $signed(reg1357[(4'h9):(3'h5)]))),
                  $signed(reg1305)};
            end
          else
            begin
              reg1375 <= $signed(reg1369[(5'h17):(1'h1)]);
              reg1376 <= (7'h4a);
            end
        end
      if ($unsigned($signed($unsigned((7'h47)))))
        begin
          reg1377 <= reg1282[(2'h3):(1'h1)];
          if ((reg1242[(1'h1):(1'h1)] & $unsigned(reg1341)))
            begin
              reg1378 = (~reg1369[(5'h18):(4'hb)]);
              reg1379 <= (~^wire1228[(4'he):(2'h2)]);
              reg1380 = (^(~|$signed({$unsigned(reg1264)})));
              reg1381 = (^~reg1254[(4'hc):(4'hc)]);
              reg1382 <= reg1373;
            end
          else
            begin
              reg1379 <= reg1369[(4'hb):(3'h5)];
            end
          reg1383 = $unsigned($unsigned(reg1373[(3'h5):(3'h4)]));
          for (forvar1384 = (1'h0); (forvar1384 < (2'h3)); forvar1384 = (forvar1384 + (1'h1)))
            begin
              reg1385 <= (reg1240[(3'h5):(1'h0)] ?
                  (+$signed(reg1335)) : $unsigned({($unsigned(reg1374) + $unsigned(reg1276))}));
              reg1386 <= wire1296;
              reg1387 <= $unsigned($unsigned({(-(reg1314 - (8'hb0))),
                  $signed(reg1339[(2'h2):(2'h2)])}));
              reg1388 = ($unsigned((8'haa)) ?
                  (|reg1246) : {$signed((reg1369[(3'h7):(3'h4)] == reg1381[(2'h2):(1'h1)])),
                      (~&reg1309[(3'h7):(1'h0)])});
              reg1389 = $signed($unsigned($unsigned(reg1346)));
            end
          for (forvar1390 = (1'h0); (forvar1390 < (1'h1)); forvar1390 = (forvar1390 + (1'h1)))
            begin
              reg1391 <= (~^$unsigned(($unsigned({wire1229}) ^~ reg1335[(1'h0):(1'h0)])));
              reg1392 <= ((~|reg1375) <= reg1378);
              reg1393 <= $unsigned($unsigned(({forvar1390[(1'h1):(1'h1)],
                  $signed(reg1289)} < reg1270[(1'h1):(1'h0)])));
            end
        end
      else
        begin
          if ((|{reg1249[(4'h8):(3'h4)]}))
            begin
              reg1378 = {$signed(($signed($signed(reg1387)) ?
                      ((^~(8'hbe)) ^~ $unsigned(reg1392)) : (~^reg1387[(1'h0):(1'h0)])))};
            end
          else
            begin
              reg1377 <= (^~reg1294[(5'h12):(4'ha)]);
              reg1378 = reg1379[(3'h4):(3'h4)];
            end
          reg1379 <= (^~(8'ha6));
        end
    end
  always
    @(posedge clk) begin
      for (forvar1394 = (1'h0); (forvar1394 < (2'h2)); forvar1394 = (forvar1394 + (1'h1)))
        begin
          if (reg1357[(3'h6):(3'h5)])
            begin
              reg1395 = (-reg1364[(3'h6):(1'h1)]);
            end
          else
            begin
              reg1395 = (-((+(wire1232 ?
                  {reg1391} : reg1280[(2'h2):(1'h1)])) <= reg1302[(3'h6):(3'h5)]));
            end
          if ($signed(wire1232[(1'h0):(1'h0)]))
            begin
              reg1396 <= $signed((reg1315[(1'h0):(1'h0)] & (reg1310[(3'h5):(3'h5)] | {{reg1356}})));
              reg1397 <= (^(~(~&(~|(reg1396 ? wire1232 : reg1294)))));
              reg1398 = ($signed((&($unsigned(reg1362) == reg1377))) ^~ (~^reg1294[(5'h13):(2'h2)]));
            end
          else
            begin
              reg1398 = ({wire1230[(1'h1):(1'h1)]} - reg1314);
            end
          reg1399 = ((reg1289 ?
              reg1261[(4'ha):(3'h7)] : ($unsigned(reg1312[(2'h2):(1'h1)]) ?
                  {wire1229[(2'h2):(1'h0)]} : (reg1276 >= reg1264))) ~^ reg1308);
          for (forvar1400 = (1'h0); (forvar1400 < (1'h1)); forvar1400 = (forvar1400 + (1'h1)))
            begin
              reg1401 <= reg1261[(1'h1):(1'h0)];
              reg1402 = $signed((~&((reg1258 + reg1376) ^ $signed((-reg1261)))));
              reg1403 = reg1289[(4'hc):(4'hb)];
              reg1404 = (~&((&({reg1386, forvar1394} ?
                      reg1382[(3'h6):(2'h2)] : (|forvar1394))) ?
                  {$signed({(7'h40)}),
                      $unsigned((8'h9e))} : reg1376[(1'h0):(1'h0)]));
              reg1405 <= ((reg1310[(3'h6):(3'h6)] ?
                  $signed(wire1228[(4'hb):(3'h4)]) : $unsigned(reg1294[(5'h10):(2'h2)])) <= (reg1377[(4'hf):(1'h1)] != $signed($signed({reg1404}))));
            end
          if (reg1297)
            begin
              reg1406 = (^{($signed({reg1351}) ?
                      (reg1253[(2'h3):(2'h2)] ?
                          {reg1267} : (reg1369 != reg1337)) : $signed($unsigned(reg1289))),
                  (reg1309 ?
                      wire1326 : ($unsigned(reg1264) >>> $unsigned(reg1396)))});
              reg1407 <= $signed((8'h9f));
              reg1408 <= (((8'hbb) ?
                      $signed(((reg1294 < wire1244) ?
                          reg1334 : {reg1320,
                              reg1404})) : (($unsigned((8'hb6)) + (reg1311 <<< reg1407)) != reg1346[(3'h7):(1'h0)])) ?
                  $signed((7'h47)) : reg1258);
              reg1409 = (reg1276 * reg1397);
            end
          else
            begin
              reg1407 <= $unsigned($signed((reg1310[(2'h3):(2'h2)] ?
                  reg1251[(3'h6):(2'h3)] : ({reg1315} ?
                      (|reg1347) : (reg1405 <= (7'h48))))));
            end
        end
      reg1410 <= reg1356[(3'h6):(3'h6)];
      for (forvar1411 = (1'h0); (forvar1411 < (2'h3)); forvar1411 = (forvar1411 + (1'h1)))
        begin
          for (forvar1412 = (1'h0); (forvar1412 < (2'h2)); forvar1412 = (forvar1412 + (1'h1)))
            begin
              reg1413 <= (!reg1369[(5'h17):(4'h9)]);
              reg1414 <= (^~(reg1393 ?
                  ($signed($unsigned(reg1353)) ?
                      reg1357[(4'h8):(3'h4)] : $unsigned({reg1240})) : (reg1341 ?
                      ((8'hba) == (reg1269 && reg1302)) : reg1312[(3'h4):(1'h0)])));
              reg1415 <= {$unsigned($unsigned((^{reg1386}))),
                  ((((!reg1238) ?
                              reg1357[(4'ha):(3'h5)] : ((7'h42) ?
                                  reg1375 : reg1341)) ?
                          $unsigned(reg1269[(3'h5):(3'h4)]) : $unsigned((reg1410 < reg1254))) ?
                      $signed(reg1254[(2'h2):(2'h2)]) : $signed(reg1305))};
            end
          reg1416 = reg1242[(5'h10):(4'hb)];
          for (forvar1417 = (1'h0); (forvar1417 < (2'h2)); forvar1417 = (forvar1417 + (1'h1)))
            begin
              reg1418 <= reg1395;
              reg1419 <= $unsigned((({(+reg1312)} | reg1406[(2'h2):(2'h2)]) ?
                  ($signed((+wire1326)) ?
                      reg1314[(2'h2):(2'h2)] : $signed($signed(reg1300))) : $signed((((8'hba) ?
                          reg1386 : (8'h9d)) ?
                      (~wire1296) : $unsigned(reg1254)))));
              reg1420 <= $unsigned($signed(wire1244[(1'h0):(1'h0)]));
            end
        end
    end
  assign wire1421 = reg1330[(1'h1):(1'h0)];
  assign wire1422 = (^reg1420);
  assign wire1423 = wire1326[(4'h8):(3'h7)];
  always
    @(posedge clk) begin
      reg1424 = $unsigned(wire1422);
    end
  assign wire1425 = (reg1376[(1'h0):(1'h0)] ?
                        reg1258[(5'h15):(1'h0)] : $signed($signed($unsigned((wire1296 * reg1376)))));
  always
    @(posedge clk) begin
      reg1426 <= $unsigned($signed(reg1415));
      for (forvar1427 = (1'h0); (forvar1427 < (2'h3)); forvar1427 = (forvar1427 + (1'h1)))
        begin
          if (reg1238)
            begin
              reg1428 = reg1376;
              reg1429 = (($unsigned(({reg1302, wire1421} ?
                  (^reg1237) : (reg1379 ? (8'ha6) : reg1305))) + (~(wire1326 ?
                  $signed(reg1346) : reg1280[(3'h7):(3'h7)]))) >>> ({$unsigned(((8'ha0) ?
                      reg1397 : (8'ha3)))} != (reg1375 ^~ reg1241)));
              reg1430 <= $unsigned(reg1385[(2'h3):(1'h1)]);
            end
          else
            begin
              reg1428 = reg1362;
              reg1430 <= (reg1420 & (reg1382[(3'h6):(1'h0)] > ((reg1309[(4'ha):(4'h8)] ?
                  wire1232[(1'h0):(1'h0)] : $unsigned(reg1396)) == {(7'h42),
                  reg1264})));
              reg1431 = (((wire1230 ? reg1305 : wire1230) | (7'h49)) ?
                  reg1393 : reg1293[(4'hf):(3'h4)]);
              reg1432 = (~(((8'ha1) >> (8'h9d)) ?
                  ({$unsigned(reg1410), (reg1414 ? reg1309 : reg1430)} ?
                      (reg1429 & (^reg1305)) : ((wire1296 ?
                          reg1428 : reg1234) ^ (reg1337 > reg1293))) : (~^{reg1305[(3'h7):(2'h3)]})));
            end
          for (forvar1433 = (1'h0); (forvar1433 < (1'h1)); forvar1433 = (forvar1433 + (1'h1)))
            begin
              reg1434 = ($signed($signed((reg1375 * wire1228))) >> reg1302[(3'h4):(1'h1)]);
            end
          for (forvar1435 = (1'h0); (forvar1435 < (3'h4)); forvar1435 = (forvar1435 + (1'h1)))
            begin
              reg1436 <= ($unsigned($signed(reg1317)) ?
                  $unsigned((($unsigned(reg1267) ?
                          (^~reg1420) : $signed(wire1296)) ?
                      (reg1242[(2'h3):(1'h1)] - reg1353[(2'h2):(2'h2)]) : ((reg1241 ?
                          reg1317 : reg1311) << reg1300[(3'h4):(2'h3)]))) : reg1413[(3'h4):(1'h1)]);
              reg1437 <= reg1351;
            end
          if ($unsigned({$unsigned($unsigned((reg1254 - reg1317))),
              reg1261[(1'h1):(1'h0)]}))
            begin
              reg1438 <= (wire1228[(4'ha):(4'h8)] + {reg1310[(4'h8):(2'h2)]});
              reg1439 = $unsigned(((8'h9e) * forvar1435[(3'h4):(1'h0)]));
              reg1440 <= reg1320;
              reg1441 <= $signed(((&(&reg1364)) || reg1434));
              reg1442 <= $unsigned((-({$signed(reg1304), {reg1337}} ?
                  ($unsigned((8'hb0)) ?
                      (reg1415 << reg1293) : (reg1351 ^ reg1405)) : ($signed(reg1405) ?
                      reg1357[(3'h4):(3'h4)] : reg1414))));
            end
          else
            begin
              reg1439 = (-{reg1312,
                  ($unsigned(reg1364[(2'h2):(2'h2)]) || (reg1261 ?
                      reg1387[(1'h1):(1'h0)] : reg1347[(3'h5):(3'h5)]))});
              reg1440 <= (((~^forvar1433) && (!reg1337)) > reg1340);
              reg1443 = reg1274[(3'h5):(2'h2)];
              reg1444 = reg1401[(1'h0):(1'h0)];
              reg1445 = (((8'hae) ?
                  $signed($unsigned((8'ha4))) : reg1434) ~^ {reg1294,
                  $unsigned(reg1379[(4'hb):(2'h2)])});
            end
        end
      for (forvar1446 = (1'h0); (forvar1446 < (1'h0)); forvar1446 = (forvar1446 + (1'h1)))
        begin
          if ({reg1282[(1'h0):(1'h0)]})
            begin
              reg1447 <= {(($unsigned(wire1228) + ((reg1240 ?
                      (8'ha4) : (8'hb4)) == reg1310[(1'h0):(1'h0)])) < (|(~&(^~reg1397))))};
            end
          else
            begin
              reg1448 = reg1413[(2'h3):(2'h3)];
              reg1449 = (8'hb9);
            end
        end
      reg1450 <= $unsigned((($unsigned((^reg1428)) ?
              ((reg1293 ^ reg1254) & $unsigned(reg1251)) : $unsigned(reg1249[(3'h5):(3'h4)])) ?
          ($signed(reg1251[(3'h6):(2'h2)]) ?
              reg1334 : $signed((reg1447 < reg1410))) : (reg1393 || (7'h42))));
      reg1451 = (^(!$unsigned((~^(reg1434 ~^ reg1294)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module903
#(parameter param1065 = (^~(&(!((~|(8'hb2)) && ((8'hac) > (8'hb7)))))))
(y, clk, wire907, wire906, wire905, wire904);
  output wire [(32'h7b5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire907;
  input wire [(3'h5):(1'h0)] wire906;
  input wire signed [(5'h18):(1'h0)] wire905;
  input wire [(4'ha):(1'h0)] wire904;
  wire signed [(3'h7):(1'h0)] wire996;
  wire signed [(5'h10):(1'h0)] wire995;
  wire [(5'h15):(1'h0)] wire972;
  wire signed [(5'h17):(1'h0)] wire965;
  wire [(3'h5):(1'h0)] wire964;
  wire [(5'h10):(1'h0)] wire963;
  wire signed [(3'h5):(1'h0)] wire908;
  reg [(5'h10):(1'h0)] reg1063 = (1'h0);
  reg [(5'h18):(1'h0)] reg1061 = (1'h0);
  reg [(2'h2):(1'h0)] reg1059 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1057 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1056 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1053 = (1'h0);
  reg [(4'ha):(1'h0)] reg1051 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1041 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1052 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1046 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1045 = (1'h0);
  reg [(3'h6):(1'h0)] reg1044 = (1'h0);
  reg [(4'ha):(1'h0)] reg1043 = (1'h0);
  reg [(4'h9):(1'h0)] reg1038 = (1'h0);
  reg [(3'h5):(1'h0)] reg1035 = (1'h0);
  reg [(4'hd):(1'h0)] reg1034 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1031 = (1'h0);
  reg [(4'hf):(1'h0)] reg1030 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1028 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1027 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1026 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1023 = (1'h0);
  reg [(5'h12):(1'h0)] reg1022 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1021 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1019 = (1'h0);
  reg [(4'he):(1'h0)] reg1018 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1015 = (1'h0);
  reg [(4'h8):(1'h0)] reg1014 = (1'h0);
  reg [(4'h9):(1'h0)] reg1008 = (1'h0);
  reg [(5'h10):(1'h0)] reg1010 = (1'h0);
  reg [(4'ha):(1'h0)] reg1009 = (1'h0);
  reg [(4'hb):(1'h0)] reg1007 = (1'h0);
  reg [(4'h9):(1'h0)] reg1005 = (1'h0);
  reg [(2'h2):(1'h0)] reg1002 = (1'h0);
  reg [(3'h5):(1'h0)] reg998 = (1'h0);
  reg [(4'h8):(1'h0)] reg994 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg993 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg992 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg991 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg988 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg987 = (1'h0);
  reg [(4'h8):(1'h0)] reg983 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg985 = (1'h0);
  reg [(3'h4):(1'h0)] reg984 = (1'h0);
  reg [(3'h5):(1'h0)] reg980 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg978 = (1'h0);
  reg [(3'h7):(1'h0)] reg977 = (1'h0);
  reg [(5'h10):(1'h0)] reg976 = (1'h0);
  reg [(5'h17):(1'h0)] reg971 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg959 = (1'h0);
  reg [(4'hf):(1'h0)] reg957 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg951 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg956 = (1'h0);
  reg signed [(4'he):(1'h0)] reg955 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg952 = (1'h0);
  reg [(5'h17):(1'h0)] reg949 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg948 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg947 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg946 = (1'h0);
  reg [(5'h14):(1'h0)] reg944 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg943 = (1'h0);
  reg [(4'h9):(1'h0)] reg941 = (1'h0);
  reg [(4'hb):(1'h0)] reg938 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg936 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg935 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg933 = (1'h0);
  reg [(5'h10):(1'h0)] reg930 = (1'h0);
  reg [(2'h2):(1'h0)] reg929 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg928 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg926 = (1'h0);
  reg [(4'hc):(1'h0)] reg924 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg923 = (1'h0);
  reg [(2'h3):(1'h0)] reg919 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg916 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg914 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg913 = (1'h0);
  reg [(4'hd):(1'h0)] reg912 = (1'h0);
  reg [(4'hc):(1'h0)] reg910 = (1'h0);
  reg [(5'h11):(1'h0)] reg1064 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1062 = (1'h0);
  reg [(2'h3):(1'h0)] reg1060 = (1'h0);
  reg [(5'h13):(1'h0)] reg1058 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1055 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1054 = (1'h0);
  reg [(4'h9):(1'h0)] reg1047 = (1'h0);
  reg [(3'h6):(1'h0)] reg1039 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1038 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1051 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1050 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1049 = (1'h0);
  reg [(2'h2):(1'h0)] reg1048 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1047 = (1'h0);
  reg [(2'h2):(1'h0)] reg1042 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1041 = (1'h0);
  reg [(5'h16):(1'h0)] reg1040 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1039 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1037 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1036 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1033 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1032 = (1'h0);
  reg [(4'hf):(1'h0)] reg1029 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1025 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1025 = (1'h0);
  reg [(4'hc):(1'h0)] reg1024 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1020 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1017 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1016 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1013 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1008 = (1'h0);
  reg [(3'h5):(1'h0)] reg1006 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1004 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1003 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1001 = (1'h0);
  reg [(3'h6):(1'h0)] reg1000 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg999 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar997 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg990 = (1'h0);
  reg [(5'h17):(1'h0)] reg989 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg986 = (1'h0);
  reg [(2'h2):(1'h0)] forvar983 = (1'h0);
  reg [(4'h9):(1'h0)] reg982 = (1'h0);
  reg [(5'h12):(1'h0)] reg981 = (1'h0);
  reg [(3'h4):(1'h0)] forvar979 = (1'h0);
  reg [(3'h5):(1'h0)] forvar975 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg974 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg973 = (1'h0);
  reg [(4'h8):(1'h0)] reg970 = (1'h0);
  reg [(2'h2):(1'h0)] reg969 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg968 = (1'h0);
  reg [(4'hb):(1'h0)] forvar967 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar966 = (1'h0);
  reg [(3'h5):(1'h0)] reg962 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg961 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg960 = (1'h0);
  reg [(5'h17):(1'h0)] reg958 = (1'h0);
  reg signed [(4'he):(1'h0)] reg954 = (1'h0);
  reg [(4'hf):(1'h0)] reg953 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar951 = (1'h0);
  reg [(5'h14):(1'h0)] reg950 = (1'h0);
  reg [(4'he):(1'h0)] reg945 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg942 = (1'h0);
  reg [(3'h4):(1'h0)] reg940 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg939 = (1'h0);
  reg signed [(4'he):(1'h0)] reg937 = (1'h0);
  reg [(5'h16):(1'h0)] forvar934 = (1'h0);
  reg [(4'hb):(1'h0)] reg932 = (1'h0);
  reg [(5'h15):(1'h0)] reg931 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg927 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg925 = (1'h0);
  reg [(5'h12):(1'h0)] reg920 = (1'h0);
  reg [(3'h7):(1'h0)] reg922 = (1'h0);
  reg [(3'h6):(1'h0)] reg921 = (1'h0);
  reg [(2'h2):(1'h0)] forvar920 = (1'h0);
  reg [(5'h13):(1'h0)] reg918 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg917 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar915 = (1'h0);
  reg [(5'h12):(1'h0)] forvar911 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg909 = (1'h0);
  assign y = {wire996,
                 wire995,
                 wire972,
                 wire965,
                 wire964,
                 wire963,
                 wire908,
                 reg1063,
                 reg1061,
                 reg1059,
                 reg1057,
                 reg1056,
                 reg1053,
                 reg1051,
                 reg1041,
                 reg1052,
                 reg1046,
                 reg1045,
                 reg1044,
                 reg1043,
                 reg1038,
                 reg1035,
                 reg1034,
                 reg1031,
                 reg1030,
                 reg1028,
                 reg1027,
                 reg1026,
                 reg1023,
                 reg1022,
                 reg1021,
                 reg1019,
                 reg1018,
                 reg1015,
                 reg1014,
                 reg1008,
                 reg1010,
                 reg1009,
                 reg1007,
                 reg1005,
                 reg1002,
                 reg998,
                 reg994,
                 reg993,
                 reg992,
                 reg991,
                 reg988,
                 reg987,
                 reg983,
                 reg985,
                 reg984,
                 reg980,
                 reg978,
                 reg977,
                 reg976,
                 reg971,
                 reg959,
                 reg957,
                 reg951,
                 reg956,
                 reg955,
                 reg952,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 reg944,
                 reg943,
                 reg941,
                 reg938,
                 reg936,
                 reg935,
                 reg933,
                 reg930,
                 reg929,
                 reg928,
                 reg926,
                 reg924,
                 reg923,
                 reg919,
                 reg916,
                 reg914,
                 reg913,
                 reg912,
                 reg910,
                 reg1064,
                 forvar1062,
                 reg1060,
                 reg1058,
                 forvar1055,
                 forvar1054,
                 reg1047,
                 reg1039,
                 forvar1038,
                 forvar1051,
                 reg1050,
                 reg1049,
                 reg1048,
                 forvar1047,
                 reg1042,
                 forvar1041,
                 reg1040,
                 forvar1039,
                 reg1037,
                 reg1036,
                 reg1033,
                 reg1032,
                 reg1029,
                 reg1025,
                 forvar1025,
                 reg1024,
                 reg1020,
                 reg1017,
                 forvar1016,
                 reg1013,
                 reg1012,
                 reg1011,
                 forvar1008,
                 reg1006,
                 forvar1004,
                 reg1003,
                 reg1001,
                 reg1000,
                 reg999,
                 forvar997,
                 reg990,
                 reg989,
                 reg986,
                 forvar983,
                 reg982,
                 reg981,
                 forvar979,
                 forvar975,
                 reg974,
                 reg973,
                 reg970,
                 reg969,
                 reg968,
                 forvar967,
                 forvar966,
                 reg962,
                 reg961,
                 reg960,
                 reg958,
                 reg954,
                 reg953,
                 forvar951,
                 reg950,
                 reg945,
                 reg942,
                 reg940,
                 reg939,
                 reg937,
                 forvar934,
                 reg932,
                 reg931,
                 reg927,
                 reg925,
                 reg920,
                 reg922,
                 reg921,
                 forvar920,
                 reg918,
                 reg917,
                 forvar915,
                 forvar911,
                 reg909,
                 (1'h0)};
  assign wire908 = (wire907 && (^wire907[(4'h9):(2'h2)]));
  always
    @(posedge clk) begin
      reg909 = ($signed(($unsigned((wire905 ? (8'hb2) : (8'hbf))) ?
              $unsigned((wire904 ?
                  (8'hb2) : wire908)) : (~|wire904[(1'h1):(1'h1)]))) ?
          (wire906[(1'h1):(1'h0)] ?
              (wire906 ?
                  (wire907 ?
                      (^wire905) : (wire904 || wire906)) : $unsigned(wire908)) : (($signed((8'hb1)) ?
                  $signed(wire908) : (~&wire907)) > wire904)) : (8'haa));
      reg910 <= $unsigned((|$signed(wire908[(2'h3):(1'h0)])));
      for (forvar911 = (1'h0); (forvar911 < (2'h3)); forvar911 = (forvar911 + (1'h1)))
        begin
          reg912 <= $unsigned((wire904 ? wire906 : reg910));
          reg913 <= (8'hb2);
          reg914 <= $unsigned((($unsigned(wire906) ?
              (reg913 >> wire907[(3'h6):(3'h4)]) : reg913) <= wire905));
          for (forvar915 = (1'h0); (forvar915 < (2'h3)); forvar915 = (forvar915 + (1'h1)))
            begin
              reg916 <= wire905[(5'h11):(4'hc)];
            end
        end
      reg917 = $unsigned(reg912);
    end
  always
    @(posedge clk) begin
      reg918 = {({wire907[(3'h6):(3'h4)]} ?
              ($signed({(7'h4a)}) ?
                  ((+(8'h9e)) + $signed(reg914)) : wire905[(1'h0):(1'h0)]) : (~|((wire904 <<< reg916) ?
                  $signed(wire907) : (reg912 & reg916)))),
          (-(8'hb9))};
      if (reg916[(4'hc):(4'hb)])
        begin
          reg919 <= (|((~|(|((7'h42) ?
              reg914 : (7'h45)))) <= $signed((wire907 | $unsigned(reg916)))));
          for (forvar920 = (1'h0); (forvar920 < (2'h3)); forvar920 = (forvar920 + (1'h1)))
            begin
              reg921 = (^(reg913[(4'ha):(4'h9)] ?
                  (~&(reg916[(3'h4):(1'h0)] ?
                      $signed((7'h48)) : {wire905})) : reg919));
              reg922 = reg916[(4'hb):(3'h6)];
              reg923 <= {((($unsigned((8'hae)) ?
                      (wire905 ?
                          (8'hb8) : reg916) : wire908[(1'h0):(1'h0)]) <<< reg910[(4'h9):(1'h1)]) < (wire907[(4'ha):(3'h6)] >> ((reg912 ?
                          wire904 : reg914) ?
                      (reg919 ^ wire904) : $unsigned(wire904))))};
              reg924 <= wire908;
            end
        end
      else
        begin
          reg920 = reg924;
          if (reg912)
            begin
              reg921 = (~^$signed((($signed(wire906) ~^ (^reg910)) | $unsigned((8'hb5)))));
            end
          else
            begin
              reg923 <= ($unsigned((reg924[(3'h4):(2'h2)] ?
                  reg924 : (reg924[(3'h6):(2'h2)] >= forvar920[(2'h2):(1'h1)]))) ^ reg914[(3'h4):(2'h2)]);
              reg924 <= {(~^(-$unsigned(reg918)))};
              reg925 = $signed(($signed(wire906[(3'h5):(2'h3)]) ?
                  $signed(((reg914 ? reg921 : reg919) ?
                      (|wire904) : ((8'had) ? wire908 : (8'ha3)))) : (8'h9f)));
              reg926 <= reg925;
            end
          if ($signed(forvar920[(1'h0):(1'h0)]))
            begin
              reg927 = reg920[(2'h2):(2'h2)];
              reg928 <= (wire908[(3'h4):(2'h3)] ?
                  $signed(({{reg925,
                          (8'hb5)}} >>> reg923[(2'h3):(2'h3)])) : $signed($signed($unsigned((reg910 ?
                      wire905 : (7'h42))))));
              reg929 <= (8'hb0);
              reg930 <= (($unsigned($unsigned((-reg918))) > $unsigned($signed($unsigned(reg919)))) ?
                  $signed($signed(((reg927 >>> wire906) * wire908))) : reg913);
            end
          else
            begin
              reg928 <= (-(^~{reg920}));
              reg931 = reg930[(1'h1):(1'h1)];
            end
          reg932 = $signed((($signed(reg910) << (+{reg930, reg929})) ?
              $signed(reg922) : $signed((+$unsigned(wire905)))));
          reg933 <= {(reg921 - $unsigned(reg929[(1'h0):(1'h0)])),
              ((reg925[(4'hc):(2'h3)] <= (((8'had) < reg924) <= {reg922})) ?
                  (reg931[(4'hc):(3'h7)] ?
                      (((7'h42) >> (7'h44)) ?
                          $signed(reg912) : reg928[(3'h7):(2'h2)]) : ((^(8'hac)) ?
                          reg924[(3'h5):(2'h2)] : reg918[(2'h2):(1'h1)])) : reg919)};
        end
    end
  always
    @(posedge clk) begin
      for (forvar934 = (1'h0); (forvar934 < (3'h4)); forvar934 = (forvar934 + (1'h1)))
        begin
          if (((!(((|reg919) << {reg916}) ?
                  $unsigned((reg919 + (8'h9c))) : reg924[(4'h9):(2'h3)])) ?
              $unsigned(((8'h9f) >>> (|(|wire906)))) : ($unsigned($unsigned({reg933})) >>> $unsigned(wire906[(2'h3):(1'h1)]))))
            begin
              reg935 <= wire906[(3'h5):(2'h3)];
              reg936 <= reg919[(1'h1):(1'h1)];
              reg937 = wire908;
              reg938 <= {$unsigned(reg910[(4'hc):(2'h2)])};
            end
          else
            begin
              reg937 = forvar934[(2'h2):(2'h2)];
              reg938 <= $signed(((8'ha6) ?
                  (($signed(reg938) ?
                      {reg933, reg928} : (reg937 ?
                          wire908 : reg924)) >= reg937[(2'h2):(1'h1)]) : reg919));
            end
          reg939 = (+(~{$signed((reg935 ~^ reg913)), (-(~|reg914))}));
          if (reg926[(2'h2):(1'h0)])
            begin
              reg940 = $unsigned($signed(reg924));
              reg941 <= {wire905};
            end
          else
            begin
              reg940 = (^$unsigned((reg938[(3'h6):(3'h6)] >= (|reg924[(4'h9):(3'h4)]))));
              reg942 = ((^~{reg912,
                  $signed(reg940[(2'h3):(1'h1)])}) ^~ $unsigned(($unsigned((reg938 ?
                  reg929 : reg926)) >= forvar934)));
              reg943 <= $unsigned(reg924[(4'h8):(1'h0)]);
              reg944 <= (8'hbf);
              reg945 = reg926;
            end
          reg946 <= $signed(((-((wire907 ?
              reg913 : reg926) == reg924[(3'h6):(1'h0)])) + (8'ha7)));
          if ($signed(reg942))
            begin
              reg947 <= {((({reg943, reg943} ^~ (^~reg923)) ?
                          (((8'hbb) >= reg937) ^ reg942[(1'h0):(1'h0)]) : wire907[(4'ha):(4'h8)]) ?
                      reg944[(4'hc):(4'hb)] : {((reg939 || reg910) ?
                              $unsigned(reg938) : $signed(wire905)),
                          (&(^reg942))})};
            end
          else
            begin
              reg947 <= (reg939 ?
                  ((|reg939[(4'h9):(3'h5)]) >>> reg923) : reg923);
              reg948 <= (|(({(reg916 ? reg939 : reg944),
                  $unsigned(reg930)} || ($signed(reg930) != $unsigned(reg937))) < (~reg928)));
            end
        end
      reg949 <= ($signed(($unsigned({reg919,
          reg928}) >>> reg914[(2'h3):(2'h3)])) >> $unsigned((&(-$signed(reg928)))));
      reg950 = $unsigned(wire908[(2'h2):(1'h1)]);
    end
  always
    @(posedge clk) begin
      if ((({$unsigned((reg913 ? reg947 : reg933))} ?
          {{(!reg919),
                  {(8'had),
                      reg919}}} : $signed((~&$unsigned(wire904)))) ^ ($unsigned(reg926) | ({{wire905}} ?
          $signed($unsigned(wire908)) : ((+reg912) <= reg912)))))
        begin
          for (forvar951 = (1'h0); (forvar951 < (2'h3)); forvar951 = (forvar951 + (1'h1)))
            begin
              reg952 <= reg941[(1'h0):(1'h0)];
              reg953 = $unsigned($unsigned($unsigned({(~reg944)})));
              reg954 = reg933;
              reg955 <= ($signed(((8'hbf) || wire905[(2'h3):(1'h1)])) ?
                  (-reg953[(3'h6):(3'h6)]) : $signed(reg954[(3'h7):(3'h6)]));
              reg956 <= forvar951[(1'h1):(1'h1)];
            end
        end
      else
        begin
          reg951 <= reg935[(2'h3):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned((reg913 ~^ {reg949, (!$unsigned((8'ha0)))})))
        begin
          reg957 <= ({{$signed((|(8'hb6)))}} ? (&$signed((8'hbc))) : reg933);
        end
      else
        begin
          reg957 <= reg941;
          reg958 = ((($unsigned(reg951[(3'h7):(3'h4)]) ?
                      ((reg948 >> reg912) ?
                          reg948 : (wire906 ? wire904 : reg943)) : ((~^reg947) ?
                          (8'ha9) : (reg956 ? reg910 : reg952))) ?
                  (wire905 ?
                      $signed((8'hbf)) : $signed((reg929 ?
                          reg944 : reg948))) : reg933) ?
              (8'h9f) : ($signed(((reg913 || reg947) ?
                  (+wire908) : wire904)) ^ ($signed((reg948 ?
                  reg912 : reg913)) <= ((wire905 ^~ reg924) ?
                  (reg948 ? wire908 : reg930) : (~^reg948)))));
          if ((8'ha4))
            begin
              reg959 <= reg930[(3'h4):(1'h1)];
              reg960 = (~|reg955[(3'h6):(3'h6)]);
              reg961 = ((~^reg933) || $unsigned((~$signed(reg924[(2'h2):(1'h1)]))));
              reg962 = (reg923 || wire906[(2'h2):(1'h1)]);
            end
          else
            begin
              reg960 = ($signed(wire904) ?
                  {((&$unsigned(reg913)) & ((reg924 & reg914) ?
                          $unsigned(reg933) : reg924)),
                      ($signed(reg928) ?
                          (wire907[(2'h3):(1'h0)] ?
                              ((7'h48) ?
                                  reg910 : reg959) : reg955[(2'h3):(2'h3)]) : (-$signed(wire904)))} : (wire905[(2'h2):(1'h0)] ?
                      ($unsigned((~reg960)) ?
                          {{reg913}} : ((reg951 ? wire907 : reg919) ?
                              $unsigned(reg955) : (wire907 ^~ wire908))) : $signed(($signed(reg948) ?
                          wire904[(3'h6):(1'h0)] : ((8'hb1) >>> reg962)))));
              reg961 = $signed((&$signed(reg947[(3'h7):(3'h5)])));
            end
        end
    end
  assign wire963 = $signed(reg929);
  assign wire964 = reg947;
  assign wire965 = (7'h44);
  always
    @(posedge clk) begin
      for (forvar966 = (1'h0); (forvar966 < (3'h4)); forvar966 = (forvar966 + (1'h1)))
        begin
          for (forvar967 = (1'h0); (forvar967 < (2'h2)); forvar967 = (forvar967 + (1'h1)))
            begin
              reg968 = reg929;
              reg969 = $signed($signed($unsigned((wire904 ?
                  reg933 : wire964))));
              reg970 = $unsigned({(({(8'ha2)} >> $signed(reg944)) > $signed({reg910}))});
              reg971 <= reg959;
            end
        end
    end
  assign wire972 = reg951[(4'h8):(3'h7)];
  always
    @(posedge clk) begin
      reg973 = $unsigned((|(((reg947 <<< reg926) ?
          wire905 : {reg926}) ^~ (|(reg959 ? (8'ha6) : reg946)))));
      reg974 = (^~((wire965 ?
          {wire908[(1'h1):(1'h0)], $signed(reg916)} : ((reg947 ?
              reg928 : reg947) * (^reg914))) & (wire908[(1'h0):(1'h0)] == $unsigned((&wire907)))));
      for (forvar975 = (1'h0); (forvar975 < (3'h4)); forvar975 = (forvar975 + (1'h1)))
        begin
          reg976 <= (^$signed(reg944[(4'he):(4'hc)]));
          reg977 <= wire964[(1'h1):(1'h0)];
          reg978 <= $signed(reg971[(3'h6):(3'h6)]);
          for (forvar979 = (1'h0); (forvar979 < (2'h3)); forvar979 = (forvar979 + (1'h1)))
            begin
              reg980 <= $unsigned(({wire965,
                  reg977} ^ $signed($unsigned($signed((8'hbf))))));
              reg981 = (reg980 ?
                  forvar979[(1'h0):(1'h0)] : $unsigned($signed(((reg913 * reg955) >= (reg947 != reg955)))));
            end
        end
      if ($unsigned(((~(7'h40)) || $unsigned(($signed(wire964) <= (reg947 ?
          wire963 : (7'h41)))))))
        begin
          reg982 = (($signed(reg941[(3'h4):(2'h2)]) ?
              $signed(reg941) : (8'had)) & (~|(8'ha2)));
          for (forvar983 = (1'h0); (forvar983 < (2'h2)); forvar983 = (forvar983 + (1'h1)))
            begin
              reg984 <= ((($signed((^reg952)) + reg941) ?
                      $signed(($signed(forvar975) - (reg910 ?
                          reg982 : wire906))) : {(reg913[(4'hb):(1'h1)] ?
                              {(8'ha2)} : reg948[(4'hc):(1'h1)]),
                          $signed({reg971})}) ?
                  {$unsigned(((reg944 ? forvar983 : reg952) || reg935)),
                      (reg959 <= $signed((reg980 < reg919)))} : $unsigned((8'ha2)));
              reg985 <= $signed((!$unsigned({wire905[(5'h17):(4'h8)],
                  {wire908, reg912}})));
            end
        end
      else
        begin
          reg983 <= reg959;
          if (reg973[(4'ha):(3'h6)])
            begin
              reg984 <= (~&reg938[(4'h9):(1'h0)]);
              reg986 = $signed(({$signed((reg983 ? reg930 : wire905)),
                  ((!reg974) ?
                      ((8'haf) ?
                          reg916 : wire907) : (wire972 | reg936))} == reg919));
              reg987 <= $unsigned(reg944[(4'hb):(2'h2)]);
              reg988 <= ($unsigned(((wire963[(4'hf):(1'h1)] > reg959) ?
                  $unsigned((~(8'hb0))) : reg987)) << reg951[(2'h3):(1'h1)]);
              reg989 = ((8'ha6) ?
                  $signed((~^$unsigned(reg941))) : (~|wire905[(5'h10):(3'h6)]));
            end
          else
            begin
              reg984 <= (($unsigned(((8'hb2) ?
                      (reg941 << (7'h45)) : (reg951 - reg913))) >> reg943) ?
                  $unsigned(reg943[(4'hb):(2'h2)]) : ((+$unsigned(reg982[(3'h5):(1'h0)])) >> ($signed($unsigned((8'ha3))) >> reg941)));
              reg986 = reg985[(2'h3):(1'h0)];
              reg987 <= wire906;
              reg988 <= $unsigned(reg912);
            end
          reg990 = (reg985 ^~ wire972);
          if (((($unsigned({reg919}) ? reg959[(1'h1):(1'h0)] : reg944) ?
                  reg971[(4'h8):(3'h6)] : ((8'hb3) != reg914[(4'ha):(4'ha)])) ?
              (~^{$unsigned(reg949)}) : $signed($unsigned(reg980))))
            begin
              reg991 <= wire904;
              reg992 <= $unsigned(reg936[(4'ha):(4'ha)]);
              reg993 <= (~^reg926[(1'h0):(1'h0)]);
              reg994 <= ((8'ha3) >>> ({reg949[(4'h8):(2'h2)],
                      $unsigned((!reg949))} ?
                  reg928[(2'h3):(2'h2)] : $unsigned($unsigned((forvar979 <<< reg912)))));
            end
          else
            begin
              reg991 <= {({$unsigned($unsigned((8'h9c))), (^$signed(reg946))} ?
                      reg944[(1'h1):(1'h0)] : wire907),
                  ({(reg994[(3'h5):(3'h5)] ?
                          $unsigned(wire965) : reg923)} << $unsigned($unsigned((reg938 ?
                      reg938 : reg982))))};
            end
        end
    end
  assign wire995 = ({({(reg936 ? reg938 : reg952)} >>> reg910[(2'h3):(1'h1)]),
                           reg933} ?
                       $signed($signed($signed(reg928))) : ($unsigned(({(8'hbf)} ?
                               $signed(reg955) : $signed(reg978))) ?
                           reg976 : (~^$unsigned({reg952, reg928}))));
  assign wire996 = ($signed(reg976) ?
                       (reg992 ?
                           (((reg914 << (8'h9c)) ?
                                   $unsigned(reg951) : $unsigned(wire907)) ?
                               reg956 : ($unsigned(wire905) >= {(8'haa),
                                   reg978})) : (({reg938} > reg957) >>> {(reg943 ?
                                   (8'hae) : reg983),
                               (reg988 * reg914)})) : {$unsigned({(reg985 ?
                                   wire963 : reg948)}),
                           wire965});
  always
    @(posedge clk) begin
      for (forvar997 = (1'h0); (forvar997 < (1'h1)); forvar997 = (forvar997 + (1'h1)))
        begin
          if ($unsigned(reg949[(5'h16):(5'h12)]))
            begin
              reg998 <= (8'hb3);
              reg999 = ((reg993 ~^ (&reg946[(1'h0):(1'h0)])) ?
                  wire906 : (~&wire906));
              reg1000 = wire996;
              reg1001 = (~|(reg992 ?
                  (^~({reg992} ?
                      $signed(reg992) : {reg949,
                          reg952})) : (reg991[(3'h7):(2'h3)] ?
                      {(^~(8'hbe))} : ($unsigned(reg924) * $unsigned(reg947)))));
              reg1002 <= {reg947[(2'h3):(2'h2)], reg944[(4'hc):(2'h2)]};
            end
          else
            begin
              reg999 = reg941[(2'h3):(2'h2)];
              reg1000 = (reg930[(3'h4):(1'h1)] ?
                  (reg928[(2'h3):(1'h1)] >> wire905) : reg928[(3'h6):(2'h3)]);
            end
          reg1003 = (reg998[(1'h1):(1'h1)] ?
              $unsigned((reg994 * reg923[(2'h3):(2'h3)])) : (!$unsigned(reg916)));
        end
      for (forvar1004 = (1'h0); (forvar1004 < (1'h0)); forvar1004 = (forvar1004 + (1'h1)))
        begin
          reg1005 <= (^$unsigned($signed($signed((reg916 ?
              reg998 : (7'h43))))));
          reg1006 = (~&(reg1001[(2'h3):(1'h1)] ?
              reg977 : (^~reg1002[(1'h0):(1'h0)])));
          reg1007 <= (+reg928[(3'h5):(1'h0)]);
        end
      if ($signed($unsigned($unsigned(wire907[(3'h4):(2'h2)]))))
        begin
          for (forvar1008 = (1'h0); (forvar1008 < (2'h3)); forvar1008 = (forvar1008 + (1'h1)))
            begin
              reg1009 <= {reg959, reg944[(3'h5):(3'h5)]};
              reg1010 <= reg951[(4'h9):(3'h6)];
              reg1011 = reg923[(2'h2):(1'h0)];
              reg1012 = $signed(reg984[(2'h2):(1'h1)]);
              reg1013 = wire964;
            end
        end
      else
        begin
          reg1008 <= reg991[(4'h9):(3'h5)];
        end
    end
  always
    @(posedge clk) begin
      if (reg956[(1'h1):(1'h0)])
        begin
          reg1014 <= (+$signed(({$signed(reg928)} ?
              $signed($signed((7'h4a))) : reg924[(1'h1):(1'h1)])));
          reg1015 <= $unsigned((~({((8'hb5) ? wire996 : reg993)} ?
              (~^$unsigned(reg1008)) : {reg1010[(3'h6):(1'h1)],
                  reg926[(1'h1):(1'h1)]})));
        end
      else
        begin
          reg1014 <= $signed(($unsigned((|((8'had) ? (8'hb7) : (8'hb8)))) ?
              reg980[(1'h0):(1'h0)] : ($unsigned(reg952[(3'h4):(3'h4)]) >> $signed($signed(reg944)))));
        end
      for (forvar1016 = (1'h0); (forvar1016 < (3'h4)); forvar1016 = (forvar1016 + (1'h1)))
        begin
          reg1017 = $signed((8'ha4));
          if (wire906[(3'h5):(2'h2)])
            begin
              reg1018 <= (-(~^{$signed((reg993 <<< reg1005))}));
              reg1019 <= $unsigned(((wire964[(3'h5):(3'h5)] == $signed({reg991})) ?
                  $unsigned($signed((wire963 ?
                      reg984 : reg978))) : $signed($signed(reg1005))));
            end
          else
            begin
              reg1018 <= $unsigned((wire965 ?
                  (((8'hb1) ?
                      (reg1019 ?
                          reg914 : (8'hb5)) : (reg944 && wire964)) != $unsigned((reg929 ?
                      reg947 : reg1008))) : reg978[(4'h8):(2'h2)]));
            end
          reg1020 = (7'h42);
          reg1021 <= $signed($signed({reg1008[(1'h1):(1'h1)]}));
          reg1022 <= ((~$signed((~&(reg913 ? reg991 : wire972)))) ?
              (reg971[(4'hd):(3'h4)] == ($signed($signed(reg1019)) <<< $signed($unsigned(reg991)))) : $unsigned((reg978[(4'hd):(4'ha)] ^~ (~&reg987))));
        end
      if ((^wire905))
        begin
          reg1023 <= (~$signed(reg928[(3'h6):(1'h0)]));
          reg1024 = $unsigned((!$signed($signed((reg943 || (8'ha4))))));
          for (forvar1025 = (1'h0); (forvar1025 < (2'h3)); forvar1025 = (forvar1025 + (1'h1)))
            begin
              reg1026 <= (&$signed($signed(((~&(8'hb6)) | (~^reg1009)))));
              reg1027 <= (7'h43);
              reg1028 <= reg983;
            end
        end
      else
        begin
          if ((!reg941))
            begin
              reg1023 <= {($unsigned(((~|reg985) || reg987)) ?
                      $signed(reg928[(3'h6):(1'h1)]) : (($signed(reg983) ?
                              reg1008 : $unsigned(reg924)) ?
                          ((wire907 ? reg947 : reg984) ?
                              (^~(8'hab)) : (~^reg1007)) : $unsigned((reg1017 ?
                              (8'ha0) : reg949))))};
              reg1024 = $signed((~^(^~$unsigned(reg985))));
              reg1025 = (~|$unsigned((((-(8'haf)) || (^reg936)) ^ (reg928[(2'h2):(1'h1)] <= reg984[(1'h1):(1'h1)]))));
              reg1029 = $signed((~&reg947));
            end
          else
            begin
              reg1024 = {(~|reg991[(4'hd):(2'h3)]),
                  (reg1020 ?
                      (&$unsigned(reg1023[(4'hd):(2'h2)])) : $unsigned($unsigned($signed(reg1018))))};
            end
          if (($signed(reg978) ~^ $signed((!($unsigned(reg930) ?
              reg955[(2'h3):(1'h1)] : reg1028[(3'h6):(1'h0)])))))
            begin
              reg1030 <= $unsigned(reg957);
              reg1031 <= ((!(~^$unsigned((reg977 >>> (8'haa))))) ?
                  $unsigned((^(reg944 << (reg1014 <= reg1021)))) : $signed(reg1021));
              reg1032 = $signed(($unsigned(reg1020[(3'h6):(2'h2)]) ?
                  (!(^$signed(reg1028))) : reg1019));
            end
          else
            begin
              reg1032 = $signed((($signed(reg924) ?
                  ({(8'ha2), forvar1025} ?
                      (~&wire972) : (+reg1020)) : {(reg959 <= reg1023)}) <<< reg987[(3'h5):(1'h1)]));
              reg1033 = $signed(reg928);
              reg1034 <= {(reg1017 * (reg1022 || (~&reg952))),
                  (-((~&{reg971, reg1008}) ?
                      ((reg1008 >>> reg959) | reg936) : $signed((reg980 || reg976))))};
            end
          reg1035 <= $signed(reg998);
          reg1036 = ((reg926[(3'h4):(1'h0)] ?
                  (reg1035 < $unsigned(reg943[(3'h5):(3'h5)])) : (8'hb7)) ?
              $unsigned(({$unsigned(reg935),
                  $signed(reg948)} ~^ (((8'haa) && wire908) ^~ $unsigned(reg924)))) : $unsigned(wire906[(3'h4):(2'h2)]));
          reg1037 = (((reg913 * reg913[(1'h0):(1'h0)]) | reg1022) ?
              {((~&reg1014) + ($unsigned(reg1017) & (-reg1002))),
                  (forvar1016[(5'h12):(1'h0)] ?
                      (reg1022 ?
                          (+reg1002) : $unsigned(reg912)) : wire963[(4'h9):(3'h4)])} : reg935);
        end
      if ((-reg938))
        begin
          reg1038 <= reg984[(3'h4):(2'h3)];
          for (forvar1039 = (1'h0); (forvar1039 < (1'h1)); forvar1039 = (forvar1039 + (1'h1)))
            begin
              reg1040 = $unsigned(wire905);
            end
          for (forvar1041 = (1'h0); (forvar1041 < (2'h3)); forvar1041 = (forvar1041 + (1'h1)))
            begin
              reg1042 = (-reg991);
              reg1043 <= {(reg1017 <= {reg913,
                      $signed(reg1031[(2'h3):(1'h0)])})};
              reg1044 <= reg946[(3'h5):(3'h4)];
              reg1045 <= reg1007[(3'h7):(1'h0)];
              reg1046 <= (&$signed(($signed(reg1023[(4'h8):(3'h4)]) ?
                  {{(8'hb5), reg1014}, $signed(wire964)} : reg1010)));
            end
          for (forvar1047 = (1'h0); (forvar1047 < (1'h0)); forvar1047 = (forvar1047 + (1'h1)))
            begin
              reg1048 = $unsigned($signed((+$signed(reg1019))));
              reg1049 = $unsigned((8'hb9));
              reg1050 = {wire907, forvar1025[(4'hd):(4'hb)]};
            end
          for (forvar1051 = (1'h0); (forvar1051 < (1'h0)); forvar1051 = (forvar1051 + (1'h1)))
            begin
              reg1052 <= ($unsigned((^{(reg1026 <= reg910),
                      $unsigned(reg1026)})) ?
                  (((&forvar1051) ?
                      (&(8'hbc)) : (~^(~^reg913))) ^~ reg1031[(3'h5):(2'h2)]) : (((!$signed(reg1023)) ?
                          (~$signed(reg952)) : ((reg998 >>> forvar1051) >> (reg1005 ?
                              (8'hac) : (8'hb6)))) ?
                      ({$unsigned(reg991)} ?
                          wire906 : ((reg983 >>> reg935) ?
                              reg952[(1'h0):(1'h0)] : (~&reg1027))) : ({$signed(wire965),
                              (|reg983)} ?
                          $unsigned(reg1031[(3'h5):(3'h4)]) : (~|(reg984 ?
                              reg1014 : reg1029)))));
            end
        end
      else
        begin
          for (forvar1038 = (1'h0); (forvar1038 < (1'h1)); forvar1038 = (forvar1038 + (1'h1)))
            begin
              reg1039 = $unsigned((((reg1018 < reg1037) ?
                      $signed(reg946[(3'h4):(3'h4)]) : ({reg924} + reg926[(1'h0):(1'h0)])) ?
                  ((!{reg1037, reg928}) ?
                      reg1023 : wire972) : $unsigned(reg928[(3'h5):(3'h5)])));
              reg1041 <= reg980[(1'h1):(1'h1)];
              reg1043 <= $unsigned($unsigned(reg1032[(4'hc):(4'h8)]));
              reg1047 = $signed((~^reg1032));
              reg1051 <= wire963;
            end
          if (({reg1044[(1'h1):(1'h0)]} ?
              reg935 : $unsigned((reg984 ?
                  (+$unsigned(reg947)) : (reg1051[(1'h0):(1'h0)] + $signed(reg993))))))
            begin
              reg1052 <= (reg1017[(1'h0):(1'h0)] ?
                  $unsigned(reg929) : $signed((reg919[(1'h0):(1'h0)] >> (8'hb3))));
            end
          else
            begin
              reg1052 <= (^~($unsigned((~$unsigned(forvar1047))) ~^ $signed($unsigned(reg923[(1'h0):(1'h0)]))));
              reg1053 <= $unsigned($unsigned((^reg1023[(3'h7):(3'h7)])));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1054 = (1'h0); (forvar1054 < (2'h2)); forvar1054 = (forvar1054 + (1'h1)))
        begin
          for (forvar1055 = (1'h0); (forvar1055 < (1'h1)); forvar1055 = (forvar1055 + (1'h1)))
            begin
              reg1056 <= $unsigned($signed($unsigned($signed($unsigned(reg946)))));
              reg1057 <= (reg936 ^ ($signed((|(^reg992))) ?
                  ($signed($signed(reg919)) ?
                      (8'h9f) : $signed(reg1030[(3'h6):(3'h5)])) : $unsigned(({wire972} && (|reg916)))));
              reg1058 = reg978[(4'hb):(3'h6)];
              reg1059 <= (~^$unsigned((~^$signed(wire963[(4'h9):(2'h3)]))));
              reg1060 = reg985;
            end
          reg1061 <= ({$signed($unsigned($unsigned(reg928))),
                  (reg1046[(2'h3):(2'h3)] & $unsigned($unsigned(reg938)))} ?
              (!(^~reg1022[(4'hc):(4'ha)])) : {reg977[(3'h6):(1'h0)],
                  wire972[(3'h7):(3'h6)]});
        end
      for (forvar1062 = (1'h0); (forvar1062 < (1'h0)); forvar1062 = (forvar1062 + (1'h1)))
        begin
          reg1063 <= ($signed({reg926, reg1038}) ?
              {(&((reg947 && reg1021) ?
                      reg949 : (reg926 <= (7'h49))))} : reg976[(4'h9):(3'h5)]);
        end
      reg1064 = wire995;
    end
endmodule