module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h2ad):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire4;
  input wire [(5'h14):(1'h0)] wire3;
  input wire [(5'h14):(1'h0)] wire2;
  input wire signed [(5'h14):(1'h0)] wire1;
  input wire signed [(4'he):(1'h0)] wire0;
  wire [(4'h8):(1'h0)] wire257;
  wire signed [(5'h14):(1'h0)] wire5;
  assign y = {wire257,
                 wire5,
                 (1'h0)};
  assign wire5 = $signed((wire4[(3'h4):(1'h0)] || {"fMR8T1MNO8l",
                     (^~(wire0 != wire1))}));
  module6 #() modinst258 (wire257, clk, wire1, wire0, wire5, wire3, wire2);

endmodule

module module6
#(parameter param256 = (8'hbe))
(y, clk, wire7, wire8, wire9, wire10, wire11);
  output wire [(32'h111):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire7;
  input wire signed [(4'hb):(1'h0)] wire8;
  input wire [(5'h14):(1'h0)] wire9;
  input wire [(4'hf):(1'h0)] wire10;
  input wire signed [(5'h14):(1'h0)] wire11;
  wire signed [(4'hd):(1'h0)] wire255;
  wire signed [(4'ha):(1'h0)] wire253;
  wire [(5'h12):(1'h0)] wire12;
  wire [(5'h10):(1'h0)] wire13;
  wire signed [(5'h11):(1'h0)] wire16;
  wire [(5'h11):(1'h0)] wire18;
  wire [(4'hf):(1'h0)] wire19;
  wire [(5'h14):(1'h0)] wire23;
  wire signed [(4'h8):(1'h0)] wire50;
  wire [(4'hd):(1'h0)] wire131;
  wire signed [(4'he):(1'h0)] wire133;
  wire [(3'h6):(1'h0)] wire134;
  wire signed [(4'hb):(1'h0)] wire135;
  wire [(4'h8):(1'h0)] wire136;
  wire [(4'hd):(1'h0)] wire139;
  wire signed [(2'h2):(1'h0)] wire221;
  reg [(3'h7):(1'h0)] reg137 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg14 = (1'h0);
  reg [(5'h13):(1'h0)] reg15 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg20 = (1'h0);
  reg [(2'h3):(1'h0)] reg22 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg138 = (1'h0);
  reg [(3'h5):(1'h0)] reg21 = (1'h0);
  assign y = {wire255,
                 wire253,
                 wire12,
                 wire13,
                 wire16,
                 wire18,
                 wire19,
                 wire23,
                 wire50,
                 wire131,
                 wire133,
                 wire134,
                 wire135,
                 wire136,
                 wire139,
                 wire221,
                 reg137,
                 reg14,
                 reg15,
                 reg17,
                 reg20,
                 reg22,
                 reg138,
                 reg21,
                 (1'h0)};
  assign wire12 = (|((8'ha6) ?
                      (wire9[(4'h8):(3'h6)] ?
                          {(+wire9)} : ($signed((8'hbb)) << "exAC")) : (wire8 ?
                          $unsigned("ET0uu6eXoYw4Tm3Q3") : (8'ha7))));
  assign wire13 = wire7[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg14 <= (|{(~wire12)});
      reg15 <= ($unsigned(reg14) ? wire12[(3'h4):(1'h0)] : (8'h9e));
    end
  assign wire16 = $unsigned((reg15 >> reg15[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      reg17 <= $unsigned($unsigned($signed($signed(wire16[(1'h1):(1'h0)]))));
    end
  assign wire18 = reg15[(4'ha):(1'h0)];
  assign wire19 = $unsigned(("cKoSmJ48qorGRxCb03" && ""));
  always
    @(posedge clk) begin
      reg20 <= wire10[(2'h3):(2'h2)];
      reg21 = (8'hbb);
      reg22 <= (8'hbd);
    end
  assign wire23 = ($unsigned(((8'hae) ? (8'hb2) : (~&$unsigned(reg20)))) ?
                      reg15 : (+"erJwkHhAHrMS"));
  module24 #() modinst51 (wire50, clk, wire11, wire16, wire18, reg22, wire12);
endmodule


module module24
#(parameter param48 = (8'hb9), 
parameter param49 = param48)
(y, clk, wire29, wire28, wire27, wire26, wire25);
  output wire [(32'hc8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire29;
  input wire signed [(4'hf):(1'h0)] wire28;
  input wire signed [(4'h8):(1'h0)] wire27;
  input wire [(2'h3):(1'h0)] wire26;
  input wire signed [(4'h9):(1'h0)] wire25;
  wire signed [(4'he):(1'h0)] wire47;
  wire [(4'ha):(1'h0)] wire30;
  reg signed [(5'h13):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg44 = (1'h0);
  reg [(4'h8):(1'h0)] reg43 = (1'h0);
  reg [(5'h15):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg41 = (1'h0);
  reg [(4'hd):(1'h0)] reg33 = (1'h0);
  reg [(4'hb):(1'h0)] reg38 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg37 = (1'h0);
  reg [(2'h2):(1'h0)] reg36 = (1'h0);
  reg [(3'h6):(1'h0)] reg35 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg34 = (1'h0);
  reg [(4'ha):(1'h0)] reg32 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg31 = (1'h0);
  reg [(2'h2):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg39 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar32 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar33 = (1'h0);
  assign y = {wire47,
                 wire30,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg33,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg32,
                 reg31,
                 reg40,
                 reg39,
                 forvar32,
                 forvar33,
                 (1'h0)};
  assign wire30 = wire25[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg31 <= ("f" ? wire27 : wire25[(3'h5):(3'h4)]);
      if ((~wire27[(3'h4):(2'h2)]))
        begin
          reg32 <= "OKvPnakTnuXarhK1wAIK";
          for (forvar33 = (1'h0); (forvar33 < (1'h1)); forvar33 = (forvar33 + (1'h1)))
            begin
              reg34 <= $signed((8'hba));
              reg35 <= ({(8'ha0)} ?
                  (((8'hac) ? (~^(8'ha6)) : $signed("hvTZ")) ?
                      "gyL4A" : wire28[(3'h5):(1'h0)]) : {wire29[(5'h11):(4'he)]});
              reg36 <= $signed(((|"VRr98") ?
                  wire29[(4'h8):(3'h6)] : ((~"IXQQKq4Gf") * "IPprfQ")));
              reg37 <= wire25;
            end
          reg38 <= $signed((&((8'ha1) ?
              (+(~(8'h9c))) : ((8'hba) ~^ $signed((8'ha3))))));
        end
      else
        begin
          for (forvar32 = (1'h0); (forvar32 < (3'h4)); forvar32 = (forvar32 + (1'h1)))
            begin
              reg33 <= ((8'hb7) >> $unsigned((("baK8CeDy3" ?
                  wire26[(2'h3):(1'h1)] : reg35) - "PIs")));
              reg34 <= (($unsigned("20YFNpwfzC57Naby8c") ~^ (forvar32[(2'h2):(1'h1)] ?
                  "Edo7Qh59cy4fNVd" : $signed((-(8'h9e))))) && (8'hbc));
              reg35 <= ((|(reg34[(3'h4):(3'h4)] * (8'ha5))) > reg32[(4'h8):(1'h1)]);
              reg36 <= $unsigned({$unsigned(($signed((8'h9e)) <= "3nKt89FXd8Py7pDlZc"))});
            end
          reg39 = reg31[(2'h2):(1'h0)];
          reg40 = ({"BWBTbPyxN", $unsigned($signed($signed((8'ha3))))} ?
              wire29 : $unsigned(wire26));
          reg41 <= $signed({(~^$unsigned({(8'hb8)})), forvar33});
        end
    end
  always
    @(posedge clk) begin
      reg42 <= (~^(wire29[(3'h7):(1'h0)] >> wire29));
      reg43 <= (7'h40);
      reg44 <= (8'hb8);
      reg45 <= (~|(({"x6Xb8PkD3"} ?
              (reg43 ?
                  $unsigned((7'h40)) : reg42[(3'h7):(1'h0)]) : (^~{(8'h9c)})) ?
          $unsigned((+$signed((8'h9e)))) : reg38[(1'h1):(1'h1)]));
      reg46 <= reg34[(1'h1):(1'h0)];
    end
  assign wire47 = {wire29[(3'h6):(3'h6)], (wire28[(2'h3):(1'h1)] > wire29)};
endmodule
