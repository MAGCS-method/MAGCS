(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param1471 = (+{(7'h43), ((^~((8'hb6) ? (8'hb5) : (8'ha9))) ~^ (((7'h46) ? (8'hbb) : (8'hb7)) >= ((8'hb9) - (8'hbd))))}))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h677):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire0;
  input wire [(5'h12):(1'h0)] wire1;
  input wire signed [(5'h15):(1'h0)] wire2;
  input wire signed [(4'hc):(1'h0)] wire3;
  input wire [(4'hc):(1'h0)] wire4;
  wire signed [(3'h5):(1'h0)] wire1451;
  wire [(5'h12):(1'h0)] wire54;
  wire signed [(5'h15):(1'h0)] wire55;
  wire signed [(3'h5):(1'h0)] wire56;
  wire signed [(4'hd):(1'h0)] wire103;
  wire [(4'hf):(1'h0)] wire104;
  wire signed [(4'hd):(1'h0)] wire190;
  wire signed [(4'hf):(1'h0)] wire1469;
  reg signed [(5'h17):(1'h0)] reg1468 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1467 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1466 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1462 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1461 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1460 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1459 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1458 = (1'h0);
  reg [(3'h6):(1'h0)] reg1457 = (1'h0);
  reg [(5'h14):(1'h0)] reg1456 = (1'h0);
  reg [(5'h16):(1'h0)] reg93 = (1'h0);
  reg [(3'h7):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg101 = (1'h0);
  reg [(4'he):(1'h0)] reg97 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg92 = (1'h0);
  reg [(5'h14):(1'h0)] reg90 = (1'h0);
  reg [(5'h11):(1'h0)] reg87 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg86 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg80 = (1'h0);
  reg [(4'hf):(1'h0)] reg75 = (1'h0);
  reg [(5'h11):(1'h0)] reg72 = (1'h0);
  reg [(3'h6):(1'h0)] reg69 = (1'h0);
  reg [(5'h17):(1'h0)] reg68 = (1'h0);
  reg signed [(4'he):(1'h0)] reg67 = (1'h0);
  reg [(4'hf):(1'h0)] reg65 = (1'h0);
  reg [(5'h14):(1'h0)] reg64 = (1'h0);
  reg [(5'h15):(1'h0)] reg53 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg51 = (1'h0);
  reg [(5'h12):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg49 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg48 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg44 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg39 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg37 = (1'h0);
  reg [(4'hf):(1'h0)] reg31 = (1'h0);
  reg [(3'h4):(1'h0)] reg30 = (1'h0);
  reg [(3'h7):(1'h0)] reg29 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg28 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg24 = (1'h0);
  reg [(4'hb):(1'h0)] reg20 = (1'h0);
  reg [(5'h14):(1'h0)] reg18 = (1'h0);
  reg [(5'h10):(1'h0)] reg15 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg14 = (1'h0);
  reg [(4'hc):(1'h0)] reg11 = (1'h0);
  reg [(5'h15):(1'h0)] reg8 = (1'h0);
  reg [(5'h15):(1'h0)] reg5 = (1'h0);
  reg [(5'h14):(1'h0)] reg1465 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1464 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1463 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1455 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1454 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1453 = (1'h0);
  reg [(5'h18):(1'h0)] forvar89 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg88 = (1'h0);
  reg [(3'h5):(1'h0)] forvar100 = (1'h0);
  reg [(5'h11):(1'h0)] reg99 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg98 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg95 = (1'h0);
  reg [(5'h10):(1'h0)] reg94 = (1'h0);
  reg [(4'hc):(1'h0)] forvar93 = (1'h0);
  reg [(2'h3):(1'h0)] reg91 = (1'h0);
  reg [(5'h12):(1'h0)] reg89 = (1'h0);
  reg [(4'hb):(1'h0)] forvar88 = (1'h0);
  reg signed [(4'he):(1'h0)] reg85 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar84 = (1'h0);
  reg [(4'he):(1'h0)] reg83 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg82 = (1'h0);
  reg [(4'hd):(1'h0)] reg81 = (1'h0);
  reg [(5'h11):(1'h0)] reg79 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar78 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg76 = (1'h0);
  reg [(4'ha):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg73 = (1'h0);
  reg [(4'h9):(1'h0)] reg71 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg70 = (1'h0);
  reg [(5'h11):(1'h0)] reg66 = (1'h0);
  reg [(5'h11):(1'h0)] reg63 = (1'h0);
  reg [(4'ha):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg61 = (1'h0);
  reg [(5'h17):(1'h0)] forvar60 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg [(5'h16):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar57 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar47 = (1'h0);
  reg [(4'hf):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg43 = (1'h0);
  reg [(5'h10):(1'h0)] reg41 = (1'h0);
  reg [(4'h9):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg38 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg36 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg35 = (1'h0);
  reg [(3'h7):(1'h0)] reg34 = (1'h0);
  reg [(5'h16):(1'h0)] reg33 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg32 = (1'h0);
  reg [(4'hd):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg26 = (1'h0);
  reg [(2'h3):(1'h0)] reg25 = (1'h0);
  reg [(4'hf):(1'h0)] reg23 = (1'h0);
  reg [(5'h15):(1'h0)] forvar22 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg21 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg16 = (1'h0);
  reg [(5'h14):(1'h0)] reg13 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg12 = (1'h0);
  reg [(5'h18):(1'h0)] forvar10 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg9 = (1'h0);
  reg [(5'h14):(1'h0)] reg7 = (1'h0);
  reg [(2'h2):(1'h0)] reg6 = (1'h0);
  assign y = {wire1451,
                 wire54,
                 wire55,
                 wire56,
                 wire103,
                 wire104,
                 wire190,
                 wire1469,
                 reg1468,
                 reg1467,
                 reg1466,
                 reg1462,
                 reg1461,
                 reg1460,
                 reg1459,
                 reg1458,
                 reg1457,
                 reg1456,
                 reg93,
                 reg102,
                 reg101,
                 reg97,
                 reg92,
                 reg90,
                 reg87,
                 reg86,
                 reg80,
                 reg75,
                 reg72,
                 reg69,
                 reg68,
                 reg67,
                 reg65,
                 reg64,
                 reg53,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg45,
                 reg44,
                 reg42,
                 reg39,
                 reg37,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg24,
                 reg20,
                 reg18,
                 reg15,
                 reg14,
                 reg11,
                 reg8,
                 reg5,
                 reg1465,
                 reg1464,
                 forvar1463,
                 reg1455,
                 reg1454,
                 forvar1453,
                 forvar89,
                 reg88,
                 forvar100,
                 reg99,
                 reg98,
                 reg96,
                 reg95,
                 reg94,
                 forvar93,
                 reg91,
                 reg89,
                 forvar88,
                 reg85,
                 forvar84,
                 reg83,
                 reg82,
                 reg81,
                 reg79,
                 forvar78,
                 reg77,
                 reg76,
                 reg74,
                 reg73,
                 reg71,
                 reg70,
                 reg66,
                 reg63,
                 reg62,
                 reg61,
                 forvar60,
                 reg59,
                 reg58,
                 forvar57,
                 reg52,
                 forvar47,
                 reg46,
                 reg43,
                 reg41,
                 reg40,
                 reg38,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg27,
                 reg26,
                 reg25,
                 reg23,
                 forvar22,
                 reg21,
                 reg19,
                 reg17,
                 reg16,
                 reg13,
                 reg12,
                 forvar10,
                 reg9,
                 reg7,
                 reg6,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg5 <= wire1;
      if ((reg5 != ((($signed(wire4) ?
              (wire0 != wire1) : wire0[(2'h2):(2'h2)]) ?
          wire4 : $unsigned((!reg5))) + $signed((wire0[(2'h2):(2'h2)] >= (wire4 == wire1))))))
        begin
          reg6 = $unsigned((-$unsigned(wire4)));
          reg7 = reg5;
        end
      else
        begin
          reg8 <= {$unsigned((^(reg5 < $unsigned(reg7)))), $unsigned(wire4)};
          reg9 = (&(!$signed(reg8)));
          for (forvar10 = (1'h0); (forvar10 < (2'h2)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg11 <= ((wire3 || ((|wire3[(1'h1):(1'h1)]) << reg9[(1'h0):(1'h0)])) ?
                  (-$unsigned(wire1)) : forvar10[(1'h0):(1'h0)]);
              reg12 = reg11;
              reg13 = {$signed($unsigned((!$unsigned(reg12)))),
                  ($signed($signed($signed(reg8))) - forvar10[(5'h15):(3'h4)])};
              reg14 <= $signed((|wire4));
            end
          if ($signed((reg14 ?
              $signed((!(reg9 << reg12))) : (({reg11} ?
                  $unsigned((8'hbd)) : (-wire0)) - ($signed(wire2) ?
                  wire4 : reg12)))))
            begin
              reg15 <= (^(({reg13} ?
                      (8'hb8) : (reg13[(1'h1):(1'h0)] ?
                          (8'ha0) : (reg9 ? reg14 : reg8))) ?
                  reg6 : (^~forvar10)));
            end
          else
            begin
              reg16 = (reg6 >= $signed((reg9 <= (wire1[(4'ha):(4'h9)] ?
                  $signed(wire2) : forvar10[(4'he):(4'he)]))));
            end
        end
      reg17 = ($signed(reg6) < {reg5[(3'h5):(1'h0)]});
      if ($signed(reg17[(4'hf):(1'h0)]))
        begin
          reg18 <= (reg8[(5'h10):(4'hd)] < ((((~wire3) >= (~reg7)) == $signed({reg17,
              forvar10})) ^ {$unsigned((+wire4))}));
          reg19 = $signed(reg6);
        end
      else
        begin
          if ($unsigned($signed($signed($unsigned($signed(reg6))))))
            begin
              reg19 = forvar10[(4'hf):(4'h9)];
            end
          else
            begin
              reg18 <= (((^$signed(wire3)) ? $unsigned((8'h9e)) : (-reg11)) ?
                  {reg16, reg6[(1'h0):(1'h0)]} : (reg7[(5'h11):(1'h1)] ?
                      (8'ha0) : {$signed((wire4 ? reg5 : reg14)),
                          forvar10[(4'h8):(2'h3)]}));
              reg20 <= (+(^$signed(reg16[(2'h3):(1'h1)])));
              reg21 = (((reg18[(5'h14):(3'h4)] >= ($unsigned(reg15) || $unsigned(reg7))) << wire2) ?
                  wire4[(4'hc):(4'h8)] : $signed((^~reg20)));
            end
          for (forvar22 = (1'h0); (forvar22 < (2'h2)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 = reg21;
              reg24 <= wire0[(2'h2):(2'h2)];
              reg25 = reg17;
            end
          reg26 = (~(reg12 ? reg17[(1'h0):(1'h0)] : (&(!$unsigned(reg16)))));
          reg27 = (reg20 ^~ ($unsigned(reg5[(4'h8):(3'h5)]) ?
              (((reg11 != reg9) <<< (wire3 + forvar22)) | ({reg6} >>> (reg9 <<< reg17))) : (!{reg7,
                  {reg25}})));
        end
      reg28 <= ((reg5 ?
          {reg18} : ({reg18} | $unsigned(wire4))) | ({forvar22[(3'h6):(1'h0)],
          (-(^reg27))} - {$signed((reg23 ? reg27 : reg25)),
          (forvar22[(4'hb):(4'h8)] ? (reg6 ? (8'hb8) : (8'hb3)) : reg25)}));
    end
  always
    @(posedge clk) begin
      reg29 <= (~|({(~&(wire2 & reg28))} <= $unsigned(wire0)));
      reg30 <= $signed(($unsigned(((reg5 <= wire2) <= (reg8 ? wire4 : reg29))) ?
          reg14 : reg18[(2'h2):(1'h1)]));
      if ($unsigned($signed(((&(wire3 || reg28)) || (wire0 + reg14)))))
        begin
          reg31 <= $signed(reg29);
          if (reg15[(4'hd):(2'h2)])
            begin
              reg32 = {$signed(reg30)};
              reg33 = $unsigned((|($signed((+wire2)) ?
                  reg15 : ((8'h9e) ? {wire1} : ((8'ha3) <= (8'hb6))))));
              reg34 = (reg11 >>> {reg30[(2'h3):(1'h0)],
                  $signed({$signed(reg32)})});
              reg35 = $unsigned(reg14);
              reg36 = ((|$signed($signed((reg11 ?
                  (8'haa) : reg18)))) & (|((((7'h47) & reg24) & {reg32}) ?
                  ((wire3 ?
                      reg32 : wire0) * reg18[(4'he):(2'h3)]) : (reg30 <<< $signed(reg31)))));
            end
          else
            begin
              reg37 <= (&reg33);
              reg38 = ($signed($signed(((~^reg37) <<< (reg34 >>> wire4)))) ?
                  $signed($signed($unsigned(reg37[(2'h2):(1'h0)]))) : ((reg35[(1'h0):(1'h0)] - $signed($unsigned(reg24))) ?
                      $signed(reg34) : {{(reg35 ? reg29 : reg5), (^~reg36)}}));
            end
        end
      else
        begin
          reg31 <= $unsigned($signed(reg18[(3'h5):(2'h3)]));
          if (reg11[(1'h0):(1'h0)])
            begin
              reg32 = (reg38[(4'hb):(4'ha)] ?
                  ((~^$unsigned(reg18[(4'he):(2'h3)])) <<< reg20[(1'h1):(1'h0)]) : reg32[(1'h1):(1'h0)]);
              reg33 = ({reg29} <<< $unsigned(({$signed((8'h9e)), reg33} ?
                  ((wire4 ^ wire1) ?
                      (reg38 | (8'hb0)) : $unsigned(reg34)) : ((+(8'had)) ?
                      (reg35 != reg34) : $unsigned(reg31)))));
              reg37 <= reg11[(4'h8):(3'h6)];
              reg39 <= $signed($signed(({(wire0 ? (8'h9d) : reg38)} ?
                  (~(^reg29)) : reg33[(3'h5):(3'h5)])));
            end
          else
            begin
              reg32 = reg24[(4'hf):(4'hb)];
              reg33 = reg24[(4'h9):(1'h1)];
            end
          if ($unsigned({($unsigned($unsigned(reg33)) <= (reg24 ^ reg37)),
              reg39[(4'ha):(3'h5)]}))
            begin
              reg40 = ($unsigned(reg37[(3'h6):(2'h2)]) ?
                  (((wire3 + (reg24 ^ reg28)) ? reg14 : (-(reg20 >> reg32))) ?
                      ((&$unsigned(reg34)) > $signed((reg18 <<< (8'hbb)))) : $signed(reg35[(4'hc):(4'h8)])) : $unsigned(reg18));
              reg41 = wire3[(4'ha):(3'h6)];
              reg42 <= reg29[(3'h7):(3'h7)];
              reg43 = $signed((reg5 && ((^(wire0 ?
                  reg11 : wire1)) | reg15[(4'hd):(4'ha)])));
              reg44 <= {(((wire0[(1'h0):(1'h0)] < (~^reg35)) ?
                      ((reg41 ?
                          reg35 : (7'h42)) | {reg29}) : reg30[(2'h3):(2'h3)]) <= $unsigned($unsigned((reg33 ?
                      reg15 : reg41)))),
                  $signed(reg40[(3'h6):(1'h0)])};
            end
          else
            begin
              reg42 <= {((((wire0 ? reg39 : reg42) ?
                      $unsigned(reg28) : $signed((7'h46))) || wire4[(3'h7):(3'h4)]) >>> (((reg43 ?
                              reg30 : reg43) ?
                          ((8'ha2) ? reg18 : reg36) : (reg24 ?
                              (8'hb5) : wire0)) ?
                      (^(reg41 ? (8'had) : wire3)) : (~^reg11)))};
              reg43 = ((-$unsigned(reg44[(3'h4):(2'h3)])) ?
                  reg30[(2'h2):(2'h2)] : (~&(7'h46)));
              reg44 <= wire4[(1'h1):(1'h0)];
              reg45 <= ((8'hbe) ? (+wire1[(1'h0):(1'h0)]) : (~^{{reg37}}));
            end
          reg46 = ({($unsigned($signed(wire0)) - (8'hbb)),
              $signed({(reg37 ? reg34 : reg11),
                  reg39[(3'h5):(1'h0)]})} | (^reg32));
          for (forvar47 = (1'h0); (forvar47 < (2'h2)); forvar47 = (forvar47 + (1'h1)))
            begin
              reg48 <= {((reg29[(3'h4):(1'h0)] ?
                          (&(reg32 ?
                              forvar47 : reg36)) : (reg24[(2'h3):(1'h0)] ?
                              $signed(wire3) : $unsigned(reg28))) ?
                      (wire3 | (reg34 ? wire2 : (~|reg39))) : (|wire2)),
                  (~({(~^reg11), $signed(reg43)} | $signed((~^reg45))))};
              reg49 <= ({$signed((^(reg20 ? reg34 : reg37))),
                      (((~reg15) ? (reg37 == reg5) : (~|reg36)) ?
                          $signed((reg33 ^~ reg48)) : reg38[(1'h0):(1'h0)])} ?
                  reg42 : ($signed(reg41[(4'h8):(3'h5)]) << (^~(!(reg11 ?
                      reg11 : (8'hbe))))));
              reg50 <= ($signed(reg32) ?
                  $signed($signed({$unsigned(reg39),
                      (reg24 ? reg45 : wire4)})) : (8'hb8));
              reg51 <= ((&$signed((~&$unsigned(reg18)))) > $signed($unsigned(((reg32 ?
                      reg5 : reg40) ?
                  (reg50 ^ (8'ha7)) : (reg11 << reg36)))));
            end
        end
      reg52 = ((~^reg20[(3'h4):(2'h2)]) && $unsigned($signed($signed($signed(reg43)))));
      reg53 <= (reg48 + ($signed({(^~reg28), (!reg31)}) <= reg31));
    end
  assign wire54 = wire1[(3'h6):(2'h3)];
  assign wire55 = (~&(8'ha1));
  assign wire56 = (wire4 >= {(reg48 ?
                          (^(reg50 ? reg42 : (8'hba))) : {$unsigned(reg11)})});
  always
    @(posedge clk) begin
      for (forvar57 = (1'h0); (forvar57 < (1'h1)); forvar57 = (forvar57 + (1'h1)))
        begin
          reg58 = $unsigned(($signed(reg49[(1'h1):(1'h0)]) ^ reg14[(1'h1):(1'h0)]));
          reg59 = wire2[(1'h1):(1'h0)];
          for (forvar60 = (1'h0); (forvar60 < (3'h4)); forvar60 = (forvar60 + (1'h1)))
            begin
              reg61 = ($unsigned(($signed(wire3) < wire56[(1'h1):(1'h0)])) ^ $unsigned((!$signed(wire55[(1'h1):(1'h0)]))));
              reg62 = wire4;
              reg63 = (8'hb4);
              reg64 <= reg53[(3'h6):(3'h6)];
              reg65 <= wire0;
            end
          if ($signed(reg5[(4'hc):(1'h0)]))
            begin
              reg66 = reg50;
            end
          else
            begin
              reg67 <= (~reg61);
              reg68 <= $unsigned(($signed((+(reg24 << reg20))) ?
                  (8'haf) : reg49[(4'he):(3'h4)]));
            end
          reg69 <= (&(reg24 ?
              $signed(wire4) : (reg39[(5'h12):(4'h9)] ~^ (~&reg58))));
        end
      if ((|$signed(wire4[(4'hc):(3'h4)])))
        begin
          reg70 = (reg50[(4'hf):(1'h1)] ^~ wire2);
        end
      else
        begin
          if (($signed({$unsigned(wire0[(1'h0):(1'h0)])}) ?
              $unsigned((8'hb2)) : {$signed($unsigned((reg53 ^ reg28)))}))
            begin
              reg70 = ((~wire55) ? (!reg29[(2'h3):(2'h3)]) : reg69);
              reg71 = reg44;
              reg72 <= reg59[(1'h1):(1'h1)];
              reg73 = $unsigned($signed(reg62));
              reg74 = ((|reg73[(3'h5):(1'h0)]) * (reg11 ?
                  reg68 : ({(^reg5)} ?
                      (!{reg44, reg59}) : $unsigned({reg45, reg58}))));
            end
          else
            begin
              reg72 <= wire54;
              reg75 <= $signed((^$signed(($signed((8'hba)) ?
                  $signed(reg65) : $signed(wire0)))));
              reg76 = $unsigned({$unsigned(reg68)});
              reg77 = {$signed($signed(((~&reg68) ?
                      $signed(reg70) : ((8'hbb) ^~ reg11)))),
                  reg67[(1'h1):(1'h0)]};
            end
          for (forvar78 = (1'h0); (forvar78 < (3'h4)); forvar78 = (forvar78 + (1'h1)))
            begin
              reg79 = $signed(({wire56, reg15[(1'h1):(1'h0)]} ^~ reg62));
              reg80 <= reg31;
              reg81 = forvar60[(3'h4):(2'h3)];
              reg82 = (-forvar60);
            end
        end
      reg83 = ($signed(((reg15[(3'h6):(1'h1)] ^~ $signed(reg77)) << (~$signed((7'h40))))) ?
          (&$unsigned($unsigned((reg8 <<< reg5)))) : reg50[(4'h8):(3'h7)]);
      for (forvar84 = (1'h0); (forvar84 < (2'h2)); forvar84 = (forvar84 + (1'h1)))
        begin
          reg85 = wire4[(4'hb):(4'ha)];
          reg86 <= (reg28[(3'h4):(3'h4)] ?
              reg85 : ((~^$unsigned(reg37)) ~^ (reg85 ?
                  ($signed(reg69) ?
                      {wire0, forvar60} : $unsigned(reg31)) : {((8'hb1) ?
                          reg53 : reg73)})));
          reg87 <= {(&$unsigned((reg18 ? (|reg31) : $signed(reg66)))),
              (reg18 ?
                  ($unsigned((reg79 ? reg70 : wire4)) ?
                      ($signed(reg81) + (&reg86)) : wire4[(4'ha):(3'h4)]) : $signed(reg45[(1'h1):(1'h0)]))};
        end
      if (reg85[(4'hb):(2'h3)])
        begin
          for (forvar88 = (1'h0); (forvar88 < (1'h1)); forvar88 = (forvar88 + (1'h1)))
            begin
              reg89 = (&reg63);
              reg90 <= reg83[(4'hb):(3'h5)];
              reg91 = (((reg68 ~^ ((reg67 ?
                  reg39 : (7'h40)) < reg15)) ^~ $unsigned((~reg64[(3'h6):(3'h4)]))) >>> (~^{reg71}));
            end
          reg92 <= reg69[(3'h5):(3'h5)];
          for (forvar93 = (1'h0); (forvar93 < (2'h2)); forvar93 = (forvar93 + (1'h1)))
            begin
              reg94 = ($signed((~&wire0[(2'h2):(1'h1)])) ?
                  (^~(~^$signed({reg15}))) : $unsigned({$signed($unsigned(reg11))}));
              reg95 = (reg51[(1'h1):(1'h1)] <<< forvar88);
              reg96 = (((((reg85 ? reg42 : reg5) > reg87[(3'h7):(3'h4)]) ?
                  reg58 : $unsigned($signed(reg89))) < (~^(((8'hae) ?
                      (8'had) : reg59) ?
                  (7'h46) : {wire4}))) <<< (~$signed(($signed(wire3) ?
                  reg91[(2'h3):(2'h2)] : reg69[(3'h6):(2'h2)]))));
              reg97 <= reg51;
              reg98 = reg8;
            end
          reg99 = (((($unsigned(reg80) ?
                      $signed(reg53) : (forvar78 ? forvar78 : reg77)) ?
                  $signed((|(8'hb5))) : reg81) * {(wire56 >>> {reg76,
                      (8'had)})}) ?
              ($signed($unsigned({reg37})) ?
                  (~^$signed((reg42 ?
                      wire54 : forvar84))) : $signed(((wire55 >= reg18) - (^~wire0)))) : $unsigned(reg31));
          for (forvar100 = (1'h0); (forvar100 < (1'h0)); forvar100 = (forvar100 + (1'h1)))
            begin
              reg101 <= $unsigned(reg81);
              reg102 <= ($unsigned(reg5) ?
                  reg81[(4'hd):(4'hb)] : forvar88[(2'h3):(1'h0)]);
            end
        end
      else
        begin
          reg88 = ((~&{reg53[(3'h7):(3'h6)],
              {reg68[(5'h17):(4'h8)]}}) >= reg96[(3'h5):(1'h0)]);
          for (forvar89 = (1'h0); (forvar89 < (1'h0)); forvar89 = (forvar89 + (1'h1)))
            begin
              reg90 <= (^forvar93[(4'h9):(4'h9)]);
              reg91 = (~reg92[(1'h1):(1'h1)]);
              reg92 <= {(reg39 ? {wire4, $unsigned((~|reg59))} : reg14)};
              reg93 <= wire54;
            end
          reg97 <= ($signed({($signed(reg95) ?
                  reg68[(1'h1):(1'h0)] : reg62[(3'h4):(3'h4)])}) | reg20[(1'h1):(1'h0)]);
        end
    end
  assign wire103 = ({$signed(reg8[(5'h11):(4'h8)])} ?
                       $signed({(|wire55[(1'h1):(1'h0)]),
                           ((reg64 << reg14) ?
                               $unsigned(reg93) : ((8'haf) - (8'hbd)))}) : {(~&(!(reg29 ?
                               reg67 : reg102)))});
  assign wire104 = wire55[(5'h12):(4'h8)];
  module105 #() modinst191 (.wire110(reg44), .clk(clk), .wire106(reg68), .wire108(reg69), .wire109(wire56), .wire107(reg75), .y(wire190));
  module192 #() modinst1452 (wire1451, clk, wire0, reg53, reg5, reg44, reg49);
  always
    @(posedge clk) begin
      for (forvar1453 = (1'h0); (forvar1453 < (1'h1)); forvar1453 = (forvar1453 + (1'h1)))
        begin
          if (wire103[(4'hb):(3'h7)])
            begin
              reg1454 = wire4[(1'h1):(1'h1)];
              reg1455 = {wire3};
              reg1456 <= ($unsigned((-$unsigned((reg49 != reg42)))) + reg53);
              reg1457 <= (((reg42[(1'h1):(1'h0)] ?
                      $signed((~^wire54)) : reg18) ^ $unsigned($unsigned(wire54[(3'h6):(1'h1)]))) ?
                  ((!$signed(reg48[(1'h0):(1'h0)])) == reg15) : $signed((reg102[(3'h7):(3'h6)] ?
                      ({wire1451, (8'hb8)} ?
                          wire55 : reg11[(4'hc):(4'h8)]) : ($unsigned(reg20) ?
                          $signed(reg64) : $unsigned(reg53)))));
            end
          else
            begin
              reg1454 = reg72[(2'h3):(2'h2)];
              reg1455 = ((-reg45) ?
                  reg101[(4'h8):(2'h3)] : (reg8 <= $unsigned(((reg65 != reg101) ?
                      (+reg48) : reg28))));
              reg1456 <= reg31[(2'h3):(2'h3)];
              reg1457 <= (&$signed((~|($signed((7'h45)) ?
                  $unsigned(wire54) : {wire190, reg50}))));
              reg1458 <= {($unsigned(reg49[(4'hb):(4'ha)]) ?
                      ((!$unsigned(reg69)) << $signed($signed(reg24))) : wire3)};
            end
          if (reg1458)
            begin
              reg1459 <= $unsigned(($signed(((^~reg15) * $unsigned(reg37))) ?
                  $signed(wire54) : $unsigned({(~&wire1451),
                      (wire55 & reg75)})));
              reg1460 <= $unsigned((((8'hb7) ?
                      (+reg5) : reg1459[(3'h6):(3'h4)]) ?
                  (|$unsigned((-reg51))) : reg20));
              reg1461 <= $signed({reg39[(4'h8):(3'h6)]});
              reg1462 <= ((~|wire1) != ($unsigned($signed((^~reg8))) ?
                  ($signed(reg14) >>> {$signed(wire1)}) : reg11[(4'ha):(1'h1)]));
            end
          else
            begin
              reg1459 <= reg1455;
            end
          for (forvar1463 = (1'h0); (forvar1463 < (1'h0)); forvar1463 = (forvar1463 + (1'h1)))
            begin
              reg1464 = (reg45[(1'h1):(1'h1)] ?
                  reg1462 : (reg93 ?
                      $unsigned($signed((~|reg1457))) : (&$signed($signed(reg24)))));
            end
          reg1465 = $signed((($unsigned({reg1464}) ?
                  $unsigned((wire56 | reg29)) : reg1461[(4'h9):(3'h4)]) ?
              reg69 : (^((wire2 ^~ wire0) ?
                  $signed(reg24) : (wire104 ? reg101 : reg18)))));
        end
      reg1466 <= (($unsigned($unsigned((reg14 ? reg30 : (7'h47)))) ?
          $unsigned($signed((~|reg75))) : ($unsigned((reg51 ?
              wire190 : reg68)) - reg1457)) << $signed($signed($unsigned((&wire104)))));
      reg1467 <= (reg8 ? wire3 : reg67);
      reg1468 <= $unsigned(reg92);
    end
  module619 #() modinst1470 (.wire623(reg24), .wire624(reg1460), .clk(clk), .wire622(reg80), .y(wire1469), .wire621(wire54), .wire620(reg93));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module192
#(parameter param1449 = (8'hbb), 
parameter param1450 = (^{((~&(param1449 ~^ param1449)) ? (~(~^param1449)) : (((8'hb7) != param1449) ? (~^(7'h45)) : param1449))}))
(y, clk, wire193, wire194, wire195, wire196, wire197);
  output wire [(32'h368):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire193;
  input wire [(5'h15):(1'h0)] wire194;
  input wire [(5'h14):(1'h0)] wire195;
  input wire [(5'h18):(1'h0)] wire196;
  input wire [(5'h14):(1'h0)] wire197;
  wire signed [(5'h12):(1'h0)] wire1448;
  wire [(2'h2):(1'h0)] wire1447;
  wire [(3'h6):(1'h0)] wire1406;
  wire [(5'h16):(1'h0)] wire198;
  wire signed [(5'h18):(1'h0)] wire199;
  wire [(2'h2):(1'h0)] wire1381;
  reg signed [(4'he):(1'h0)] reg1446 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1445 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1444 = (1'h0);
  reg [(5'h15):(1'h0)] reg1442 = (1'h0);
  reg [(4'hf):(1'h0)] reg1440 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1439 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1438 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1433 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1431 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1430 = (1'h0);
  reg [(5'h11):(1'h0)] reg1429 = (1'h0);
  reg [(3'h7):(1'h0)] reg1428 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1426 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1425 = (1'h0);
  reg [(4'hc):(1'h0)] reg1423 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1417 = (1'h0);
  reg [(2'h2):(1'h0)] reg1416 = (1'h0);
  reg [(4'ha):(1'h0)] reg1414 = (1'h0);
  reg [(4'hc):(1'h0)] reg1411 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1409 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1404 = (1'h0);
  reg [(4'ha):(1'h0)] reg1400 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1394 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1390 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1389 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1385 = (1'h0);
  reg [(5'h13):(1'h0)] reg1443 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1441 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1439 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1437 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1436 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1435 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1434 = (1'h0);
  reg [(5'h12):(1'h0)] reg1432 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1427 = (1'h0);
  reg [(4'hf):(1'h0)] reg1424 = (1'h0);
  reg [(5'h13):(1'h0)] reg1422 = (1'h0);
  reg [(4'h9):(1'h0)] reg1421 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1420 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1419 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1418 = (1'h0);
  reg [(3'h5):(1'h0)] reg1415 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1413 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1412 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1410 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1408 = (1'h0);
  reg [(5'h16):(1'h0)] reg1407 = (1'h0);
  reg [(4'hd):(1'h0)] reg1405 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1403 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1402 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1401 = (1'h0);
  reg [(3'h6):(1'h0)] reg1399 = (1'h0);
  reg [(4'ha):(1'h0)] reg1398 = (1'h0);
  reg [(2'h3):(1'h0)] reg1397 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1396 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1395 = (1'h0);
  reg [(5'h14):(1'h0)] reg1393 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1392 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1391 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1388 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1387 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1386 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1384 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1383 = (1'h0);
  assign y = {wire1448,
                 wire1447,
                 wire1406,
                 wire198,
                 wire199,
                 wire1381,
                 reg1446,
                 reg1445,
                 reg1444,
                 reg1442,
                 reg1440,
                 reg1439,
                 reg1438,
                 reg1433,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1426,
                 reg1425,
                 reg1423,
                 reg1417,
                 reg1416,
                 reg1414,
                 reg1411,
                 reg1409,
                 reg1404,
                 reg1400,
                 reg1394,
                 reg1390,
                 reg1389,
                 reg1385,
                 reg1443,
                 reg1441,
                 forvar1439,
                 reg1437,
                 reg1436,
                 reg1435,
                 reg1434,
                 reg1432,
                 reg1427,
                 reg1424,
                 reg1422,
                 reg1421,
                 forvar1420,
                 reg1419,
                 reg1418,
                 reg1415,
                 forvar1413,
                 forvar1412,
                 reg1410,
                 forvar1408,
                 reg1407,
                 reg1405,
                 forvar1403,
                 reg1402,
                 reg1401,
                 reg1399,
                 reg1398,
                 reg1397,
                 forvar1396,
                 forvar1395,
                 reg1393,
                 reg1392,
                 reg1391,
                 forvar1388,
                 reg1387,
                 reg1386,
                 forvar1384,
                 forvar1383,
                 (1'h0)};
  assign wire198 = $signed($unsigned($signed((wire193 == wire193))));
  assign wire199 = (-$signed((^~$signed((^~wire195)))));
  module200 #() modinst1382 (.wire204(wire195), .wire202(wire193), .y(wire1381), .wire203(wire199), .wire205(wire194), .clk(clk), .wire201(wire197));
  always
    @(posedge clk) begin
      for (forvar1383 = (1'h0); (forvar1383 < (2'h2)); forvar1383 = (forvar1383 + (1'h1)))
        begin
          for (forvar1384 = (1'h0); (forvar1384 < (1'h0)); forvar1384 = (forvar1384 + (1'h1)))
            begin
              reg1385 <= (~wire1381);
              reg1386 = ($signed((wire193[(4'h9):(4'h9)] <<< $unsigned((+reg1385)))) ?
                  (((~&((8'hb7) >>> reg1385)) ~^ wire193) <= (forvar1384[(3'h7):(1'h0)] ?
                      wire195[(4'ha):(2'h3)] : wire198[(5'h15):(2'h3)])) : wire1381[(2'h2):(2'h2)]);
            end
          reg1387 = reg1385[(3'h5):(3'h5)];
          for (forvar1388 = (1'h0); (forvar1388 < (1'h0)); forvar1388 = (forvar1388 + (1'h1)))
            begin
              reg1389 <= (^$signed(wire198));
              reg1390 <= $unsigned((~|$unsigned(wire195[(5'h14):(5'h10)])));
              reg1391 = {$unsigned(wire1381),
                  (((~^{forvar1384, forvar1388}) ?
                      (|$unsigned(reg1385)) : {reg1389,
                          (wire1381 ? wire196 : reg1385)}) < forvar1384)};
              reg1392 = (~|reg1385);
            end
          reg1393 = wire195;
          reg1394 <= reg1385[(5'h10):(3'h7)];
        end
      for (forvar1395 = (1'h0); (forvar1395 < (3'h4)); forvar1395 = (forvar1395 + (1'h1)))
        begin
          for (forvar1396 = (1'h0); (forvar1396 < (3'h4)); forvar1396 = (forvar1396 + (1'h1)))
            begin
              reg1397 = (&(wire1381 ?
                  $signed(((~|forvar1388) >= (&(8'hb4)))) : wire196));
              reg1398 = forvar1383;
              reg1399 = (+(wire199 ?
                  wire198[(5'h11):(3'h5)] : reg1393[(4'hd):(4'hb)]));
              reg1400 <= {$signed(wire195), reg1389};
              reg1401 = reg1398;
            end
          reg1402 = $signed(({((forvar1388 ?
                  forvar1395 : reg1392) <<< (forvar1396 ?
                  wire196 : reg1391))} <= (&$signed(((8'ha6) >= wire195)))));
        end
      for (forvar1403 = (1'h0); (forvar1403 < (2'h3)); forvar1403 = (forvar1403 + (1'h1)))
        begin
          if ((8'ha1))
            begin
              reg1404 <= (|(~&(~|{$unsigned(wire196)})));
            end
          else
            begin
              reg1404 <= $signed(forvar1383);
            end
          reg1405 = (+wire1381);
        end
    end
  assign wire1406 = ((reg1390[(3'h7):(2'h2)] ?
                            {(~&reg1400[(3'h6):(1'h0)])} : reg1385[(5'h10):(3'h5)]) ?
                        $signed((|reg1385)) : $unsigned($unsigned((((8'ha8) ?
                                reg1390 : wire197) ?
                            wire193 : {wire1381}))));
  always
    @(posedge clk) begin
      if ((~&($signed(wire1381) * (^~wire197))))
        begin
          reg1407 = reg1394[(4'h9):(3'h7)];
          for (forvar1408 = (1'h0); (forvar1408 < (1'h0)); forvar1408 = (forvar1408 + (1'h1)))
            begin
              reg1409 <= $signed($unsigned($unsigned($unsigned($unsigned(reg1400)))));
              reg1410 = (8'hb7);
            end
        end
      else
        begin
          reg1407 = reg1389[(5'h11):(4'h8)];
        end
      reg1411 <= $unsigned({reg1407});
      for (forvar1412 = (1'h0); (forvar1412 < (1'h0)); forvar1412 = (forvar1412 + (1'h1)))
        begin
          for (forvar1413 = (1'h0); (forvar1413 < (2'h3)); forvar1413 = (forvar1413 + (1'h1)))
            begin
              reg1414 <= $unsigned((8'h9e));
              reg1415 = reg1411[(4'hb):(1'h0)];
              reg1416 <= forvar1412;
              reg1417 <= reg1414[(2'h3):(1'h1)];
              reg1418 = ($unsigned({forvar1413}) ?
                  reg1389[(4'hc):(3'h7)] : reg1394[(2'h2):(1'h0)]);
            end
          reg1419 = reg1385;
        end
      for (forvar1420 = (1'h0); (forvar1420 < (2'h3)); forvar1420 = (forvar1420 + (1'h1)))
        begin
          reg1421 = $signed($signed(forvar1412));
          if ($signed(wire193))
            begin
              reg1422 = (-(-{$signed((reg1407 ? reg1416 : reg1400))}));
              reg1423 <= (-reg1422);
              reg1424 = (^(^wire194[(4'he):(2'h2)]));
            end
          else
            begin
              reg1423 <= $unsigned(forvar1420);
              reg1424 = reg1410[(1'h0):(1'h0)];
              reg1425 <= (8'hb2);
            end
        end
      reg1426 <= ((~({reg1404[(2'h2):(1'h0)], $signed(reg1421)} ?
          reg1404 : $unsigned((!reg1390)))) >= $signed($signed(wire193)));
    end
  always
    @(posedge clk) begin
      reg1427 = $unsigned(reg1394);
      reg1428 <= $unsigned(reg1385[(1'h1):(1'h1)]);
      if (wire1406[(1'h1):(1'h1)])
        begin
          reg1429 <= ((wire195 >= ((~|$signed(wire195)) ?
                  wire199 : $signed((~|reg1385)))) ?
              (+(reg1416 * ((~|reg1409) >> $signed(reg1423)))) : {$unsigned({$unsigned(reg1409)}),
                  $unsigned(wire195[(4'hd):(3'h6)])});
          if ({(reg1389[(4'he):(1'h0)] - $signed(((wire197 ?
                      (8'hb4) : wire1381) ?
                  wire196[(4'hd):(3'h6)] : wire196[(5'h15):(5'h10)])))})
            begin
              reg1430 <= ((reg1423 < wire194[(5'h11):(3'h7)]) ?
                  $unsigned(reg1409) : $unsigned(((reg1428[(2'h3):(1'h1)] ?
                      (reg1416 ?
                          wire199 : reg1400) : $unsigned(reg1429)) * (^{reg1423,
                      reg1423}))));
              reg1431 <= (8'hae);
              reg1432 = {$signed($unsigned(reg1389[(3'h4):(2'h3)])),
                  ({((reg1426 > reg1430) >>> $signed(reg1390))} != reg1417)};
              reg1433 <= $unsigned((~&{reg1430}));
            end
          else
            begin
              reg1432 = (&(~|$signed({{reg1425, reg1433},
                  wire199[(5'h17):(2'h2)]})));
              reg1434 = $signed((reg1417[(4'ha):(4'ha)] ?
                  wire199 : ($unsigned(reg1390[(2'h2):(2'h2)]) + wire199)));
              reg1435 = $unsigned((8'h9d));
              reg1436 = $signed($unsigned((($signed(reg1417) ?
                      reg1390 : (&reg1400)) ?
                  (&(~^wire196)) : reg1414)));
              reg1437 = {reg1428[(3'h6):(3'h6)]};
            end
          reg1438 <= wire196;
        end
      else
        begin
          reg1432 = reg1435;
        end
      if (((((8'ha6) ? $signed(reg1432[(3'h4):(1'h1)]) : {$signed(reg1385)}) ?
              $unsigned(({wire197} ?
                  $unsigned((8'hb9)) : (reg1437 + reg1436))) : $signed({(reg1435 ?
                      (8'hb5) : (8'ha6))})) ?
          $unsigned(wire198) : (wire194 ?
              {{(&wire195)}} : ((^(reg1389 * reg1436)) ?
                  reg1436 : $signed(reg1435[(5'h10):(1'h0)])))))
        begin
          reg1439 <= ({reg1434[(1'h0):(1'h0)]} ?
              $unsigned((7'h42)) : $signed(reg1434[(1'h1):(1'h1)]));
          reg1440 <= (!(-($unsigned(((8'ha3) ?
              reg1400 : wire194)) >>> (~&$unsigned(wire198)))));
        end
      else
        begin
          for (forvar1439 = (1'h0); (forvar1439 < (2'h2)); forvar1439 = (forvar1439 + (1'h1)))
            begin
              reg1441 = {$signed(((wire1381[(2'h2):(2'h2)] & (-forvar1439)) || (&$unsigned(reg1400)))),
                  $signed(((+((7'h48) && reg1436)) >> reg1429[(1'h1):(1'h0)]))};
              reg1442 <= reg1438;
              reg1443 = $unsigned($signed(reg1390));
              reg1444 <= $unsigned(reg1417);
            end
          reg1445 <= reg1443;
        end
      reg1446 <= $unsigned($unsigned((+(reg1433 || (wire197 ?
          wire194 : reg1438)))));
    end
  assign wire1447 = $unsigned(((((reg1425 ?
                            wire199 : reg1442) * wire1406[(3'h4):(1'h0)]) >>> $signed(wire194[(4'hd):(3'h7)])) ?
                        reg1400 : ($signed($unsigned(reg1440)) ?
                            reg1446[(3'h5):(1'h1)] : {reg1439[(5'h10):(4'ha)],
                                (7'h45)})));
  assign wire1448 = (~&reg1440);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module105
#(parameter param188 = ((^((^~{(8'hae), (8'hb2)}) <= (((7'h43) ? (8'ha7) : (8'hb8)) ? ((8'ha5) ? (8'hbf) : (8'hbd)) : {(8'haa), (8'hb2)}))) << (((|((8'h9c) || (8'haf))) >> (~^((7'h4a) & (8'hac)))) ? ((((8'had) ? (8'hb8) : (8'hbe)) || (^(8'hb5))) ? (((8'ha6) ? (8'had) : (8'hb4)) ? (^(7'h46)) : ((8'hb3) ? (8'hab) : (8'hbd))) : ({(7'h47)} < ((8'hb2) && (8'ha1)))) : ((&{(7'h43)}) ? (((8'hb6) * (8'hae)) ? ((8'ha6) ? (7'h42) : (8'ha7)) : (~&(7'h41))) : (((8'ha0) >= (7'h49)) >= ((7'h47) ? (7'h43) : (7'h42)))))), 
parameter param189 = (((~|param188) && ((((8'ha3) ? (8'hb5) : param188) ? param188 : param188) ? ((~&param188) ? (|param188) : (~(8'ha2))) : ((~^param188) ? ((7'h42) + param188) : (~&param188)))) ? (((8'hac) ? ({param188} ^ (param188 <= param188)) : param188) ? ((^~(param188 >= param188)) + (~(^~param188))) : (({param188} || (param188 && param188)) | param188)) : (8'hbd)))
(y, clk, wire110, wire109, wire108, wire107, wire106);
  output wire [(32'h40d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire110;
  input wire signed [(2'h2):(1'h0)] wire109;
  input wire signed [(2'h3):(1'h0)] wire108;
  input wire [(4'hf):(1'h0)] wire107;
  input wire signed [(4'hf):(1'h0)] wire106;
  wire [(4'hb):(1'h0)] wire187;
  wire signed [(4'h9):(1'h0)] wire185;
  reg [(3'h5):(1'h0)] reg186 = (1'h0);
  reg [(5'h17):(1'h0)] reg184 = (1'h0);
  reg [(4'h8):(1'h0)] reg180 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg179 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg176 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg174 = (1'h0);
  reg [(4'h9):(1'h0)] reg172 = (1'h0);
  reg [(5'h15):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg166 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg157 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg154 = (1'h0);
  reg [(4'hf):(1'h0)] reg152 = (1'h0);
  reg [(4'h8):(1'h0)] reg138 = (1'h0);
  reg [(4'ha):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg148 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg145 = (1'h0);
  reg [(4'h9):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg141 = (1'h0);
  reg [(5'h10):(1'h0)] reg139 = (1'h0);
  reg [(5'h12):(1'h0)] reg135 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg134 = (1'h0);
  reg [(2'h3):(1'h0)] reg130 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg129 = (1'h0);
  reg [(5'h18):(1'h0)] reg126 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg124 = (1'h0);
  reg [(4'hb):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg117 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg114 = (1'h0);
  reg [(3'h6):(1'h0)] reg113 = (1'h0);
  reg [(3'h6):(1'h0)] forvar183 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg181 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar178 = (1'h0);
  reg [(5'h18):(1'h0)] reg177 = (1'h0);
  reg [(3'h7):(1'h0)] reg175 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar173 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar171 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg170 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg169 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar167 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg165 = (1'h0);
  reg [(5'h10):(1'h0)] forvar164 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar163 = (1'h0);
  reg [(4'h8):(1'h0)] reg162 = (1'h0);
  reg [(2'h3):(1'h0)] reg161 = (1'h0);
  reg [(5'h17):(1'h0)] reg160 = (1'h0);
  reg [(5'h17):(1'h0)] reg158 = (1'h0);
  reg [(5'h18):(1'h0)] reg156 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar155 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg153 = (1'h0);
  reg [(4'hf):(1'h0)] forvar151 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar141 = (1'h0);
  reg [(3'h7):(1'h0)] reg149 = (1'h0);
  reg [(4'hf):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg144 = (1'h0);
  reg [(5'h17):(1'h0)] reg143 = (1'h0);
  reg [(5'h15):(1'h0)] reg140 = (1'h0);
  reg [(4'hd):(1'h0)] forvar138 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg137 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg136 = (1'h0);
  reg [(4'hd):(1'h0)] reg133 = (1'h0);
  reg signed [(4'he):(1'h0)] reg132 = (1'h0);
  reg [(3'h4):(1'h0)] reg131 = (1'h0);
  reg [(5'h17):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar119 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg121 = (1'h0);
  reg [(4'he):(1'h0)] reg120 = (1'h0);
  reg [(4'ha):(1'h0)] reg119 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg116 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar112 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar111 = (1'h0);
  assign y = {wire187,
                 wire185,
                 reg186,
                 reg184,
                 reg180,
                 reg179,
                 reg176,
                 reg174,
                 reg172,
                 reg168,
                 reg166,
                 reg159,
                 reg157,
                 reg154,
                 reg152,
                 reg138,
                 reg150,
                 reg148,
                 reg145,
                 reg142,
                 reg141,
                 reg139,
                 reg135,
                 reg134,
                 reg130,
                 reg129,
                 reg126,
                 reg124,
                 reg123,
                 reg117,
                 reg114,
                 reg113,
                 forvar183,
                 reg182,
                 reg181,
                 forvar178,
                 reg177,
                 reg175,
                 forvar173,
                 forvar171,
                 reg170,
                 reg169,
                 forvar167,
                 reg165,
                 forvar164,
                 forvar163,
                 reg162,
                 reg161,
                 reg160,
                 reg158,
                 reg156,
                 forvar155,
                 reg153,
                 forvar151,
                 forvar141,
                 reg149,
                 reg147,
                 reg146,
                 reg144,
                 reg143,
                 reg140,
                 forvar138,
                 reg137,
                 reg136,
                 reg133,
                 reg132,
                 reg131,
                 reg128,
                 reg127,
                 forvar119,
                 reg125,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg116,
                 reg115,
                 forvar112,
                 forvar111,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar111 = (1'h0); (forvar111 < (3'h4)); forvar111 = (forvar111 + (1'h1)))
        begin
          for (forvar112 = (1'h0); (forvar112 < (2'h3)); forvar112 = (forvar112 + (1'h1)))
            begin
              reg113 <= wire106[(4'hc):(2'h3)];
              reg114 <= wire107;
              reg115 = wire110[(4'h9):(4'h9)];
            end
          if ($unsigned($unsigned((&wire107[(1'h1):(1'h0)]))))
            begin
              reg116 = (~$signed(((~^(!forvar112)) < (!$unsigned(wire109)))));
            end
          else
            begin
              reg117 <= ((|$signed($unsigned($unsigned(reg116)))) ^~ (!$unsigned($signed(wire109[(1'h1):(1'h1)]))));
            end
          reg118 = ($signed(reg115[(2'h3):(1'h1)]) ^ {forvar111[(2'h3):(1'h0)]});
        end
      if ($unsigned((((~&reg116) ?
              (wire107 ?
                  wire109[(2'h2):(1'h1)] : (wire109 ?
                      forvar112 : (8'hbd))) : {(reg115 & wire107)}) ?
          (wire108[(1'h0):(1'h0)] >> (wire107[(4'hd):(4'h9)] ?
              forvar111 : $unsigned(wire106))) : {wire108,
              $signed((reg113 >>> wire110))})))
        begin
          if ($unsigned(wire110[(3'h6):(3'h5)]))
            begin
              reg119 = ($unsigned($unsigned({reg113[(1'h0):(1'h0)]})) ?
                  $unsigned((-(reg114 ?
                      reg117 : reg113))) : $signed(forvar111[(1'h0):(1'h0)]));
              reg120 = (wire110[(3'h7):(3'h7)] ?
                  (reg114[(4'ha):(3'h4)] ~^ forvar112) : (8'hae));
              reg121 = wire106;
              reg122 = reg118;
              reg123 <= ({$signed($signed($unsigned(reg113))),
                  (reg117 ?
                      reg115 : (~|(reg121 ? reg116 : (7'h46))))} << reg120);
            end
          else
            begin
              reg119 = $signed(wire109);
              reg123 <= (($signed((wire109 ? reg115 : reg119[(2'h2):(1'h1)])) ?
                  reg119[(3'h7):(2'h2)] : {reg113[(3'h4):(1'h0)]}) & (|reg121));
              reg124 <= (~wire106);
              reg125 = reg116;
              reg126 <= reg115[(3'h7):(1'h1)];
            end
        end
      else
        begin
          for (forvar119 = (1'h0); (forvar119 < (2'h3)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg123 <= $unsigned($unsigned(((reg121 <= (~&reg114)) ?
                  wire109 : $unsigned((wire106 <<< reg123)))));
            end
          if ($unsigned(({$unsigned((reg126 != wire109)),
                  (~&reg120[(2'h3):(2'h3)])} ?
              ($unsigned((7'h44)) ^~ reg120[(4'ha):(3'h5)]) : ($signed((+(8'had))) ^~ forvar111[(3'h4):(3'h4)]))))
            begin
              reg125 = $signed(forvar119);
              reg126 <= forvar111[(2'h3):(1'h0)];
              reg127 = (^~$unsigned(($signed({forvar112}) ~^ (reg120[(4'hd):(4'h9)] < ((7'h43) >> reg125)))));
            end
          else
            begin
              reg124 <= $unsigned($unsigned(reg122));
              reg125 = (|(reg121 ? reg123 : forvar119));
              reg127 = {$signed((8'hbb)),
                  ($unsigned(reg114) ?
                      ({(wire106 ? wire110 : forvar119)} ?
                          $signed((+reg113)) : reg126[(3'h6):(3'h4)]) : forvar119)};
              reg128 = $unsigned(reg127[(4'hc):(3'h6)]);
              reg129 <= reg122;
            end
          if (wire110[(4'hb):(4'ha)])
            begin
              reg130 <= (^$unsigned(reg114[(3'h6):(2'h2)]));
            end
          else
            begin
              reg130 <= $signed(reg122[(1'h0):(1'h0)]);
              reg131 = ((!$unsigned({(!wire107), forvar119[(4'hb):(4'ha)]})) ?
                  $unsigned($signed(reg115)) : ($signed(reg124[(4'h8):(2'h2)]) << ((7'h46) ?
                      reg123 : $unsigned((forvar119 != wire108)))));
              reg132 = ($unsigned((~&((wire109 ~^ forvar111) ?
                  (reg128 >> reg116) : (forvar119 && wire109)))) <= {(reg119[(4'h8):(2'h2)] <= (^~reg119[(1'h0):(1'h0)]))});
              reg133 = wire110[(2'h2):(1'h1)];
            end
          reg134 <= forvar112[(4'ha):(3'h4)];
          reg135 <= $signed($unsigned(reg122));
        end
      reg136 = (~wire110);
      if (((!$unsigned($unsigned({reg114,
          reg113}))) == $unsigned((~^(!((8'ha7) ? (8'ha5) : wire106))))))
        begin
          reg137 = {$unsigned($signed((~^forvar111)))};
          for (forvar138 = (1'h0); (forvar138 < (2'h3)); forvar138 = (forvar138 + (1'h1)))
            begin
              reg139 <= reg124;
              reg140 = reg129[(3'h5):(2'h3)];
            end
          if (((~{((7'h44) * $signed(reg120)), wire108[(2'h2):(1'h0)]}) ?
              $signed(reg124[(1'h1):(1'h0)]) : (((~&$signed(reg114)) * ((reg122 >>> (8'ha9)) ?
                      (^~forvar111) : {(8'hb1)})) ?
                  reg139[(2'h3):(1'h0)] : (!($signed(forvar111) ?
                      (reg132 ? forvar111 : wire109) : ((8'ha2) ~^ wire110))))))
            begin
              reg141 <= (&(+reg133));
              reg142 <= ((8'ha3) | $signed(reg113));
              reg143 = $unsigned(($signed(reg119[(4'ha):(3'h4)]) ?
                  (&((8'hbb) ?
                      (reg127 ?
                          reg129 : wire109) : (reg130 == reg140))) : (((~reg136) ^~ $unsigned(reg129)) ?
                      (8'haf) : reg142)));
              reg144 = reg117[(5'h13):(4'hc)];
            end
          else
            begin
              reg143 = (~^((~&$signed($unsigned(reg133))) ?
                  $signed((~|(reg123 << forvar138))) : $signed($signed($unsigned(reg130)))));
              reg144 = $signed({($unsigned($unsigned(reg129)) ?
                      $unsigned((reg136 <= wire106)) : ({reg136, (8'hb9)} ?
                          {reg131} : $signed(reg128)))});
              reg145 <= $signed({{($unsigned(reg124) ?
                          reg128[(5'h14):(3'h5)] : {forvar119, reg136})},
                  reg119[(4'h8):(3'h5)]});
              reg146 = reg134[(2'h2):(1'h1)];
            end
          if ((!(forvar111[(2'h3):(2'h2)] ?
              (^~reg117[(3'h5):(3'h4)]) : $unsigned(($signed(reg122) >> ((7'h45) != reg131))))))
            begin
              reg147 = ({{(^((8'ha1) ? reg136 : reg128)),
                      ({wire110} ?
                          (reg136 ?
                              wire110 : (8'hb5)) : reg146[(4'hc):(2'h2)])},
                  {$signed(reg144[(1'h1):(1'h0)])}} != reg114[(1'h0):(1'h0)]);
              reg148 <= (~^(($unsigned(((8'hb7) >> reg116)) >> reg145[(1'h1):(1'h1)]) ?
                  (~^(forvar119[(4'hc):(1'h1)] * $unsigned(reg139))) : $signed((reg133 ?
                      reg135 : reg144))));
              reg149 = (-((-(-(^~reg134))) ?
                  $unsigned((~|(wire109 ?
                      (8'ha9) : reg128))) : $signed(((+reg113) & $signed(reg147)))));
            end
          else
            begin
              reg147 = $signed(reg114[(3'h5):(3'h4)]);
              reg148 <= reg127;
              reg149 = $signed(((reg135[(2'h2):(1'h1)] ?
                      $unsigned(reg149) : reg139) ?
                  ($signed((~^reg120)) <= $signed($signed(reg132))) : $signed((^reg120[(2'h2):(1'h0)]))));
              reg150 <= ($unsigned(({reg139[(1'h0):(1'h0)],
                  (reg118 | reg149)} | reg127[(4'hb):(3'h4)])) + (((~&$signed((8'hb7))) ?
                  (~$signed(forvar111)) : reg130[(2'h3):(2'h3)]) != $unsigned(reg118)));
            end
        end
      else
        begin
          reg137 = ($signed(forvar111[(3'h4):(2'h2)]) ? reg129 : (8'hbb));
          reg138 <= (+(((-(reg114 ^ reg125)) ?
              ((reg144 ? forvar111 : reg120) ?
                  reg116[(4'ha):(4'h9)] : $signed(wire106)) : ((reg119 ^~ wire108) ?
                  {(7'h47), wire107} : reg116)) >= reg118[(4'hc):(3'h5)]));
          reg140 = reg127[(3'h7):(1'h0)];
          for (forvar141 = (1'h0); (forvar141 < (2'h2)); forvar141 = (forvar141 + (1'h1)))
            begin
              reg143 = ({(8'haf)} ^~ reg138);
            end
        end
      for (forvar151 = (1'h0); (forvar151 < (3'h4)); forvar151 = (forvar151 + (1'h1)))
        begin
          reg152 <= reg149[(3'h4):(2'h3)];
          reg153 = reg133[(3'h6):(2'h2)];
          reg154 <= reg138;
          for (forvar155 = (1'h0); (forvar155 < (2'h3)); forvar155 = (forvar155 + (1'h1)))
            begin
              reg156 = reg145[(3'h5):(2'h2)];
              reg157 <= ((((7'h49) + reg127[(3'h4):(2'h2)]) < $signed(reg146)) ?
                  reg135 : $unsigned((-((reg118 == reg139) && (~|reg121)))));
            end
          if ((~(reg148 ? (~|$unsigned({reg116, reg123})) : wire108)))
            begin
              reg158 = (~$unsigned((reg121[(1'h1):(1'h1)] <= ({reg149} >= (&reg149)))));
              reg159 <= ((8'hbe) != (8'ha6));
              reg160 = $signed(reg137);
            end
          else
            begin
              reg158 = reg153[(1'h0):(1'h0)];
              reg159 <= (({($signed(forvar151) ?
                      forvar112 : (&reg136))} && (~reg157[(4'he):(4'h9)])) * ({$unsigned((reg134 ?
                      reg133 : reg152)),
                  $signed((reg127 >= reg145))} * reg114));
              reg160 = $unsigned(forvar138);
              reg161 = $signed(wire110[(1'h1):(1'h1)]);
              reg162 = reg115[(4'h8):(2'h3)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar163 = (1'h0); (forvar163 < (3'h4)); forvar163 = (forvar163 + (1'h1)))
        begin
          for (forvar164 = (1'h0); (forvar164 < (2'h2)); forvar164 = (forvar164 + (1'h1)))
            begin
              reg165 = $signed((~^reg145[(2'h2):(2'h2)]));
            end
          reg166 <= $signed((!wire109));
          for (forvar167 = (1'h0); (forvar167 < (1'h1)); forvar167 = (forvar167 + (1'h1)))
            begin
              reg168 <= (~&$unsigned((8'haf)));
              reg169 = $unsigned(reg150);
              reg170 = reg130;
            end
          for (forvar171 = (1'h0); (forvar171 < (1'h1)); forvar171 = (forvar171 + (1'h1)))
            begin
              reg172 <= (~|$unsigned($unsigned(reg168)));
            end
        end
      for (forvar173 = (1'h0); (forvar173 < (2'h3)); forvar173 = (forvar173 + (1'h1)))
        begin
          reg174 <= (|$signed(reg172[(3'h4):(2'h3)]));
          reg175 = (~^(|($signed($unsigned(reg166)) <= $unsigned((reg130 ?
              reg170 : reg123)))));
        end
    end
  always
    @(posedge clk) begin
      if (reg168[(3'h5):(1'h0)])
        begin
          reg176 <= ((reg157 < $unsigned($signed((-reg154)))) <= reg152[(4'h9):(1'h1)]);
          reg177 = ((&reg145) ?
              (^~reg135) : ((wire108[(1'h1):(1'h0)] && $signed((+reg166))) ?
                  (8'hb5) : {reg138[(1'h1):(1'h0)],
                      ((wire106 >> reg138) ?
                          (&reg174) : reg130[(1'h0):(1'h0)])}));
          for (forvar178 = (1'h0); (forvar178 < (2'h2)); forvar178 = (forvar178 + (1'h1)))
            begin
              reg179 <= ((~|($signed((-reg134)) ?
                  (^(reg168 - reg154)) : ($signed(reg174) ^~ reg172[(3'h4):(2'h2)]))) * reg135[(1'h0):(1'h0)]);
              reg180 <= forvar178;
              reg181 = ((!wire110) << ((|reg113) < reg123[(4'hb):(1'h0)]));
            end
          reg182 = (((~((!wire108) >>> (reg150 ?
                  wire109 : (8'hb8)))) <<< (reg159[(2'h3):(2'h3)] ?
                  $signed((reg141 ?
                      reg124 : reg150)) : reg114[(4'h8):(3'h7)])) ?
              ($signed(($unsigned((8'hb6)) >>> $unsigned((8'ha3)))) ?
                  ($signed(((8'hbd) ?
                      reg180 : wire106)) ^~ (~&reg134[(1'h1):(1'h0)])) : $signed((forvar178[(3'h5):(3'h5)] | reg134[(1'h1):(1'h1)]))) : $signed((!reg126)));
          for (forvar183 = (1'h0); (forvar183 < (1'h0)); forvar183 = (forvar183 + (1'h1)))
            begin
              reg184 <= ($signed((~(~reg126))) < reg145);
            end
        end
      else
        begin
          reg176 <= {(|(~&((!reg126) ?
                  (reg129 ? reg148 : (8'haa)) : {reg180, reg159})))};
        end
    end
  assign wire185 = reg126;
  always
    @(posedge clk) begin
      reg186 <= $unsigned($unsigned($signed(reg180)));
    end
  assign wire187 = ((reg186[(2'h3):(2'h2)] ?
                       (^~($signed(reg150) <<< (8'ha4))) : $unsigned($unsigned((reg114 > reg186)))) < reg150[(4'h9):(3'h7)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module200  (y, clk, wire201, wire202, wire203, wire204, wire205);
  output wire [(32'h927):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire201;
  input wire [(5'h15):(1'h0)] wire202;
  input wire [(5'h18):(1'h0)] wire203;
  input wire [(3'h6):(1'h0)] wire204;
  input wire signed [(2'h3):(1'h0)] wire205;
  wire [(4'hd):(1'h0)] wire1380;
  wire [(2'h3):(1'h0)] wire1243;
  wire [(4'he):(1'h0)] wire872;
  wire signed [(5'h14):(1'h0)] wire829;
  wire [(4'hb):(1'h0)] wire828;
  wire signed [(2'h3):(1'h0)] wire827;
  wire [(4'he):(1'h0)] wire786;
  wire signed [(5'h12):(1'h0)] wire206;
  wire [(5'h10):(1'h0)] wire254;
  wire signed [(4'ha):(1'h0)] wire616;
  wire signed [(4'hf):(1'h0)] wire1378;
  reg [(5'h18):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg898 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg897 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg894 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg891 = (1'h0);
  reg [(3'h4):(1'h0)] reg890 = (1'h0);
  reg [(4'hc):(1'h0)] reg885 = (1'h0);
  reg [(5'h10):(1'h0)] reg880 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg878 = (1'h0);
  reg [(2'h2):(1'h0)] reg876 = (1'h0);
  reg [(5'h13):(1'h0)] reg871 = (1'h0);
  reg [(4'hb):(1'h0)] reg864 = (1'h0);
  reg [(2'h2):(1'h0)] reg859 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg869 = (1'h0);
  reg [(4'hb):(1'h0)] reg867 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg866 = (1'h0);
  reg [(4'he):(1'h0)] reg863 = (1'h0);
  reg [(5'h10):(1'h0)] reg861 = (1'h0);
  reg [(2'h3):(1'h0)] reg855 = (1'h0);
  reg [(5'h16):(1'h0)] reg854 = (1'h0);
  reg [(5'h10):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg849 = (1'h0);
  reg [(3'h5):(1'h0)] reg843 = (1'h0);
  reg [(3'h5):(1'h0)] reg842 = (1'h0);
  reg [(5'h11):(1'h0)] reg841 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg838 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg836 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg834 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg825 = (1'h0);
  reg [(5'h13):(1'h0)] reg824 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg819 = (1'h0);
  reg [(4'hd):(1'h0)] reg816 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg823 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg818 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg814 = (1'h0);
  reg [(4'he):(1'h0)] reg812 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg797 = (1'h0);
  reg [(5'h12):(1'h0)] reg808 = (1'h0);
  reg [(5'h15):(1'h0)] reg807 = (1'h0);
  reg [(4'h8):(1'h0)] reg806 = (1'h0);
  reg [(3'h7):(1'h0)] reg804 = (1'h0);
  reg [(5'h17):(1'h0)] reg800 = (1'h0);
  reg [(2'h3):(1'h0)] reg795 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg793 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg790 = (1'h0);
  reg [(5'h17):(1'h0)] reg788 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg253 = (1'h0);
  reg [(5'h13):(1'h0)] reg252 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg246 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg245 = (1'h0);
  reg [(5'h18):(1'h0)] reg244 = (1'h0);
  reg [(4'h9):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg240 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg239 = (1'h0);
  reg [(5'h10):(1'h0)] reg238 = (1'h0);
  reg [(3'h6):(1'h0)] reg236 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg235 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg230 = (1'h0);
  reg [(4'he):(1'h0)] reg229 = (1'h0);
  reg [(3'h5):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg224 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg223 = (1'h0);
  reg [(5'h18):(1'h0)] reg213 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg210 = (1'h0);
  reg [(5'h16):(1'h0)] reg618 = (1'h0);
  reg [(4'hc):(1'h0)] reg899 = (1'h0);
  reg [(4'ha):(1'h0)] reg896 = (1'h0);
  reg [(5'h13):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar893 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg892 = (1'h0);
  reg [(4'he):(1'h0)] reg889 = (1'h0);
  reg [(3'h7):(1'h0)] reg888 = (1'h0);
  reg [(5'h15):(1'h0)] reg887 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg886 = (1'h0);
  reg [(2'h2):(1'h0)] reg884 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg883 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg882 = (1'h0);
  reg [(3'h5):(1'h0)] reg881 = (1'h0);
  reg [(5'h10):(1'h0)] reg879 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg877 = (1'h0);
  reg [(4'h8):(1'h0)] forvar875 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg874 = (1'h0);
  reg [(3'h5):(1'h0)] forvar873 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg868 = (1'h0);
  reg [(4'ha):(1'h0)] forvar860 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg870 = (1'h0);
  reg [(2'h3):(1'h0)] forvar868 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg865 = (1'h0);
  reg [(2'h3):(1'h0)] forvar864 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg862 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg860 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar859 = (1'h0);
  reg [(5'h18):(1'h0)] reg858 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg857 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg856 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg853 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg852 = (1'h0);
  reg [(3'h5):(1'h0)] reg850 = (1'h0);
  reg [(4'ha):(1'h0)] reg848 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg847 = (1'h0);
  reg [(5'h15):(1'h0)] reg846 = (1'h0);
  reg [(5'h14):(1'h0)] forvar845 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg844 = (1'h0);
  reg [(5'h16):(1'h0)] reg840 = (1'h0);
  reg [(4'h8):(1'h0)] forvar839 = (1'h0);
  reg [(5'h11):(1'h0)] forvar837 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg835 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg833 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg832 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar831 = (1'h0);
  reg [(3'h4):(1'h0)] forvar830 = (1'h0);
  reg [(5'h18):(1'h0)] reg826 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar813 = (1'h0);
  reg [(3'h4):(1'h0)] reg822 = (1'h0);
  reg [(4'he):(1'h0)] reg821 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg820 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar819 = (1'h0);
  reg [(4'h9):(1'h0)] reg817 = (1'h0);
  reg [(4'he):(1'h0)] forvar816 = (1'h0);
  reg [(4'hf):(1'h0)] reg815 = (1'h0);
  reg [(5'h17):(1'h0)] reg813 = (1'h0);
  reg [(4'hf):(1'h0)] reg811 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar810 = (1'h0);
  reg [(5'h10):(1'h0)] forvar809 = (1'h0);
  reg [(5'h17):(1'h0)] forvar802 = (1'h0);
  reg [(5'h11):(1'h0)] forvar798 = (1'h0);
  reg [(5'h14):(1'h0)] reg805 = (1'h0);
  reg [(4'h8):(1'h0)] reg803 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg802 = (1'h0);
  reg [(2'h2):(1'h0)] reg801 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg799 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg798 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar797 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg796 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar790 = (1'h0);
  reg [(4'he):(1'h0)] reg794 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg792 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg791 = (1'h0);
  reg [(3'h4):(1'h0)] reg789 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg251 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg250 = (1'h0);
  reg [(5'h18):(1'h0)] reg249 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg248 = (1'h0);
  reg [(4'hc):(1'h0)] reg247 = (1'h0);
  reg [(2'h2):(1'h0)] forvar239 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg243 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg242 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg237 = (1'h0);
  reg [(5'h18):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg233 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar232 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg231 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar228 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg226 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar222 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar221 = (1'h0);
  reg [(4'h9):(1'h0)] reg220 = (1'h0);
  reg [(4'h8):(1'h0)] reg219 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg218 = (1'h0);
  reg [(3'h5):(1'h0)] forvar217 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg216 = (1'h0);
  reg [(3'h6):(1'h0)] reg208 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg215 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg214 = (1'h0);
  reg [(3'h5):(1'h0)] forvar212 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg211 = (1'h0);
  reg [(4'hf):(1'h0)] reg209 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar208 = (1'h0);
  reg [(3'h7):(1'h0)] reg207 = (1'h0);
  assign y = {wire1380,
                 wire1243,
                 wire872,
                 wire829,
                 wire828,
                 wire827,
                 wire786,
                 wire206,
                 wire254,
                 wire616,
                 wire1378,
                 reg900,
                 reg898,
                 reg897,
                 reg894,
                 reg891,
                 reg890,
                 reg885,
                 reg880,
                 reg878,
                 reg876,
                 reg871,
                 reg864,
                 reg859,
                 reg869,
                 reg867,
                 reg866,
                 reg863,
                 reg861,
                 reg855,
                 reg854,
                 reg851,
                 reg849,
                 reg843,
                 reg842,
                 reg841,
                 reg838,
                 reg836,
                 reg834,
                 reg825,
                 reg824,
                 reg819,
                 reg816,
                 reg823,
                 reg818,
                 reg814,
                 reg812,
                 reg797,
                 reg808,
                 reg807,
                 reg806,
                 reg804,
                 reg800,
                 reg795,
                 reg793,
                 reg790,
                 reg788,
                 reg253,
                 reg252,
                 reg246,
                 reg245,
                 reg244,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg236,
                 reg235,
                 reg230,
                 reg229,
                 reg227,
                 reg225,
                 reg224,
                 reg223,
                 reg213,
                 reg210,
                 reg618,
                 reg899,
                 reg896,
                 reg895,
                 forvar893,
                 reg892,
                 reg889,
                 reg888,
                 reg887,
                 reg886,
                 reg884,
                 reg883,
                 reg882,
                 reg881,
                 reg879,
                 reg877,
                 forvar875,
                 reg874,
                 forvar873,
                 reg868,
                 forvar860,
                 reg870,
                 forvar868,
                 reg865,
                 forvar864,
                 reg862,
                 reg860,
                 forvar859,
                 reg858,
                 reg857,
                 reg856,
                 reg853,
                 reg852,
                 reg850,
                 reg848,
                 reg847,
                 reg846,
                 forvar845,
                 reg844,
                 reg840,
                 forvar839,
                 forvar837,
                 reg835,
                 reg833,
                 reg832,
                 forvar831,
                 forvar830,
                 reg826,
                 forvar813,
                 reg822,
                 reg821,
                 reg820,
                 forvar819,
                 reg817,
                 forvar816,
                 reg815,
                 reg813,
                 reg811,
                 forvar810,
                 forvar809,
                 forvar802,
                 forvar798,
                 reg805,
                 reg803,
                 reg802,
                 reg801,
                 reg799,
                 reg798,
                 forvar797,
                 reg796,
                 forvar790,
                 reg794,
                 reg792,
                 reg791,
                 reg789,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 forvar239,
                 reg243,
                 reg242,
                 reg237,
                 reg234,
                 reg233,
                 forvar232,
                 reg231,
                 forvar228,
                 reg226,
                 forvar222,
                 forvar221,
                 reg220,
                 reg219,
                 reg218,
                 forvar217,
                 reg216,
                 reg208,
                 reg215,
                 reg214,
                 forvar212,
                 reg211,
                 reg209,
                 forvar208,
                 reg207,
                 (1'h0)};
  assign wire206 = wire203[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg207 = ((8'hae) && ($unsigned({{wire204}}) ?
          $signed($unsigned((~(8'hb6)))) : $signed(wire205)));
      if (reg207[(2'h3):(1'h0)])
        begin
          for (forvar208 = (1'h0); (forvar208 < (2'h2)); forvar208 = (forvar208 + (1'h1)))
            begin
              reg209 = wire203[(2'h2):(1'h1)];
              reg210 <= {{$unsigned(($unsigned(wire202) <<< $signed(wire201)))},
                  $signed({(~&wire206[(4'ha):(3'h5)])})};
            end
          reg211 = $signed({(8'ha3)});
          for (forvar212 = (1'h0); (forvar212 < (3'h4)); forvar212 = (forvar212 + (1'h1)))
            begin
              reg213 <= $signed($signed((^(&reg210[(4'h8):(3'h6)]))));
              reg214 = (wire205[(2'h3):(2'h2)] ?
                  (^$signed({(reg211 ? wire201 : reg209),
                      reg207[(3'h5):(3'h4)]})) : $unsigned($unsigned((~&$unsigned(reg207)))));
              reg215 = $signed((~&$signed({$unsigned(forvar208),
                  $signed((7'h48))})));
            end
        end
      else
        begin
          reg208 = (&(&$unsigned(wire206)));
        end
      reg216 = ((~(($unsigned(wire205) < (~&wire203)) + reg213[(5'h14):(4'hc)])) ?
          $unsigned(reg214[(2'h3):(1'h0)]) : $signed((8'h9e)));
      for (forvar217 = (1'h0); (forvar217 < (1'h1)); forvar217 = (forvar217 + (1'h1)))
        begin
          reg218 = {$signed((~^reg211[(4'he):(4'h9)])),
              ((^~reg214[(3'h7):(3'h5)]) ?
                  ((~^{wire202}) == ((8'hab) ?
                      {(8'ha0)} : (&reg211))) : (($signed(wire202) ^ (wire201 ?
                          reg214 : wire201)) ?
                      (~^(reg209 ? (7'h4a) : reg209)) : ((8'ha4) ?
                          $signed(reg213) : {wire202, reg209})))};
        end
    end
  always
    @(posedge clk) begin
      if ((^($unsigned(wire204[(3'h6):(2'h2)]) >> ((wire203[(1'h1):(1'h1)] && (reg213 ?
          wire204 : wire202)) >= $signed($signed(wire206))))))
        begin
          reg219 = $unsigned((($unsigned((~^wire202)) == wire202) ?
              $unsigned(((reg213 * reg213) ?
                  wire202[(2'h2):(1'h1)] : (^reg210))) : reg210[(1'h0):(1'h0)]));
        end
      else
        begin
          reg219 = wire205[(1'h0):(1'h0)];
        end
      reg220 = wire203[(2'h3):(2'h3)];
      for (forvar221 = (1'h0); (forvar221 < (1'h1)); forvar221 = (forvar221 + (1'h1)))
        begin
          for (forvar222 = (1'h0); (forvar222 < (1'h0)); forvar222 = (forvar222 + (1'h1)))
            begin
              reg223 <= wire201[(2'h2):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg224 <= (wire203 ?
          (!(!((-(8'ha3)) ?
              reg210 : (wire204 ?
                  wire202 : wire201)))) : $unsigned((~&(wire202[(4'h9):(4'h8)] ?
              $unsigned(reg213) : (wire204 << wire204)))));
      reg225 <= reg210;
      reg226 = $signed((&reg223[(2'h3):(1'h0)]));
      reg227 <= wire204;
    end
  always
    @(posedge clk) begin
      for (forvar228 = (1'h0); (forvar228 < (1'h1)); forvar228 = (forvar228 + (1'h1)))
        begin
          reg229 <= reg223;
          reg230 <= $unsigned((reg213[(4'hb):(3'h4)] ?
              (({reg229} || {reg213}) + {(-reg227)}) : (-wire205[(2'h2):(1'h0)])));
          reg231 = ((8'hbd) ?
              ($signed((7'h41)) + reg227[(2'h2):(2'h2)]) : {$signed((-((7'h44) ?
                      reg227 : wire204)))});
          for (forvar232 = (1'h0); (forvar232 < (2'h3)); forvar232 = (forvar232 + (1'h1)))
            begin
              reg233 = reg230;
              reg234 = reg224;
              reg235 <= reg223;
              reg236 <= (reg210 ?
                  $unsigned($unsigned(reg223)) : $signed(wire203[(1'h0):(1'h0)]));
            end
        end
      reg237 = ($signed($signed(reg231[(3'h5):(2'h3)])) ^~ wire202[(5'h15):(2'h3)]);
      if (reg235)
        begin
          reg238 <= ((^~(^~wire204[(3'h4):(2'h2)])) > (~&({$unsigned((8'hb5)),
                  $signed(reg229)} ?
              ({wire203,
                  (8'ha6)} - $unsigned(reg227)) : (reg236[(2'h3):(1'h1)] < (reg229 || reg230)))));
          reg239 <= (((forvar232 ?
                  $unsigned(reg223[(2'h2):(1'h1)]) : {(reg234 != reg237),
                      ((7'h49) == reg234)}) * $unsigned(reg210[(1'h0):(1'h0)])) ?
              $unsigned(reg231) : reg210[(2'h3):(2'h3)]);
          if ($unsigned(reg231[(2'h2):(2'h2)]))
            begin
              reg240 <= $signed({reg229[(4'ha):(1'h0)],
                  {reg237[(1'h0):(1'h0)], (-(|wire203))}});
              reg241 <= (~|((7'h40) ?
                  {$signed(reg213)} : {$signed(reg229[(4'hb):(4'ha)]),
                      $unsigned({wire203, reg233})}));
            end
          else
            begin
              reg240 <= {(wire205[(1'h0):(1'h0)] * $unsigned((-(~&reg235))))};
              reg242 = ($signed(forvar232[(1'h1):(1'h1)]) >>> $signed({(!$unsigned(wire205)),
                  (|$unsigned(reg234))}));
              reg243 = $unsigned(reg242);
              reg244 <= ((reg210 != reg229[(4'he):(4'h9)]) || reg224);
            end
        end
      else
        begin
          reg238 <= {((((7'h47) <<< (forvar228 >> (8'ha2))) ?
                      forvar232[(1'h1):(1'h0)] : $unsigned(reg238[(3'h6):(1'h1)])) ?
                  (^~reg231) : ({$unsigned((8'hb5)), (-reg225)} - ((reg240 ?
                          reg238 : reg230) ?
                      {wire202, reg244} : (reg244 ~^ reg241)))),
              reg224[(4'hd):(3'h6)]};
          for (forvar239 = (1'h0); (forvar239 < (1'h1)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg240 <= wire201[(4'h9):(1'h0)];
              reg242 = $unsigned($unsigned(wire201[(4'ha):(2'h3)]));
              reg243 = {(reg210[(4'h8):(2'h3)] || $signed((!{reg237, reg235}))),
                  ($signed($unsigned((!reg239))) ?
                      $unsigned({$unsigned(reg231),
                          (|reg244)}) : (($signed(wire203) - reg223[(3'h7):(3'h7)]) - {$signed(wire202),
                          (reg213 == (8'hae))}))};
              reg244 <= reg236;
            end
          if ($signed($unsigned(reg224)))
            begin
              reg245 <= $unsigned({wire205});
              reg246 <= $signed(reg227);
            end
          else
            begin
              reg245 <= (reg213 >= (forvar228[(2'h3):(1'h0)] << ((~|(!forvar239)) ?
                  (~|(reg244 ? (8'hae) : wire202)) : reg227)));
              reg246 <= (wire206[(2'h2):(1'h0)] ?
                  (^~(~((+reg245) ?
                      (reg210 ?
                          reg229 : forvar232) : reg245[(4'ha):(2'h2)]))) : (reg241[(3'h7):(3'h7)] << reg229[(2'h2):(2'h2)]));
            end
          if ({($signed(((^wire203) * $signed(reg237))) | ((reg223 == {(8'haf)}) > $signed({reg243})))})
            begin
              reg247 = reg230;
              reg248 = $unsigned(((((reg229 >> wire202) ?
                          $signed(wire203) : (~|reg236)) ?
                      (reg224[(1'h0):(1'h0)] ?
                          $unsigned(reg245) : $signed(reg247)) : (&(reg240 ^~ forvar232))) ?
                  (reg223[(1'h0):(1'h0)] - ($unsigned(reg224) >= (^wire205))) : (+reg241)));
              reg249 = {reg245, $unsigned(reg236)};
              reg250 = {(7'h41),
                  (reg213[(3'h6):(1'h0)] ?
                      wire205 : ((reg236 > reg235[(2'h3):(1'h0)]) + (+((8'ha3) ?
                          forvar239 : (8'hbe)))))};
              reg251 = $signed($unsigned((reg248 ~^ (~$unsigned((7'h45))))));
            end
          else
            begin
              reg247 = $signed((!({$unsigned((8'ha0)),
                  $signed(reg246)} <= ((reg236 ?
                  reg213 : reg242) ~^ reg242[(3'h4):(2'h3)]))));
              reg248 = reg247[(3'h5):(3'h5)];
              reg249 = $unsigned({{$signed((reg237 ? wire205 : reg231))}});
              reg250 = $unsigned((7'h48));
            end
          reg252 <= ($signed($unsigned($unsigned($signed(reg236)))) ?
              (((reg241[(3'h7):(3'h6)] ?
                      reg236[(2'h3):(1'h1)] : $signed(reg210)) != $signed(((8'hb2) ?
                      reg235 : reg230))) ?
                  (&reg231) : reg240[(1'h0):(1'h0)]) : wire203);
        end
      reg253 <= $signed(reg227[(2'h2):(1'h0)]);
    end
  assign wire254 = $unsigned($unsigned((~|(^reg223))));
  module255 #() modinst617 (wire616, clk, wire203, reg225, reg238, reg223);
  always
    @(posedge clk) begin
      reg618 <= {reg235,
          (({reg213[(4'ha):(3'h7)]} ? $signed($signed(wire616)) : reg223) ?
              (~&(-(reg210 ? reg230 : reg210))) : (wire206 ?
                  {(wire206 < reg236), reg244[(3'h4):(2'h2)]} : reg213))};
    end
  module619 #() modinst787 (wire786, clk, reg224, reg227, wire203, wire206, reg252);
  always
    @(posedge clk) begin
      if ((reg239[(3'h7):(3'h6)] && (($unsigned(((8'h9d) ? reg241 : reg223)) ?
          reg236[(3'h6):(1'h1)] : reg239) + $signed({reg252,
          ((7'h46) && wire201)}))))
        begin
          reg788 <= (&{(~^((reg227 ? (8'ha3) : reg236) ?
                  wire205[(2'h2):(2'h2)] : {reg236})),
              (|wire202)});
          if (reg210)
            begin
              reg789 = $signed((reg229 ?
                  (~^$unsigned($unsigned(wire201))) : {(|{reg213})}));
              reg790 <= (^wire254[(2'h2):(1'h1)]);
              reg791 = ({(8'hb0), $signed(reg618)} ?
                  (8'hb3) : (~$unsigned(wire203[(4'hb):(3'h7)])));
            end
          else
            begin
              reg790 <= wire206[(3'h7):(2'h3)];
              reg791 = {(!reg229[(2'h2):(1'h1)])};
              reg792 = (^~wire202[(3'h4):(2'h2)]);
              reg793 <= (~&$signed($signed(wire786)));
              reg794 = (-wire203);
            end
          reg795 <= reg230;
        end
      else
        begin
          reg788 <= $signed((~^(reg793[(4'h9):(3'h4)] < $unsigned($unsigned(wire616)))));
          reg789 = {$unsigned((~reg240[(4'hc):(2'h3)]))};
          for (forvar790 = (1'h0); (forvar790 < (1'h0)); forvar790 = (forvar790 + (1'h1)))
            begin
              reg791 = wire204[(1'h1):(1'h0)];
              reg793 <= (forvar790 ? wire201[(3'h6):(2'h2)] : (7'h45));
              reg794 = (((|((~reg245) ? reg788 : (!wire254))) == (((~^reg227) ?
                          $signed(wire786) : {reg788}) ?
                      (|reg618) : (^{reg253}))) ?
                  reg245 : (reg788[(4'hb):(4'h8)] ?
                      reg790[(5'h11):(4'hb)] : ((~|reg225) ^ ($unsigned(forvar790) ^~ $signed(reg252)))));
              reg796 = wire203;
            end
        end
      if (((~|reg252) ?
          (($signed((~^reg253)) ^ (~^(|reg618))) <<< reg213[(5'h12):(4'hb)]) : {$unsigned(((reg792 || reg246) && $unsigned((7'h45)))),
              (-reg795[(2'h2):(2'h2)])}))
        begin
          for (forvar797 = (1'h0); (forvar797 < (3'h4)); forvar797 = (forvar797 + (1'h1)))
            begin
              reg798 = reg253;
              reg799 = {({reg227[(1'h0):(1'h0)]} < ($unsigned($signed(reg238)) ?
                      (~(reg229 ? reg210 : (8'hb5))) : ((~&wire204) ?
                          reg230[(3'h6):(2'h3)] : reg239))),
                  reg796};
              reg800 <= $signed(reg241);
            end
          reg801 = wire786;
          if (reg235[(2'h3):(1'h1)])
            begin
              reg802 = reg229;
              reg803 = (&($unsigned(reg225) <= (8'ha2)));
              reg804 <= ($unsigned(reg245[(1'h0):(1'h0)]) - (reg802[(4'he):(4'h8)] ?
                  reg800[(3'h6):(3'h5)] : reg238));
              reg805 = reg213[(5'h11):(4'hd)];
              reg806 <= $unsigned($signed(wire201));
            end
          else
            begin
              reg804 <= (8'ha1);
              reg805 = (({(reg789[(3'h4):(1'h0)] ?
                          $signed(reg246) : {(7'h45), reg799})} ?
                  reg236 : (reg794 + (reg252[(4'hd):(4'h9)] <<< {reg798}))) > (~|(8'hac)));
              reg806 <= reg806[(3'h6):(1'h1)];
              reg807 <= reg245[(1'h1):(1'h0)];
              reg808 <= (~&forvar797[(4'h8):(3'h7)]);
            end
        end
      else
        begin
          reg797 <= ((&reg804[(3'h4):(1'h0)]) <= reg245[(4'hb):(3'h5)]);
          for (forvar798 = (1'h0); (forvar798 < (3'h4)); forvar798 = (forvar798 + (1'h1)))
            begin
              reg799 = reg800[(5'h12):(4'hf)];
              reg800 <= (reg802[(4'he):(4'h9)] && (^~wire786));
              reg801 = reg235;
            end
          for (forvar802 = (1'h0); (forvar802 < (1'h1)); forvar802 = (forvar802 + (1'h1)))
            begin
              reg804 <= reg210[(2'h3):(2'h2)];
              reg805 = ($unsigned((-$unsigned((reg239 >> (8'haa))))) ?
                  (^~$unsigned(($unsigned(wire254) ?
                      $signed(reg788) : {forvar797}))) : forvar797);
              reg806 <= $unsigned((reg790 ?
                  $unsigned(((|reg252) != (wire616 >>> reg807))) : (((~&wire202) ^ reg227[(2'h2):(1'h0)]) >>> (forvar790[(4'hf):(3'h7)] ?
                      reg791 : $signed(wire204)))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar809 = (1'h0); (forvar809 < (1'h1)); forvar809 = (forvar809 + (1'h1)))
        begin
          for (forvar810 = (1'h0); (forvar810 < (3'h4)); forvar810 = (forvar810 + (1'h1)))
            begin
              reg811 = reg227[(1'h1):(1'h1)];
            end
          reg812 <= $unsigned((^forvar810[(3'h5):(3'h5)]));
        end
      if ({($signed($unsigned($signed((8'hb9)))) | (^~wire206[(2'h3):(2'h3)])),
          ($unsigned(reg808) <<< reg241)})
        begin
          if ((^~($signed($signed((|(8'hbe)))) ?
              (8'ha7) : (((reg808 ? reg230 : wire201) == {reg225,
                  reg223}) ~^ {(^reg244)}))))
            begin
              reg813 = ($unsigned(((forvar810[(3'h6):(3'h4)] ?
                          (forvar810 ?
                              wire616 : reg797) : reg246[(3'h5):(3'h4)]) ?
                      ($signed((7'h45)) == wire203[(4'hd):(3'h7)]) : $unsigned($signed(reg241)))) ?
                  reg240[(1'h0):(1'h0)] : $unsigned((+{(reg229 < reg811)})));
              reg814 <= $unsigned(((!reg225) && {(^{reg224}),
                  ((reg235 ? reg245 : reg223) <<< (^~reg788))}));
            end
          else
            begin
              reg813 = reg800[(5'h10):(3'h4)];
              reg814 <= (&$unsigned((~(~&reg236[(1'h1):(1'h0)]))));
              reg815 = (|reg795);
            end
          for (forvar816 = (1'h0); (forvar816 < (2'h2)); forvar816 = (forvar816 + (1'h1)))
            begin
              reg817 = ({reg814[(2'h3):(2'h2)]} ^ (((~(+wire205)) ?
                  $signed($unsigned(wire786)) : reg807) * (^(!(wire202 && forvar810)))));
              reg818 <= ((reg806 & reg813) ?
                  $unsigned({reg213}) : ($unsigned((+$signed(forvar810))) <= (((reg213 | reg225) ?
                      $signed((8'haf)) : reg253[(3'h5):(3'h4)]) >= {wire204[(2'h2):(1'h1)]})));
            end
          for (forvar819 = (1'h0); (forvar819 < (1'h1)); forvar819 = (forvar819 + (1'h1)))
            begin
              reg820 = reg808;
              reg821 = reg807[(4'h9):(2'h2)];
              reg822 = ($unsigned(wire206) ^ {(reg815[(3'h7):(3'h4)] ?
                      reg804[(2'h2):(2'h2)] : {((8'ha2) >> wire206)})});
            end
          reg823 <= wire203[(3'h4):(1'h0)];
        end
      else
        begin
          for (forvar813 = (1'h0); (forvar813 < (1'h0)); forvar813 = (forvar813 + (1'h1)))
            begin
              reg815 = (($signed(reg227) ?
                      $unsigned($unsigned($signed(reg236))) : {(((8'ha0) ?
                                  reg797 : reg229) ?
                              {(8'hb0), wire205} : (^~reg811)),
                          ((8'hb0) ^ (reg795 ? wire205 : reg618))}) ?
                  $unsigned($signed($unsigned((reg244 >= wire203)))) : reg821[(4'ha):(3'h4)]);
              reg816 <= (8'hbf);
              reg818 <= (+(($signed((~^reg808)) * (reg223[(1'h1):(1'h0)] ?
                  (8'hb4) : (|reg800))) >>> ($signed($unsigned(reg811)) ^~ $signed((^reg823)))));
              reg819 <= reg618[(4'hf):(1'h1)];
              reg823 <= $signed((~&(^~({reg229, (8'hb4)} ?
                  (+reg818) : reg807[(5'h11):(5'h10)]))));
            end
        end
      reg824 <= $signed(reg245[(4'hb):(2'h2)]);
      reg825 <= {$signed(reg811),
          (~|$unsigned((reg820 + (reg213 ? reg807 : reg240))))};
      reg826 = ((+$unsigned(wire786[(4'he):(4'hc)])) ? reg808 : wire201);
    end
  assign wire827 = $unsigned((^~(((reg253 & reg227) ^ reg823) ?
                       wire203 : ((~|reg229) & (wire205 | (8'hb6))))));
  assign wire828 = $unsigned($signed($unsigned($signed(reg804[(3'h7):(2'h2)]))));
  assign wire829 = $unsigned((7'h49));
  always
    @(posedge clk) begin
      for (forvar830 = (1'h0); (forvar830 < (2'h3)); forvar830 = (forvar830 + (1'h1)))
        begin
          for (forvar831 = (1'h0); (forvar831 < (2'h2)); forvar831 = (forvar831 + (1'h1)))
            begin
              reg832 = ((reg800 ?
                  reg825[(2'h2):(2'h2)] : $unsigned($unsigned($signed(reg823)))) - wire254[(3'h7):(1'h1)]);
              reg833 = $unsigned(($unsigned((~&(reg808 == reg818))) >= (~(reg825[(1'h0):(1'h0)] ?
                  reg241 : wire206[(4'hb):(1'h0)]))));
              reg834 <= reg229[(2'h3):(1'h1)];
              reg835 = (reg795[(1'h0):(1'h0)] ?
                  ($signed($unsigned({reg807})) ?
                      reg812 : (+reg824[(4'h9):(2'h3)])) : (reg812[(4'hb):(2'h2)] | reg252[(3'h6):(2'h2)]));
              reg836 <= (+$signed((|{(reg834 ? forvar830 : reg797),
                  (~^wire786)})));
            end
        end
      for (forvar837 = (1'h0); (forvar837 < (1'h1)); forvar837 = (forvar837 + (1'h1)))
        begin
          reg838 <= $signed(reg816);
          for (forvar839 = (1'h0); (forvar839 < (2'h3)); forvar839 = (forvar839 + (1'h1)))
            begin
              reg840 = forvar837[(4'h9):(1'h0)];
              reg841 <= reg823;
              reg842 <= (~^$signed((^~((~reg239) <<< $signed(reg800)))));
            end
          reg843 <= $unsigned(reg235[(3'h5):(3'h5)]);
          reg844 = (((($unsigned(reg824) ?
                  (wire254 != (8'ha5)) : reg836[(2'h3):(2'h3)]) <<< (^wire202[(4'hc):(4'ha)])) ^~ $unsigned(((reg788 ?
                      reg618 : reg227) ?
                  $unsigned(wire254) : reg246[(3'h5):(1'h0)]))) ?
              {$unsigned(reg241[(3'h4):(1'h1)]),
                  (((reg824 ? reg814 : wire201) ?
                          $unsigned(reg840) : $unsigned(forvar837)) ?
                      ($signed(reg223) & ((8'ha0) == reg236)) : ((^~reg833) || wire616))} : (~^$unsigned({(!(8'hb0)),
                  (reg230 ? wire201 : reg618)})));
        end
      for (forvar845 = (1'h0); (forvar845 < (3'h4)); forvar845 = (forvar845 + (1'h1)))
        begin
          reg846 = (wire828 > reg814);
          if ((($signed($unsigned({(8'hbb),
                  wire201})) < $unsigned(reg804[(2'h3):(2'h2)])) ?
              (wire202 ?
                  ((reg253 ?
                      $unsigned(reg819) : reg227[(1'h0):(1'h0)]) && ($unsigned(reg806) ?
                      reg797[(1'h0):(1'h0)] : $signed(forvar837))) : ($signed(wire616) ?
                      $unsigned((reg788 ~^ forvar837)) : (8'had))) : reg808[(4'hb):(2'h2)]))
            begin
              reg847 = ($unsigned($unsigned(({reg213} ?
                      {reg793} : $unsigned(reg833)))) ?
                  reg824 : $signed($unsigned((~^$signed(reg790)))));
              reg848 = (reg840 ?
                  (({wire206[(4'h9):(3'h6)]} ?
                      reg252[(2'h3):(2'h3)] : reg843[(2'h2):(2'h2)]) * (~&reg227)) : reg841[(4'hc):(1'h1)]);
              reg849 <= (forvar831[(2'h3):(2'h3)] ?
                  reg804 : $unsigned($signed($signed($unsigned((8'hbb))))));
            end
          else
            begin
              reg847 = (($signed($unsigned(reg244[(5'h10):(4'hc)])) == (reg818 | reg224)) ?
                  {($unsigned(reg235[(4'h8):(3'h7)]) ?
                          $signed((reg240 >> (8'ha1))) : $unsigned(reg252[(4'h9):(2'h3)]))} : (reg239 ?
                      (~^reg808) : $signed($unsigned(reg253))));
              reg848 = ($signed(reg835) ? forvar837[(3'h4):(1'h0)] : reg844);
              reg850 = reg238[(2'h2):(1'h1)];
            end
          if ($unsigned(reg833[(2'h2):(1'h1)]))
            begin
              reg851 <= (wire616[(4'h9):(4'h8)] | (8'ha3));
              reg852 = $unsigned(reg235[(1'h1):(1'h0)]);
              reg853 = {(!$unsigned((+$unsigned(wire616)))),
                  reg844[(1'h1):(1'h0)]};
              reg854 <= ((((!(~|reg846)) ^ $signed((reg843 ?
                      reg239 : reg618))) ?
                  {reg235[(4'ha):(2'h2)]} : {((reg229 ?
                          reg851 : wire786) ^~ $unsigned((8'hb1)))}) && reg835);
              reg855 <= ({(~^wire206),
                      ((-(~|reg818)) ?
                          $unsigned($signed(wire829)) : (+(reg841 <= forvar831)))} ?
                  $signed(reg844) : ($signed(($signed((8'haa)) != (wire206 <= forvar839))) ?
                      {$signed($unsigned(wire828))} : (8'ha1)));
            end
          else
            begin
              reg851 <= {(reg838[(1'h1):(1'h0)] ?
                      ($unsigned((reg245 ? reg241 : reg847)) ?
                          ($signed(wire202) << reg824) : (8'hb1)) : $unsigned((~^$unsigned((8'haf)))))};
              reg854 <= reg816[(4'hc):(1'h1)];
            end
          reg856 = {reg236[(3'h4):(2'h3)]};
        end
      if ($unsigned({reg851}))
        begin
          reg857 = (^~(^reg846[(4'hc):(2'h3)]));
          reg858 = $signed(reg855[(2'h3):(1'h1)]);
          for (forvar859 = (1'h0); (forvar859 < (2'h2)); forvar859 = (forvar859 + (1'h1)))
            begin
              reg860 = ($unsigned($signed(($unsigned(forvar831) != {wire204}))) < ($signed(((wire206 ?
                      (8'had) : (8'h9d)) && $unsigned(reg848))) ?
                  {$signed($unsigned(wire828))} : reg800));
              reg861 <= (8'hab);
              reg862 = ($signed(reg847[(3'h7):(2'h2)]) >> reg836[(2'h2):(2'h2)]);
              reg863 <= $unsigned(($signed(reg833) ?
                  (8'h9e) : reg253[(1'h1):(1'h0)]));
            end
          for (forvar864 = (1'h0); (forvar864 < (2'h2)); forvar864 = (forvar864 + (1'h1)))
            begin
              reg865 = (wire206 ? wire202 : $signed(forvar845));
              reg866 <= reg797[(3'h5):(2'h3)];
              reg867 <= reg853;
            end
          for (forvar868 = (1'h0); (forvar868 < (2'h3)); forvar868 = (forvar868 + (1'h1)))
            begin
              reg869 <= $unsigned($signed((~^$signed({reg239, reg797}))));
              reg870 = $signed($signed((~|(~|$signed(reg240)))));
            end
        end
      else
        begin
          reg859 <= (reg843[(1'h1):(1'h0)] <= (~reg807[(4'hb):(1'h1)]));
          for (forvar860 = (1'h0); (forvar860 < (1'h0)); forvar860 = (forvar860 + (1'h1)))
            begin
              reg862 = ((reg841 ?
                  reg850 : ((^~$signed(reg854)) ?
                      reg814[(2'h3):(2'h3)] : $signed((forvar837 ?
                          reg245 : reg788)))) <= reg834[(4'hb):(4'hb)]);
              reg863 <= {(reg618[(2'h2):(1'h1)] ?
                      reg825 : {$unsigned((8'hbc)), reg860})};
              reg864 <= (({reg843[(3'h5):(1'h1)]} || ({(reg842 ?
                          (7'h48) : reg225)} <= (^~(reg238 - reg861)))) ?
                  $unsigned((((-reg819) >= (reg224 ?
                      forvar864 : reg870)) <<< ($signed(wire204) ?
                      (reg245 ?
                          wire828 : reg818) : (^reg816)))) : (~^(((reg240 <<< reg849) ?
                          (~&reg865) : (wire205 ? reg855 : reg224)) ?
                      $unsigned((reg854 ? reg229 : reg797)) : reg825)));
              reg866 <= reg863;
              reg868 = reg847;
            end
          reg869 <= (^~reg870[(2'h2):(1'h1)]);
        end
      reg871 <= reg853;
    end
  assign wire872 = reg252[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar873 = (1'h0); (forvar873 < (2'h3)); forvar873 = (forvar873 + (1'h1)))
        begin
          reg874 = (reg808[(3'h5):(1'h1)] >>> reg861);
          for (forvar875 = (1'h0); (forvar875 < (2'h3)); forvar875 = (forvar875 + (1'h1)))
            begin
              reg876 <= $unsigned($signed($signed((&((8'hb3) << reg210)))));
            end
          if ((^forvar873))
            begin
              reg877 = $signed((8'ha8));
              reg878 <= reg800;
              reg879 = wire616;
            end
          else
            begin
              reg878 <= $signed((wire872 >>> (|(!$unsigned((8'hb3))))));
              reg880 <= $signed((&(reg210[(3'h5):(3'h5)] ?
                  reg824[(4'hd):(3'h6)] : ($signed(reg851) ?
                      (reg227 ? wire872 : wire204) : (wire872 + (8'had))))));
              reg881 = $signed(reg223[(3'h5):(2'h3)]);
              reg882 = (~$signed((~^$signed(wire203))));
            end
          if (((reg236 ?
                  (~|(|reg239)) : (({reg804} ? {reg869} : $signed(reg867)) ?
                      reg797[(3'h4):(1'h0)] : (~&$unsigned(wire872)))) ?
              $signed(reg240) : ($unsigned($unsigned((wire616 ?
                  reg230 : (7'h48)))) + reg224)))
            begin
              reg883 = $signed((forvar873 == (+(&$unsigned(reg239)))));
              reg884 = ($unsigned($signed(reg880[(2'h2):(1'h0)])) >= $signed((($signed(reg878) >>> reg883[(4'he):(1'h1)]) | ((|reg824) ^~ $unsigned(reg241)))));
              reg885 <= (~|reg818);
            end
          else
            begin
              reg885 <= ($signed((reg823[(3'h4):(2'h3)] >>> $signed($signed(reg618)))) ?
                  reg866[(3'h7):(3'h5)] : (reg807[(3'h5):(2'h3)] ?
                      (reg235 ?
                          wire203 : ((^reg618) != $signed(wire829))) : reg245));
            end
          if ((((((reg797 ? reg823 : (8'haa)) > reg843[(1'h0):(1'h0)]) ?
                      wire786[(4'hb):(1'h0)] : (~|$signed(reg808))) ?
                  ($unsigned($signed(reg841)) ?
                      (!reg230[(1'h1):(1'h0)]) : reg824) : reg854) ?
              ($signed(reg618[(4'hf):(3'h4)]) ?
                  reg807 : reg863[(4'he):(4'he)]) : ((~{((8'ha4) << reg240),
                      (~|reg876)}) ?
                  wire206 : wire202)))
            begin
              reg886 = ({($signed($unsigned(reg244)) ?
                      $signed($unsigned(wire202)) : (~|(reg807 ?
                          reg253 : (8'hb9)))),
                  ($signed(((8'had) ?
                      wire254 : (8'hba))) - $signed($signed((8'h9e))))} >>> ($unsigned($signed(reg804[(3'h6):(3'h4)])) << $signed($unsigned(reg210))));
              reg887 = $unsigned((($signed($signed(reg236)) <<< $signed((reg253 ?
                  reg882 : reg788))) && (~|reg807[(5'h10):(3'h4)])));
              reg888 = reg882[(5'h10):(4'hf)];
              reg889 = ((((wire201[(4'h9):(3'h6)] ?
                  ((7'h4a) < reg825) : {reg834,
                      reg797}) + reg800[(1'h1):(1'h1)]) + reg235) != $signed($signed(reg880[(2'h2):(1'h1)])));
            end
          else
            begin
              reg890 <= {wire786};
            end
        end
      reg891 <= (!$signed(reg240[(1'h0):(1'h0)]));
      reg892 = $unsigned(($unsigned($unsigned(wire827)) ?
          $unsigned($signed($signed(reg230))) : $unsigned($unsigned((reg851 <= reg884)))));
      for (forvar893 = (1'h0); (forvar893 < (1'h0)); forvar893 = (forvar893 + (1'h1)))
        begin
          reg894 <= ($unsigned($signed(forvar873[(3'h4):(1'h1)])) ?
              reg863 : (reg867 ?
                  ((^~(^~reg224)) ?
                      reg793 : ((|reg223) ?
                          reg885[(2'h2):(2'h2)] : (reg886 >= reg241))) : (&reg825[(1'h0):(1'h0)])));
          reg895 = ((&wire205[(2'h3):(2'h3)]) >= $unsigned(reg797));
          reg896 = ((!$signed((-wire206))) ?
              $unsigned((|(reg808[(3'h6):(3'h5)] ?
                  (^wire201) : reg867[(2'h2):(2'h2)]))) : reg806);
          if ((reg238[(3'h4):(2'h2)] ^~ ({(~(wire204 ~^ reg818))} ^~ wire872[(2'h2):(1'h0)])))
            begin
              reg897 <= ((-(reg824[(4'hc):(3'h7)] >>> ((~^(8'h9c)) || $unsigned(reg246)))) ?
                  $unsigned(reg841) : {reg804[(2'h2):(1'h1)]});
              reg898 <= (-$unsigned($unsigned($unsigned((-reg213)))));
            end
          else
            begin
              reg899 = $unsigned($signed(reg816));
              reg900 <= {(reg887[(5'h15):(4'hf)] ~^ (reg227 ~^ ((reg239 ?
                      wire202 : reg223) * ((8'ha1) ? (7'h40) : reg880))))};
            end
        end
    end
  module901 #() modinst1244 (wire1243, clk, reg823, reg819, reg224, wire254, reg851);
  module1245 #() modinst1379 (.wire1250(reg891), .wire1249(reg235), .clk(clk), .wire1247(reg227), .y(wire1378), .wire1248(wire201), .wire1246(reg871));
  assign wire1380 = $signed($unsigned((~(^(~reg235)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1245
#(parameter param1376 = {(8'h9c), (((|((8'hbe) && (8'hab))) <<< (((8'hbc) ? (8'haf) : (8'hb4)) <<< ((8'hbd) ? (8'h9f) : (7'h40)))) & {(((7'h45) && (8'hbe)) ? (!(7'h45)) : {(8'hb5)}), (8'haa)})}, 
parameter param1377 = param1376)
(y, clk, wire1250, wire1249, wire1248, wire1247, wire1246);
  output wire [(32'h6d7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire1250;
  input wire signed [(4'hc):(1'h0)] wire1249;
  input wire signed [(4'hd):(1'h0)] wire1248;
  input wire signed [(3'h5):(1'h0)] wire1247;
  input wire [(5'h13):(1'h0)] wire1246;
  wire [(2'h2):(1'h0)] wire1349;
  wire signed [(2'h3):(1'h0)] wire1337;
  wire signed [(4'hb):(1'h0)] wire1336;
  wire signed [(5'h14):(1'h0)] wire1318;
  wire [(3'h5):(1'h0)] wire1317;
  wire [(2'h3):(1'h0)] wire1289;
  wire signed [(4'hf):(1'h0)] wire1284;
  wire [(5'h11):(1'h0)] wire1252;
  wire signed [(2'h2):(1'h0)] wire1251;
  reg signed [(5'h12):(1'h0)] reg1373 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1372 = (1'h0);
  reg [(5'h18):(1'h0)] reg1370 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1368 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1366 = (1'h0);
  reg [(2'h3):(1'h0)] reg1365 = (1'h0);
  reg [(5'h15):(1'h0)] reg1364 = (1'h0);
  reg [(5'h18):(1'h0)] reg1356 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1360 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1357 = (1'h0);
  reg [(3'h6):(1'h0)] reg1355 = (1'h0);
  reg [(4'h9):(1'h0)] reg1348 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1345 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1344 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1342 = (1'h0);
  reg [(3'h6):(1'h0)] reg1341 = (1'h0);
  reg [(4'h8):(1'h0)] reg1338 = (1'h0);
  reg [(4'hc):(1'h0)] reg1335 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1331 = (1'h0);
  reg [(5'h18):(1'h0)] reg1330 = (1'h0);
  reg [(2'h3):(1'h0)] reg1327 = (1'h0);
  reg [(4'ha):(1'h0)] reg1324 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1321 = (1'h0);
  reg [(4'h9):(1'h0)] reg1312 = (1'h0);
  reg [(2'h3):(1'h0)] reg1308 = (1'h0);
  reg [(5'h18):(1'h0)] reg1307 = (1'h0);
  reg [(5'h17):(1'h0)] reg1305 = (1'h0);
  reg [(5'h11):(1'h0)] reg1306 = (1'h0);
  reg [(5'h15):(1'h0)] reg1303 = (1'h0);
  reg [(4'h9):(1'h0)] reg1302 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1299 = (1'h0);
  reg [(4'hb):(1'h0)] reg1295 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1294 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1293 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1291 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1288 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1287 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1286 = (1'h0);
  reg [(2'h2):(1'h0)] reg1265 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1280 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1276 = (1'h0);
  reg [(3'h5):(1'h0)] reg1275 = (1'h0);
  reg [(4'h9):(1'h0)] reg1274 = (1'h0);
  reg [(4'hc):(1'h0)] reg1273 = (1'h0);
  reg [(4'h8):(1'h0)] reg1271 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1270 = (1'h0);
  reg [(5'h10):(1'h0)] reg1268 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1262 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1259 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1258 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1256 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1255 = (1'h0);
  reg [(4'hb):(1'h0)] reg1254 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1370 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1369 = (1'h0);
  reg [(4'ha):(1'h0)] reg1375 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1374 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1371 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1369 = (1'h0);
  reg [(3'h7):(1'h0)] reg1367 = (1'h0);
  reg [(4'ha):(1'h0)] reg1363 = (1'h0);
  reg [(5'h13):(1'h0)] reg1362 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1359 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1352 = (1'h0);
  reg [(5'h13):(1'h0)] reg1350 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1361 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1359 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1358 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1356 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1354 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1353 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1352 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1351 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1350 = (1'h0);
  reg [(4'hc):(1'h0)] reg1347 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1346 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1343 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1340 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1339 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1334 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1333 = (1'h0);
  reg [(5'h14):(1'h0)] reg1332 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1329 = (1'h0);
  reg [(2'h2):(1'h0)] reg1328 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1326 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1325 = (1'h0);
  reg [(3'h5):(1'h0)] reg1320 = (1'h0);
  reg [(4'hc):(1'h0)] reg1323 = (1'h0);
  reg [(4'h8):(1'h0)] reg1322 = (1'h0);
  reg [(4'he):(1'h0)] forvar1320 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1319 = (1'h0);
  reg [(4'he):(1'h0)] reg1316 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1315 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1314 = (1'h0);
  reg [(5'h11):(1'h0)] reg1313 = (1'h0);
  reg [(5'h18):(1'h0)] reg1311 = (1'h0);
  reg [(5'h11):(1'h0)] reg1310 = (1'h0);
  reg [(3'h5):(1'h0)] reg1309 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1306 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1300 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1298 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1305 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1304 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1301 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1300 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1298 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1297 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1296 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1292 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1290 = (1'h0);
  reg [(4'h9):(1'h0)] reg1285 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1283 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1282 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1281 = (1'h0);
  reg [(3'h7):(1'h0)] reg1279 = (1'h0);
  reg [(4'h8):(1'h0)] reg1278 = (1'h0);
  reg [(4'he):(1'h0)] forvar1277 = (1'h0);
  reg [(2'h3):(1'h0)] reg1272 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1269 = (1'h0);
  reg [(5'h14):(1'h0)] reg1267 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1266 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1265 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1264 = (1'h0);
  reg [(4'ha):(1'h0)] reg1263 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1261 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1260 = (1'h0);
  reg [(5'h13):(1'h0)] reg1257 = (1'h0);
  reg [(4'ha):(1'h0)] reg1253 = (1'h0);
  assign y = {wire1349,
                 wire1337,
                 wire1336,
                 wire1318,
                 wire1317,
                 wire1289,
                 wire1284,
                 wire1252,
                 wire1251,
                 reg1373,
                 reg1372,
                 reg1370,
                 reg1368,
                 reg1366,
                 reg1365,
                 reg1364,
                 reg1356,
                 reg1360,
                 reg1357,
                 reg1355,
                 reg1348,
                 reg1345,
                 reg1344,
                 reg1342,
                 reg1341,
                 reg1338,
                 reg1335,
                 reg1331,
                 reg1330,
                 reg1327,
                 reg1324,
                 reg1321,
                 reg1312,
                 reg1308,
                 reg1307,
                 reg1305,
                 reg1306,
                 reg1303,
                 reg1302,
                 reg1299,
                 reg1295,
                 reg1294,
                 reg1293,
                 reg1291,
                 reg1288,
                 reg1287,
                 reg1286,
                 reg1265,
                 reg1280,
                 reg1276,
                 reg1275,
                 reg1274,
                 reg1273,
                 reg1271,
                 reg1270,
                 reg1268,
                 reg1262,
                 reg1259,
                 reg1258,
                 reg1256,
                 reg1255,
                 reg1254,
                 forvar1370,
                 reg1369,
                 reg1375,
                 reg1374,
                 reg1371,
                 forvar1369,
                 reg1367,
                 reg1363,
                 reg1362,
                 forvar1359,
                 reg1352,
                 reg1350,
                 reg1361,
                 reg1359,
                 reg1358,
                 forvar1356,
                 reg1354,
                 reg1353,
                 forvar1352,
                 reg1351,
                 forvar1350,
                 reg1347,
                 reg1346,
                 reg1343,
                 reg1340,
                 reg1339,
                 reg1334,
                 forvar1333,
                 reg1332,
                 forvar1329,
                 reg1328,
                 reg1326,
                 reg1325,
                 reg1320,
                 reg1323,
                 reg1322,
                 forvar1320,
                 reg1319,
                 reg1316,
                 reg1315,
                 reg1314,
                 reg1313,
                 reg1311,
                 reg1310,
                 reg1309,
                 forvar1306,
                 reg1300,
                 forvar1298,
                 forvar1305,
                 reg1304,
                 reg1301,
                 forvar1300,
                 reg1298,
                 reg1297,
                 reg1296,
                 reg1292,
                 reg1290,
                 reg1285,
                 reg1283,
                 reg1282,
                 forvar1281,
                 reg1279,
                 reg1278,
                 forvar1277,
                 reg1272,
                 reg1269,
                 reg1267,
                 reg1266,
                 forvar1265,
                 reg1264,
                 reg1263,
                 reg1261,
                 reg1260,
                 reg1257,
                 reg1253,
                 (1'h0)};
  assign wire1251 = wire1248;
  assign wire1252 = wire1246;
  always
    @(posedge clk) begin
      if (wire1250)
        begin
          if ((~^({((wire1249 ^~ wire1248) ?
                      (|wire1247) : ((7'h46) || wire1251))} ?
              (((wire1250 ~^ (8'ha0)) <<< (wire1248 ?
                  wire1248 : wire1252)) && wire1249[(3'h5):(1'h0)]) : wire1248[(2'h3):(2'h2)])))
            begin
              reg1253 = (wire1249 + wire1247[(3'h5):(2'h3)]);
              reg1254 <= $unsigned(wire1251[(2'h2):(1'h1)]);
              reg1255 <= (({wire1249,
                      $signed((wire1246 ?
                          wire1249 : (8'hb8)))} | $unsigned(wire1250)) ?
                  wire1251 : {(((^~wire1249) >>> $signed(wire1249)) ?
                          reg1254 : (8'hbf)),
                      (^~$signed(reg1254))});
            end
          else
            begin
              reg1253 = $signed($signed((wire1250[(3'h6):(3'h6)] ?
                  ((wire1249 ?
                      reg1255 : wire1246) >= wire1250[(5'h12):(4'hc)]) : $unsigned(wire1246[(4'hf):(4'h8)]))));
              reg1254 <= $signed((8'ha6));
              reg1255 <= wire1247;
              reg1256 <= {reg1255, $unsigned(reg1253)};
            end
        end
      else
        begin
          reg1254 <= ((~&wire1250[(4'hb):(2'h3)]) ?
              $unsigned($unsigned({$signed(wire1250),
                  ((8'hae) * wire1246)})) : reg1254[(4'h8):(2'h2)]);
          reg1257 = $unsigned(wire1249);
          reg1258 <= wire1246[(3'h5):(3'h4)];
          if ((|$signed(wire1247[(2'h2):(1'h1)])))
            begin
              reg1259 <= ((+(((!reg1253) ?
                          (~^(7'h42)) : wire1251[(1'h0):(1'h0)]) ?
                      (-{reg1253,
                          (8'hb9)}) : (wire1247[(1'h1):(1'h1)] || wire1248))) ?
                  (^($signed((8'hbd)) ^~ $unsigned((wire1249 == wire1252)))) : {wire1248,
                      (^wire1249)});
            end
          else
            begin
              reg1260 = $unsigned($signed(((&reg1257) || reg1258)));
              reg1261 = $signed({$signed((-((8'hac) || wire1251))),
                  $unsigned($signed((&reg1256)))});
            end
        end
    end
  always
    @(posedge clk) begin
      reg1262 <= (reg1258 ?
          $unsigned(wire1247) : (($signed((|wire1248)) >= wire1247[(3'h4):(1'h0)]) >>> {($signed((7'h41)) ?
                  (wire1249 ? wire1251 : wire1246) : (^(7'h46)))}));
      reg1263 = $signed((~$signed(((reg1259 && wire1249) ?
          $signed(wire1248) : reg1256))));
    end
  always
    @(posedge clk) begin
      reg1264 = wire1246[(4'h8):(3'h4)];
    end
  always
    @(posedge clk) begin
      if (wire1251[(1'h1):(1'h0)])
        begin
          for (forvar1265 = (1'h0); (forvar1265 < (1'h0)); forvar1265 = (forvar1265 + (1'h1)))
            begin
              reg1266 = reg1262[(3'h4):(3'h4)];
              reg1267 = reg1262[(3'h7):(2'h3)];
              reg1268 <= $signed((($signed({wire1246, reg1255}) ?
                      wire1246 : ($signed(wire1251) ~^ $signed(forvar1265))) ?
                  $unsigned((^wire1251)) : $signed({(reg1258 ^~ reg1267)})));
              reg1269 = reg1258[(1'h1):(1'h1)];
              reg1270 <= wire1249;
            end
          if ($signed((reg1266 ?
              (8'h9c) : $unsigned({(reg1262 ? reg1258 : reg1269)}))))
            begin
              reg1271 <= {(~$signed($signed(reg1270[(5'h12):(5'h11)])))};
              reg1272 = {(-reg1269[(2'h2):(1'h0)]), (~|reg1254)};
              reg1273 <= $signed(reg1270);
            end
          else
            begin
              reg1272 = (reg1259 < $signed($signed(((^~forvar1265) ?
                  (+reg1256) : wire1247[(2'h2):(1'h1)]))));
              reg1273 <= (($signed(((+reg1259) ?
                      (8'h9f) : (reg1271 ~^ reg1270))) * (^((forvar1265 && reg1271) ?
                      $unsigned(wire1248) : $signed(wire1246)))) ?
                  reg1266[(1'h0):(1'h0)] : (-((^~(|reg1255)) ?
                      $unsigned(((8'hb0) ?
                          reg1262 : wire1250)) : {$signed(reg1255)})));
              reg1274 <= wire1246[(5'h13):(4'hd)];
              reg1275 <= {reg1269};
              reg1276 <= ({$signed($unsigned(forvar1265)),
                      (|$unsigned((wire1246 | reg1259)))} ?
                  reg1267 : ($unsigned($unsigned($unsigned(reg1274))) ?
                      {$unsigned(((7'h42) ?
                              (8'hb9) : forvar1265))} : $unsigned((reg1254 << $unsigned(reg1256)))));
            end
          for (forvar1277 = (1'h0); (forvar1277 < (2'h2)); forvar1277 = (forvar1277 + (1'h1)))
            begin
              reg1278 = reg1266;
            end
          reg1279 = $unsigned(wire1252[(1'h1):(1'h0)]);
          reg1280 <= reg1266[(1'h0):(1'h0)];
        end
      else
        begin
          reg1265 <= (~^reg1275[(2'h2):(2'h2)]);
          reg1268 <= {reg1254[(3'h4):(1'h0)], reg1273[(4'h8):(2'h2)]};
        end
      for (forvar1281 = (1'h0); (forvar1281 < (3'h4)); forvar1281 = (forvar1281 + (1'h1)))
        begin
          reg1282 = wire1248;
        end
    end
  always
    @(posedge clk) begin
      reg1283 = $signed($unsigned($unsigned(reg1280[(4'hc):(4'ha)])));
    end
  assign wire1284 = (^~$signed(wire1252));
  always
    @(posedge clk) begin
      if (((|reg1273[(2'h3):(1'h0)]) ?
          ($unsigned(($signed(wire1248) | (wire1247 - reg1273))) || $signed($unsigned($signed(reg1273)))) : ($unsigned($unsigned((reg1258 ?
                  reg1262 : reg1273))) ?
              ((reg1271[(1'h1):(1'h0)] || $unsigned(wire1248)) ?
                  $unsigned(wire1249[(4'hc):(3'h5)]) : (~|reg1275[(1'h1):(1'h0)])) : reg1258)))
        begin
          if (reg1255)
            begin
              reg1285 = ({(~|reg1255)} ?
                  reg1268 : $unsigned((reg1265[(1'h0):(1'h0)] >= $signed((~&reg1274)))));
              reg1286 <= (8'hbc);
            end
          else
            begin
              reg1285 = reg1259;
              reg1286 <= $unsigned(((+$signed((reg1255 ? (8'ha0) : reg1262))) ?
                  (wire1251 | $signed($unsigned(reg1273))) : reg1273[(4'hc):(4'h8)]));
              reg1287 <= reg1271;
            end
          reg1288 <= $signed(reg1276[(4'hc):(4'hc)]);
        end
      else
        begin
          reg1286 <= $unsigned(reg1271[(1'h0):(1'h0)]);
        end
    end
  assign wire1289 = ($signed((&((wire1249 ? reg1280 : reg1280) ~^ {reg1276}))) ?
                        {reg1254[(3'h7):(2'h3)],
                            (+wire1250)} : reg1258[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg1290 = wire1251;
      reg1291 <= $unsigned((!reg1288));
      if ((reg1290 ? $unsigned((!{reg1270[(5'h12):(3'h4)]})) : (~&wire1247)))
        begin
          reg1292 = $signed(reg1291[(4'h8):(2'h2)]);
          reg1293 <= reg1255;
          if ((-(wire1252[(5'h10):(4'h8)] | ((^reg1274[(3'h5):(2'h2)]) ?
              $signed((^~(8'ha9))) : (~reg1291)))))
            begin
              reg1294 <= ((!(-wire1249[(3'h5):(3'h4)])) ?
                  wire1250 : (^~(((+reg1288) < (reg1274 << reg1290)) ?
                      wire1250[(5'h10):(5'h10)] : $signed((reg1258 != (8'ha6))))));
              reg1295 <= ($signed({((reg1275 ?
                          (8'ha3) : reg1286) && (+reg1291))}) ?
                  ($unsigned($signed(reg1275)) ?
                      $signed((~|{reg1290,
                          reg1291})) : (reg1290[(4'hf):(1'h0)] + $signed(wire1250[(4'hd):(2'h2)]))) : reg1287[(4'hf):(3'h5)]);
            end
          else
            begin
              reg1294 <= $signed((8'ha4));
              reg1296 = $unsigned((~|(8'ha6)));
              reg1297 = (($unsigned(wire1284[(2'h2):(1'h1)]) ?
                      wire1252[(3'h5):(3'h5)] : $unsigned($unsigned(reg1268))) ?
                  ($signed(reg1280[(4'hb):(1'h0)]) == (!(8'hb7))) : $signed($unsigned(((reg1259 ?
                          reg1256 : (7'h40)) ?
                      (^~wire1247) : $signed(reg1262)))));
              reg1298 = (reg1295[(3'h5):(2'h2)] < $signed($unsigned((reg1294 < (~^reg1286)))));
              reg1299 <= $unsigned(reg1273);
            end
          for (forvar1300 = (1'h0); (forvar1300 < (3'h4)); forvar1300 = (forvar1300 + (1'h1)))
            begin
              reg1301 = (reg1280 ?
                  $unsigned(reg1256[(4'hd):(4'hb)]) : ({(-$signed(reg1286))} && (((forvar1300 ?
                              reg1265 : wire1252) ?
                          (wire1252 ? wire1246 : reg1270) : $signed(wire1250)) ?
                      reg1273[(4'h8):(3'h7)] : wire1250)));
              reg1302 <= $signed(reg1270[(4'hc):(4'hb)]);
              reg1303 <= reg1273;
              reg1304 = wire1289[(2'h2):(1'h0)];
            end
          for (forvar1305 = (1'h0); (forvar1305 < (3'h4)); forvar1305 = (forvar1305 + (1'h1)))
            begin
              reg1306 <= $unsigned((8'h9d));
            end
        end
      else
        begin
          if (((reg1256 ?
                  reg1273 : (($signed(reg1292) << reg1258[(2'h3):(2'h2)]) < wire1251)) ?
              ((8'hb5) ?
                  (-$signed($unsigned(reg1302))) : $signed(wire1249)) : wire1248))
            begin
              reg1292 = (+$unsigned(reg1268));
              reg1296 = (~&((~^forvar1305) ?
                  reg1292[(2'h3):(1'h1)] : {(((8'hbb) ?
                          wire1247 : forvar1305) | (8'ha8)),
                      $signed($unsigned(reg1299))}));
              reg1297 = ({reg1294[(3'h7):(3'h6)],
                      ((|(reg1295 >>> reg1296)) & (wire1248[(4'hd):(4'hb)] && ((8'hb9) ?
                          wire1247 : (8'ha0))))} ?
                  $unsigned(reg1292) : {$signed($signed((wire1247 ?
                          reg1274 : reg1259)))});
            end
          else
            begin
              reg1293 <= reg1291[(4'ha):(4'h8)];
              reg1294 <= ($unsigned($signed($signed((reg1294 ~^ reg1301)))) ?
                  reg1275[(3'h5):(3'h4)] : ({reg1265[(2'h2):(2'h2)]} <= $signed((!wire1250))));
            end
          for (forvar1298 = (1'h0); (forvar1298 < (3'h4)); forvar1298 = (forvar1298 + (1'h1)))
            begin
              reg1300 = forvar1305;
              reg1302 <= reg1268;
              reg1303 <= $signed(forvar1305[(5'h11):(4'hb)]);
              reg1305 <= forvar1305;
            end
          for (forvar1306 = (1'h0); (forvar1306 < (3'h4)); forvar1306 = (forvar1306 + (1'h1)))
            begin
              reg1307 <= ($unsigned({(reg1293[(1'h1):(1'h1)] >> $unsigned(reg1254))}) ?
                  wire1250[(3'h6):(3'h4)] : (wire1247 ?
                      reg1265 : reg1292[(2'h2):(1'h1)]));
              reg1308 <= $unsigned($signed(reg1296[(1'h1):(1'h0)]));
            end
          reg1309 = $signed($signed($unsigned(reg1307)));
          reg1310 = ($unsigned({$unsigned(((7'h40) ?
                  reg1306 : (8'hbb)))}) & wire1248);
        end
      reg1311 = $unsigned($signed((^reg1254)));
    end
  always
    @(posedge clk) begin
      reg1312 <= reg1288[(3'h6):(3'h4)];
      reg1313 = {reg1271, $unsigned($unsigned($unsigned($signed((8'ha1)))))};
      reg1314 = (~reg1305[(1'h0):(1'h0)]);
      reg1315 = reg1276;
      reg1316 = reg1313;
    end
  assign wire1317 = (-(~&wire1249[(2'h2):(1'h0)]));
  assign wire1318 = reg1276;
  always
    @(posedge clk) begin
      reg1319 = reg1274[(1'h0):(1'h0)];
      if ((|($unsigned({(-reg1291),
          (reg1293 * reg1254)}) < reg1276[(1'h0):(1'h0)])))
        begin
          for (forvar1320 = (1'h0); (forvar1320 < (1'h1)); forvar1320 = (forvar1320 + (1'h1)))
            begin
              reg1321 <= $unsigned({($signed(wire1249) >>> reg1294[(4'hc):(3'h4)]),
                  (~|($unsigned((7'h4a)) ?
                      {reg1274, wire1246} : (reg1305 ^~ reg1258)))});
              reg1322 = $signed(((~^((reg1262 >>> (8'hab)) <= (wire1247 >= reg1299))) ~^ $unsigned((reg1294 ^ (wire1246 <<< (8'hbd))))));
              reg1323 = (|reg1275);
              reg1324 <= {$unsigned((reg1270[(1'h1):(1'h0)] ?
                      (~^wire1251[(2'h2):(2'h2)]) : reg1255))};
            end
        end
      else
        begin
          if (reg1312[(1'h0):(1'h0)])
            begin
              reg1320 = $unsigned(($unsigned(($signed((8'ha0)) & $unsigned(reg1268))) ?
                  (|(wire1317[(3'h4):(1'h0)] ?
                      wire1318[(3'h5):(3'h5)] : (~|reg1265))) : (wire1249[(4'ha):(2'h2)] ?
                      (~$unsigned(reg1262)) : wire1318[(5'h10):(4'he)])));
              reg1322 = (~|($signed($unsigned(wire1251[(1'h0):(1'h0)])) ?
                  (^~{(reg1306 ? reg1291 : reg1324), wire1252}) : (reg1299 ?
                      (reg1273[(4'hb):(1'h1)] ?
                          {reg1303, reg1305} : {reg1254}) : $unsigned({reg1255,
                          reg1268}))));
              reg1324 <= (8'ha0);
              reg1325 = reg1288;
              reg1326 = reg1273;
            end
          else
            begin
              reg1321 <= reg1280;
              reg1322 = $signed((((^(~^reg1302)) ?
                      ((reg1255 ? reg1294 : reg1326) ?
                          reg1286[(1'h0):(1'h0)] : (reg1299 >> wire1249)) : $signed($signed(reg1303))) ?
                  reg1294[(4'hd):(4'hc)] : ((|reg1305[(4'hf):(2'h3)]) == reg1286)));
              reg1323 = (~|(|(reg1291 != $unsigned((wire1318 | reg1321)))));
              reg1324 <= $signed(($unsigned($signed((+reg1271))) >>> (!((reg1256 ?
                      wire1249 : reg1280) ?
                  wire1317[(3'h4):(3'h4)] : $signed(reg1287)))));
              reg1327 <= reg1324;
            end
          reg1328 = reg1262;
          for (forvar1329 = (1'h0); (forvar1329 < (2'h2)); forvar1329 = (forvar1329 + (1'h1)))
            begin
              reg1330 <= {((((reg1307 + (8'hb3)) ?
                          reg1302 : (|wire1249)) || $signed((reg1268 ?
                          reg1293 : reg1275))) ?
                      $signed(reg1254) : (7'h41))};
              reg1331 <= (&{{$unsigned((reg1270 >>> (8'hb6)))}});
              reg1332 = $unsigned({$signed({reg1308})});
            end
          for (forvar1333 = (1'h0); (forvar1333 < (2'h2)); forvar1333 = (forvar1333 + (1'h1)))
            begin
              reg1334 = $signed(forvar1329[(3'h6):(2'h2)]);
              reg1335 <= reg1323;
            end
        end
    end
  assign wire1336 = ($unsigned(((reg1303[(2'h3):(1'h1)] <<< $unsigned(wire1289)) > reg1330[(1'h1):(1'h0)])) ~^ ((((~|wire1284) * reg1321[(5'h11):(1'h1)]) <= $signed(wire1247)) ?
                        wire1250[(4'hc):(3'h7)] : $signed(((reg1274 & wire1246) * (reg1331 >> wire1248)))));
  assign wire1337 = reg1262;
  always
    @(posedge clk) begin
      reg1338 <= $unsigned(reg1307);
      reg1339 = reg1254[(1'h0):(1'h0)];
      if (($signed(($unsigned((reg1256 ^~ (7'h41))) ?
          reg1274 : reg1335)) < (wire1251 || wire1284)))
        begin
          if ((^$signed(($unsigned(reg1276[(3'h6):(1'h0)]) ?
              (~^reg1306) : (!(reg1268 ? wire1336 : (8'hae)))))))
            begin
              reg1340 = (wire1249 ?
                  ({($unsigned(reg1338) ?
                          (reg1327 ~^ wire1289) : $signed(reg1324))} != reg1308[(1'h0):(1'h0)]) : $signed((reg1312 | (~$unsigned((8'ha7))))));
              reg1341 <= wire1289;
              reg1342 <= ($unsigned(((~wire1251[(1'h1):(1'h0)]) == $signed(reg1256[(4'hb):(4'h9)]))) ?
                  ((8'hbd) ?
                      ((reg1270 ? (~&wire1250) : $unsigned(reg1259)) ?
                          reg1312 : {reg1258[(4'h8):(1'h0)]}) : ((reg1321[(1'h0):(1'h0)] ?
                              $signed(reg1273) : (reg1335 ^~ wire1337)) ?
                          ((-reg1287) ?
                              {reg1271,
                                  wire1336} : (wire1337 | reg1294)) : $unsigned((~reg1306)))) : (($unsigned($unsigned(reg1255)) ?
                      {(!(8'hbf))} : $unsigned($unsigned(reg1338))) == ((reg1262 ?
                          (reg1288 ?
                              wire1336 : reg1295) : (reg1280 & reg1259)) ?
                      $unsigned((~&reg1271)) : reg1303)));
              reg1343 = wire1246[(3'h4):(1'h0)];
            end
          else
            begin
              reg1341 <= ($signed($unsigned(({reg1324,
                  reg1268} << wire1289[(1'h1):(1'h1)]))) * wire1249);
            end
          reg1344 <= reg1262;
          reg1345 <= (|(reg1258[(2'h3):(1'h1)] << (-(8'h9d))));
        end
      else
        begin
          if (wire1318)
            begin
              reg1340 = $unsigned((~((-(reg1258 ?
                  reg1258 : wire1318)) << (~|(reg1265 * wire1251)))));
              reg1341 <= (wire1246 - (reg1335[(1'h0):(1'h0)] ?
                  reg1307 : reg1268));
            end
          else
            begin
              reg1341 <= reg1268[(1'h0):(1'h0)];
              reg1343 = (+reg1273);
            end
          reg1346 = (~($unsigned((reg1308 ? (^~reg1280) : {reg1338, reg1256})) ?
              (&((reg1270 != reg1259) - $signed(reg1339))) : {reg1293[(1'h1):(1'h0)]}));
          reg1347 = (~&(!$signed($signed({reg1342, reg1335}))));
          reg1348 <= $unsigned(reg1274);
        end
    end
  assign wire1349 = $signed((($signed(wire1337) << (reg1259[(4'hb):(3'h6)] ?
                        reg1345 : {reg1287, wire1252})) < $unsigned({(reg1342 ?
                            reg1305 : (7'h4a)),
                        (-(8'hac))})));
  always
    @(posedge clk) begin
      if (reg1262[(1'h1):(1'h0)])
        begin
          for (forvar1350 = (1'h0); (forvar1350 < (2'h3)); forvar1350 = (forvar1350 + (1'h1)))
            begin
              reg1351 = wire1251;
            end
          for (forvar1352 = (1'h0); (forvar1352 < (3'h4)); forvar1352 = (forvar1352 + (1'h1)))
            begin
              reg1353 = (reg1345 * (reg1330[(5'h15):(1'h1)] | {(^(reg1302 ?
                      wire1250 : (8'hb1)))}));
            end
          reg1354 = wire1248[(1'h0):(1'h0)];
          reg1355 <= (~&{($unsigned((reg1273 <= wire1251)) | (&(wire1250 ~^ reg1268))),
              reg1293[(1'h0):(1'h0)]});
          for (forvar1356 = (1'h0); (forvar1356 < (2'h2)); forvar1356 = (forvar1356 + (1'h1)))
            begin
              reg1357 <= {(^(((reg1355 << reg1327) ?
                      wire1289 : (reg1293 ?
                          reg1268 : (8'hac))) >= wire1251[(1'h1):(1'h1)])),
                  $signed($unsigned(reg1342[(1'h1):(1'h0)]))};
              reg1358 = reg1262[(4'hf):(3'h4)];
              reg1359 = ((reg1344 ?
                  {$signed($unsigned((8'hb2)))} : ({(wire1318 <= reg1276)} | ((reg1288 < (7'h48)) ?
                      reg1271 : {reg1254}))) <= (($signed({reg1255,
                      reg1348}) < (~^{(8'ha1)})) ?
                  (~({reg1335} ?
                      {reg1254} : reg1330)) : (reg1268[(2'h2):(1'h0)] ?
                      (~(7'h49)) : ($signed(wire1251) ?
                          $signed((8'hbc)) : $unsigned(reg1303)))));
              reg1360 <= (forvar1350 + ((&reg1359[(5'h16):(4'hf)]) ?
                  reg1306 : $signed((^~wire1251[(2'h2):(2'h2)]))));
              reg1361 = (|{(8'had),
                  (+($unsigned(reg1338) ?
                      (reg1274 ? reg1359 : reg1303) : reg1303))});
            end
        end
      else
        begin
          reg1350 = reg1321[(5'h10):(1'h1)];
          if ($unsigned(reg1299[(2'h2):(1'h1)]))
            begin
              reg1351 = $signed(($signed(reg1255[(2'h3):(1'h1)]) ~^ (((^~reg1268) ?
                      $signed(wire1250) : ((8'hab) ? reg1327 : reg1275)) ?
                  reg1256[(5'h16):(2'h3)] : $signed(wire1284[(3'h6):(1'h0)]))));
              reg1352 = ((&{forvar1356,
                      (reg1271[(4'h8):(1'h0)] ?
                          $unsigned(wire1251) : (reg1276 ^~ reg1335))}) ?
                  $unsigned(forvar1350[(1'h0):(1'h0)]) : (((((8'h9c) ^~ reg1348) ?
                              (wire1349 >= reg1280) : reg1342) ?
                          $unsigned(wire1317[(2'h2):(2'h2)]) : ((wire1246 ?
                              reg1353 : (8'hbb)) << (!reg1275))) ?
                      $signed(($unsigned((8'h9d)) ?
                          ((7'h48) + reg1305) : (reg1344 >= forvar1350))) : (wire1252 ?
                          $signed($signed(reg1331)) : reg1291[(2'h3):(2'h2)])));
              reg1355 <= {reg1287[(2'h3):(1'h1)]};
              reg1356 <= (~reg1254);
            end
          else
            begin
              reg1355 <= $signed((wire1337[(2'h3):(1'h1)] ?
                  wire1247[(2'h3):(1'h1)] : forvar1352[(4'hc):(4'ha)]));
            end
          reg1358 = ($signed(((reg1275[(1'h0):(1'h0)] ~^ {wire1318}) ?
                  $unsigned(wire1246[(5'h12):(4'h9)]) : $signed((reg1331 ?
                      reg1331 : (8'hb9))))) ?
              ((~|$signed({reg1348})) == ({$unsigned((8'h9c))} ?
                  ((reg1361 ? reg1306 : (8'hb4)) ?
                      reg1295[(3'h5):(3'h4)] : $unsigned(reg1344)) : (8'hba))) : reg1345[(1'h1):(1'h0)]);
          for (forvar1359 = (1'h0); (forvar1359 < (3'h4)); forvar1359 = (forvar1359 + (1'h1)))
            begin
              reg1361 = reg1331[(5'h17):(4'hf)];
              reg1362 = reg1360;
            end
        end
      if ($signed($signed((({reg1330, wire1247} ?
          (reg1265 || reg1305) : (reg1305 >>> wire1289)) > $signed(((8'hab) ?
          (8'hab) : reg1353))))))
        begin
          reg1363 = wire1251;
        end
      else
        begin
          reg1363 = $signed(reg1350[(5'h13):(3'h6)]);
          reg1364 <= (7'h42);
          reg1365 <= $unsigned($signed($unsigned(((8'h9f) ?
              $unsigned(wire1349) : $signed(reg1255)))));
          reg1366 <= (^(|$unsigned(reg1275)));
        end
      if ((!reg1356[(5'h14):(4'hb)]))
        begin
          reg1367 = wire1249;
          reg1368 <= forvar1359;
          for (forvar1369 = (1'h0); (forvar1369 < (1'h0)); forvar1369 = (forvar1369 + (1'h1)))
            begin
              reg1370 <= ((($unsigned((-wire1337)) ^ $unsigned($unsigned(reg1338))) ?
                  (-reg1276[(3'h6):(1'h1)]) : $unsigned(reg1321[(4'h9):(3'h5)])) <= (reg1355[(2'h3):(2'h3)] ?
                  (($signed(reg1262) >> wire1247) <<< (+reg1353[(1'h1):(1'h0)])) : $unsigned((!(reg1367 ?
                      reg1341 : wire1249)))));
            end
          if ((~&(~reg1259[(4'hc):(4'h9)])))
            begin
              reg1371 = ({$unsigned(reg1312),
                  $signed((reg1360[(2'h2):(1'h1)] && reg1254))} >>> (~|{(reg1360[(3'h6):(3'h4)] ^ (|reg1276)),
                  ((7'h47) ? (reg1335 ? (8'ha1) : reg1360) : (&reg1355))}));
              reg1372 <= (~&(reg1366 * ($signed($signed((8'ha3))) - wire1251)));
              reg1373 <= (wire1284[(4'hc):(3'h6)] >= (forvar1352 ?
                  (^((reg1254 ?
                      reg1356 : reg1291) || $unsigned(reg1308))) : reg1321[(5'h12):(4'hf)]));
              reg1374 = forvar1350[(1'h1):(1'h1)];
            end
          else
            begin
              reg1371 = reg1371;
            end
          reg1375 = {$unsigned($signed(reg1350)), reg1358[(2'h2):(2'h2)]};
        end
      else
        begin
          reg1367 = ({reg1321[(4'he):(4'ha)],
                  $unsigned(($unsigned(wire1289) > (reg1270 >= reg1321)))} ?
              ((7'h47) >= ((reg1321 ?
                      ((8'hba) ~^ reg1275) : (reg1303 ? wire1246 : reg1305)) ?
                  reg1280[(4'hb):(3'h5)] : ((reg1275 ?
                      reg1274 : reg1354) <<< reg1359))) : ($signed(reg1361[(3'h7):(2'h2)]) + $signed((reg1341[(1'h1):(1'h1)] ^~ wire1252))));
          reg1369 = ($signed((((wire1251 ? (8'hb4) : reg1370) ?
                  {reg1331} : (reg1268 ? (8'h9d) : reg1355)) && (reg1295 ?
                  reg1303 : (~reg1306)))) ?
              $unsigned(((reg1302[(1'h1):(1'h0)] < reg1270) ?
                  {$signed(reg1371),
                      reg1302[(4'h9):(2'h3)]} : (|(~^reg1312)))) : reg1268[(2'h2):(2'h2)]);
          for (forvar1370 = (1'h0); (forvar1370 < (2'h2)); forvar1370 = (forvar1370 + (1'h1)))
            begin
              reg1372 <= {forvar1370[(4'h8):(3'h7)], reg1280};
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module901
#(parameter param1242 = ((^(8'hbd)) ? (&(({(8'hb3)} || ((8'hb4) >>> (7'h41))) ? ((8'hb1) ? ((8'haa) ? (8'hbd) : (7'h47)) : {(8'h9d)}) : (&((8'hba) ? (8'hab) : (8'haa))))) : {(&(((7'h46) < (8'hbc)) ? {(8'hb0)} : (8'ha9)))}))
(y, clk, wire906, wire905, wire904, wire903, wire902);
  output wire [(32'h11b4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire906;
  input wire signed [(5'h17):(1'h0)] wire905;
  input wire [(4'hc):(1'h0)] wire904;
  input wire signed [(4'he):(1'h0)] wire903;
  input wire signed [(2'h2):(1'h0)] wire902;
  wire [(5'h18):(1'h0)] wire1220;
  wire [(3'h4):(1'h0)] wire1182;
  wire signed [(3'h4):(1'h0)] wire1181;
  wire signed [(3'h7):(1'h0)] wire1180;
  wire [(4'ha):(1'h0)] wire1179;
  wire [(4'he):(1'h0)] wire1178;
  wire signed [(2'h2):(1'h0)] wire1177;
  wire signed [(2'h3):(1'h0)] wire1153;
  wire [(2'h3):(1'h0)] wire1104;
  wire [(4'h8):(1'h0)] wire1103;
  wire signed [(2'h2):(1'h0)] wire1102;
  wire signed [(2'h3):(1'h0)] wire1101;
  wire [(5'h18):(1'h0)] wire1100;
  wire [(4'h8):(1'h0)] wire986;
  wire signed [(4'hc):(1'h0)] wire929;
  reg [(2'h3):(1'h0)] reg1240 = (1'h0);
  reg [(5'h11):(1'h0)] reg1238 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1237 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1236 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1234 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1232 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1230 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1228 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1226 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1224 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1222 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1219 = (1'h0);
  reg [(4'hc):(1'h0)] reg1218 = (1'h0);
  reg [(5'h11):(1'h0)] reg1216 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1214 = (1'h0);
  reg [(4'he):(1'h0)] reg1212 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1211 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1208 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1205 = (1'h0);
  reg [(4'he):(1'h0)] reg1202 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1200 = (1'h0);
  reg [(5'h13):(1'h0)] reg1196 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1194 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1192 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1188 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1186 = (1'h0);
  reg [(4'h8):(1'h0)] reg1185 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1173 = (1'h0);
  reg [(4'ha):(1'h0)] reg1170 = (1'h0);
  reg [(5'h18):(1'h0)] reg1168 = (1'h0);
  reg [(5'h10):(1'h0)] reg1166 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1165 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1164 = (1'h0);
  reg [(4'ha):(1'h0)] reg1163 = (1'h0);
  reg [(5'h11):(1'h0)] reg1161 = (1'h0);
  reg [(4'hf):(1'h0)] reg1155 = (1'h0);
  reg [(2'h3):(1'h0)] reg1154 = (1'h0);
  reg [(5'h15):(1'h0)] reg1152 = (1'h0);
  reg [(3'h4):(1'h0)] reg1151 = (1'h0);
  reg [(3'h5):(1'h0)] reg1146 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1144 = (1'h0);
  reg [(4'hd):(1'h0)] reg1141 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1139 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1137 = (1'h0);
  reg [(3'h5):(1'h0)] reg1136 = (1'h0);
  reg [(4'h9):(1'h0)] reg1133 = (1'h0);
  reg [(5'h13):(1'h0)] reg1132 = (1'h0);
  reg [(4'hb):(1'h0)] reg1130 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1129 = (1'h0);
  reg [(4'hf):(1'h0)] reg1124 = (1'h0);
  reg [(4'hc):(1'h0)] reg1122 = (1'h0);
  reg [(3'h6):(1'h0)] reg1119 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1116 = (1'h0);
  reg [(5'h13):(1'h0)] reg1113 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1111 = (1'h0);
  reg [(4'h8):(1'h0)] reg1109 = (1'h0);
  reg [(3'h7):(1'h0)] reg1105 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1099 = (1'h0);
  reg [(3'h5):(1'h0)] reg1097 = (1'h0);
  reg [(5'h15):(1'h0)] reg1096 = (1'h0);
  reg [(4'hf):(1'h0)] reg1094 = (1'h0);
  reg [(3'h4):(1'h0)] reg1093 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1090 = (1'h0);
  reg [(4'he):(1'h0)] reg1087 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1080 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1079 = (1'h0);
  reg [(4'hb):(1'h0)] reg1075 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1073 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1071 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1069 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1063 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1056 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1065 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1064 = (1'h0);
  reg [(4'hc):(1'h0)] reg1061 = (1'h0);
  reg [(5'h18):(1'h0)] reg1059 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1058 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1057 = (1'h0);
  reg [(5'h16):(1'h0)] reg1054 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1053 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1047 = (1'h0);
  reg [(4'h9):(1'h0)] reg1045 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1044 = (1'h0);
  reg [(4'he):(1'h0)] reg1041 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1040 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1039 = (1'h0);
  reg [(3'h6):(1'h0)] reg1036 = (1'h0);
  reg [(4'hd):(1'h0)] reg1033 = (1'h0);
  reg [(4'hd):(1'h0)] reg1031 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1030 = (1'h0);
  reg [(3'h4):(1'h0)] reg1028 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1027 = (1'h0);
  reg [(5'h11):(1'h0)] reg1024 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1022 = (1'h0);
  reg [(4'h9):(1'h0)] reg1020 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1018 = (1'h0);
  reg [(3'h5):(1'h0)] reg1017 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1016 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1014 = (1'h0);
  reg [(4'hd):(1'h0)] reg1013 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1009 = (1'h0);
  reg [(5'h14):(1'h0)] reg1008 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1005 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1002 = (1'h0);
  reg [(4'ha):(1'h0)] reg998 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg997 = (1'h0);
  reg [(5'h12):(1'h0)] reg994 = (1'h0);
  reg signed [(4'he):(1'h0)] reg992 = (1'h0);
  reg [(2'h3):(1'h0)] reg989 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg988 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg984 = (1'h0);
  reg [(3'h6):(1'h0)] reg981 = (1'h0);
  reg [(4'h8):(1'h0)] reg979 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg977 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg976 = (1'h0);
  reg [(2'h2):(1'h0)] reg975 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg974 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg971 = (1'h0);
  reg [(2'h2):(1'h0)] reg968 = (1'h0);
  reg [(4'h8):(1'h0)] reg967 = (1'h0);
  reg [(3'h5):(1'h0)] reg965 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg963 = (1'h0);
  reg [(3'h4):(1'h0)] reg962 = (1'h0);
  reg [(5'h17):(1'h0)] reg961 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg960 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg957 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg956 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg955 = (1'h0);
  reg [(5'h11):(1'h0)] reg952 = (1'h0);
  reg [(5'h13):(1'h0)] reg950 = (1'h0);
  reg [(4'hb):(1'h0)] reg949 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg948 = (1'h0);
  reg [(4'hb):(1'h0)] reg947 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg945 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg930 = (1'h0);
  reg [(4'hb):(1'h0)] reg941 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg936 = (1'h0);
  reg [(5'h13):(1'h0)] reg935 = (1'h0);
  reg [(3'h6):(1'h0)] reg933 = (1'h0);
  reg [(3'h5):(1'h0)] reg932 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg931 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg927 = (1'h0);
  reg [(5'h10):(1'h0)] reg926 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg924 = (1'h0);
  reg [(4'ha):(1'h0)] reg922 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg921 = (1'h0);
  reg [(4'he):(1'h0)] reg918 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg916 = (1'h0);
  reg [(3'h5):(1'h0)] reg915 = (1'h0);
  reg [(4'he):(1'h0)] reg914 = (1'h0);
  reg [(5'h16):(1'h0)] reg912 = (1'h0);
  reg [(5'h15):(1'h0)] reg911 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg910 = (1'h0);
  reg [(2'h3):(1'h0)] reg1241 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1239 = (1'h0);
  reg [(5'h18):(1'h0)] reg1235 = (1'h0);
  reg [(4'h8):(1'h0)] reg1233 = (1'h0);
  reg [(5'h11):(1'h0)] reg1231 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1229 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1227 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1225 = (1'h0);
  reg [(2'h2):(1'h0)] reg1223 = (1'h0);
  reg [(4'he):(1'h0)] forvar1221 = (1'h0);
  reg [(4'ha):(1'h0)] reg1217 = (1'h0);
  reg [(5'h13):(1'h0)] reg1215 = (1'h0);
  reg [(5'h18):(1'h0)] reg1213 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1210 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1209 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1207 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1206 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1204 = (1'h0);
  reg [(5'h18):(1'h0)] reg1203 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1201 = (1'h0);
  reg [(5'h13):(1'h0)] reg1199 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1198 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1197 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1195 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1193 = (1'h0);
  reg [(5'h13):(1'h0)] reg1191 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1190 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1189 = (1'h0);
  reg [(5'h12):(1'h0)] reg1187 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1184 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1183 = (1'h0);
  reg [(2'h3):(1'h0)] reg1176 = (1'h0);
  reg [(5'h15):(1'h0)] reg1175 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1174 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1172 = (1'h0);
  reg [(5'h11):(1'h0)] reg1171 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1169 = (1'h0);
  reg [(4'ha):(1'h0)] reg1167 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1162 = (1'h0);
  reg [(3'h6):(1'h0)] reg1160 = (1'h0);
  reg [(4'hd):(1'h0)] reg1159 = (1'h0);
  reg [(3'h5):(1'h0)] reg1158 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1157 = (1'h0);
  reg [(4'hc):(1'h0)] reg1156 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1149 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1148 = (1'h0);
  reg [(3'h5):(1'h0)] reg1147 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1145 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1143 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1142 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1134 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1131 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1138 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1135 = (1'h0);
  reg [(5'h16):(1'h0)] reg1134 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1131 = (1'h0);
  reg [(4'h9):(1'h0)] reg1128 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1127 = (1'h0);
  reg [(5'h15):(1'h0)] reg1126 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1125 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1123 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1121 = (1'h0);
  reg [(4'hd):(1'h0)] reg1120 = (1'h0);
  reg [(3'h5):(1'h0)] reg1118 = (1'h0);
  reg [(5'h18):(1'h0)] reg1117 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1115 = (1'h0);
  reg [(5'h13):(1'h0)] reg1114 = (1'h0);
  reg [(4'he):(1'h0)] reg1112 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1110 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1108 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1107 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1106 = (1'h0);
  reg [(3'h4):(1'h0)] reg1098 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1095 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1092 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1091 = (1'h0);
  reg [(3'h4):(1'h0)] reg1081 = (1'h0);
  reg [(4'hd):(1'h0)] reg1072 = (1'h0);
  reg [(4'hb):(1'h0)] reg1089 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1088 = (1'h0);
  reg [(5'h15):(1'h0)] reg1086 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1085 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1084 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1083 = (1'h0);
  reg [(4'hb):(1'h0)] reg1082 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1081 = (1'h0);
  reg [(4'ha):(1'h0)] reg1078 = (1'h0);
  reg [(5'h18):(1'h0)] reg1077 = (1'h0);
  reg [(3'h7):(1'h0)] reg1076 = (1'h0);
  reg [(3'h7):(1'h0)] reg1074 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1072 = (1'h0);
  reg [(3'h6):(1'h0)] reg1070 = (1'h0);
  reg [(4'h9):(1'h0)] reg1068 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1067 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1065 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1066 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1063 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1062 = (1'h0);
  reg [(5'h17):(1'h0)] reg1060 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1056 = (1'h0);
  reg [(4'h9):(1'h0)] reg1055 = (1'h0);
  reg [(5'h18):(1'h0)] reg1052 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1051 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1049 = (1'h0);
  reg [(5'h10):(1'h0)] reg1048 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1046 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1043 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1042 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1038 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1037 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1035 = (1'h0);
  reg [(5'h13):(1'h0)] reg1034 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1032 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1029 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1026 = (1'h0);
  reg [(5'h14):(1'h0)] reg1026 = (1'h0);
  reg [(5'h11):(1'h0)] reg1025 = (1'h0);
  reg [(4'hf):(1'h0)] reg1023 = (1'h0);
  reg [(4'hf):(1'h0)] reg1021 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1019 = (1'h0);
  reg [(3'h5):(1'h0)] reg1015 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1012 = (1'h0);
  reg [(5'h18):(1'h0)] reg1010 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1007 = (1'h0);
  reg [(3'h6):(1'h0)] reg1006 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1004 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1003 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1001 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg995 = (1'h0);
  reg [(2'h3):(1'h0)] reg993 = (1'h0);
  reg [(4'hf):(1'h0)] forvar992 = (1'h0);
  reg [(2'h2):(1'h0)] reg991 = (1'h0);
  reg [(5'h15):(1'h0)] reg987 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1000 = (1'h0);
  reg [(5'h10):(1'h0)] reg999 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg996 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar995 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar993 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar991 = (1'h0);
  reg [(3'h5):(1'h0)] reg990 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar987 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg985 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar983 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg982 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg980 = (1'h0);
  reg [(3'h6):(1'h0)] reg978 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar973 = (1'h0);
  reg [(3'h5):(1'h0)] reg972 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg970 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar969 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg966 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg964 = (1'h0);
  reg [(5'h11):(1'h0)] forvar956 = (1'h0);
  reg [(5'h10):(1'h0)] reg953 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg959 = (1'h0);
  reg [(3'h6):(1'h0)] reg958 = (1'h0);
  reg [(3'h7):(1'h0)] reg954 = (1'h0);
  reg [(4'h8):(1'h0)] forvar953 = (1'h0);
  reg [(4'h9):(1'h0)] reg951 = (1'h0);
  reg [(5'h15):(1'h0)] reg946 = (1'h0);
  reg [(3'h5):(1'h0)] reg944 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg943 = (1'h0);
  reg [(2'h2):(1'h0)] forvar939 = (1'h0);
  reg [(4'hf):(1'h0)] reg937 = (1'h0);
  reg [(4'h9):(1'h0)] reg942 = (1'h0);
  reg [(5'h18):(1'h0)] reg940 = (1'h0);
  reg signed [(4'he):(1'h0)] reg939 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg938 = (1'h0);
  reg [(5'h17):(1'h0)] forvar937 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg934 = (1'h0);
  reg [(2'h2):(1'h0)] forvar930 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg928 = (1'h0);
  reg [(5'h11):(1'h0)] forvar921 = (1'h0);
  reg [(5'h18):(1'h0)] reg920 = (1'h0);
  reg [(4'hf):(1'h0)] reg925 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg923 = (1'h0);
  reg [(5'h15):(1'h0)] forvar920 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg919 = (1'h0);
  reg [(5'h10):(1'h0)] reg917 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg913 = (1'h0);
  reg [(4'h8):(1'h0)] forvar909 = (1'h0);
  reg [(4'hd):(1'h0)] reg908 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg907 = (1'h0);
  assign y = {wire1220,
                 wire1182,
                 wire1181,
                 wire1180,
                 wire1179,
                 wire1178,
                 wire1177,
                 wire1153,
                 wire1104,
                 wire1103,
                 wire1102,
                 wire1101,
                 wire1100,
                 wire986,
                 wire929,
                 reg1240,
                 reg1238,
                 reg1237,
                 reg1236,
                 reg1234,
                 reg1232,
                 reg1230,
                 reg1228,
                 reg1226,
                 reg1224,
                 reg1222,
                 reg1219,
                 reg1218,
                 reg1216,
                 reg1214,
                 reg1212,
                 reg1211,
                 reg1208,
                 reg1205,
                 reg1202,
                 reg1200,
                 reg1196,
                 reg1194,
                 reg1192,
                 reg1188,
                 reg1186,
                 reg1185,
                 reg1173,
                 reg1170,
                 reg1168,
                 reg1166,
                 reg1165,
                 reg1164,
                 reg1163,
                 reg1161,
                 reg1155,
                 reg1154,
                 reg1152,
                 reg1151,
                 reg1146,
                 reg1144,
                 reg1141,
                 reg1139,
                 reg1137,
                 reg1136,
                 reg1133,
                 reg1132,
                 reg1130,
                 reg1129,
                 reg1124,
                 reg1122,
                 reg1119,
                 reg1116,
                 reg1113,
                 reg1111,
                 reg1109,
                 reg1105,
                 reg1099,
                 reg1097,
                 reg1096,
                 reg1094,
                 reg1093,
                 reg1090,
                 reg1087,
                 reg1080,
                 reg1079,
                 reg1075,
                 reg1073,
                 reg1071,
                 reg1069,
                 reg1063,
                 reg1056,
                 reg1065,
                 reg1064,
                 reg1061,
                 reg1059,
                 reg1058,
                 reg1057,
                 reg1054,
                 reg1053,
                 reg1050,
                 reg1047,
                 reg1045,
                 reg1044,
                 reg1041,
                 reg1040,
                 reg1039,
                 reg1036,
                 reg1033,
                 reg1031,
                 reg1030,
                 reg1028,
                 reg1027,
                 reg1024,
                 reg1022,
                 reg1020,
                 reg1018,
                 reg1017,
                 reg1016,
                 reg1014,
                 reg1013,
                 reg1011,
                 reg1009,
                 reg1008,
                 reg1005,
                 reg1002,
                 reg998,
                 reg997,
                 reg994,
                 reg992,
                 reg989,
                 reg988,
                 reg984,
                 reg981,
                 reg979,
                 reg977,
                 reg976,
                 reg975,
                 reg974,
                 reg971,
                 reg968,
                 reg967,
                 reg965,
                 reg963,
                 reg962,
                 reg961,
                 reg960,
                 reg957,
                 reg956,
                 reg955,
                 reg952,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 reg945,
                 reg930,
                 reg941,
                 reg936,
                 reg935,
                 reg933,
                 reg932,
                 reg931,
                 reg927,
                 reg926,
                 reg924,
                 reg922,
                 reg921,
                 reg918,
                 reg916,
                 reg915,
                 reg914,
                 reg912,
                 reg911,
                 reg910,
                 reg1241,
                 reg1239,
                 reg1235,
                 reg1233,
                 reg1231,
                 forvar1229,
                 reg1227,
                 reg1225,
                 reg1223,
                 forvar1221,
                 reg1217,
                 reg1215,
                 reg1213,
                 forvar1210,
                 forvar1209,
                 reg1207,
                 forvar1206,
                 reg1204,
                 reg1203,
                 forvar1201,
                 reg1199,
                 reg1198,
                 reg1197,
                 forvar1195,
                 reg1193,
                 reg1191,
                 forvar1190,
                 forvar1189,
                 reg1187,
                 forvar1184,
                 forvar1183,
                 reg1176,
                 reg1175,
                 reg1174,
                 reg1172,
                 reg1171,
                 reg1169,
                 reg1167,
                 reg1162,
                 reg1160,
                 reg1159,
                 reg1158,
                 reg1157,
                 reg1156,
                 reg1150,
                 forvar1149,
                 reg1148,
                 reg1147,
                 forvar1145,
                 forvar1143,
                 reg1142,
                 forvar1134,
                 forvar1131,
                 reg1140,
                 reg1138,
                 reg1135,
                 reg1134,
                 reg1131,
                 reg1128,
                 reg1127,
                 reg1126,
                 reg1125,
                 reg1123,
                 reg1121,
                 reg1120,
                 reg1118,
                 reg1117,
                 forvar1115,
                 reg1114,
                 reg1112,
                 reg1110,
                 reg1108,
                 forvar1107,
                 reg1106,
                 reg1098,
                 reg1095,
                 reg1092,
                 forvar1091,
                 reg1081,
                 reg1072,
                 reg1089,
                 reg1088,
                 reg1086,
                 reg1085,
                 reg1084,
                 reg1083,
                 reg1082,
                 forvar1081,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1074,
                 forvar1072,
                 reg1070,
                 reg1068,
                 reg1067,
                 forvar1065,
                 reg1066,
                 forvar1063,
                 reg1062,
                 reg1060,
                 forvar1056,
                 reg1055,
                 reg1052,
                 reg1051,
                 reg1049,
                 reg1048,
                 reg1046,
                 forvar1043,
                 reg1042,
                 forvar1038,
                 reg1037,
                 forvar1035,
                 reg1034,
                 reg1032,
                 reg1029,
                 forvar1026,
                 reg1026,
                 reg1025,
                 reg1023,
                 reg1021,
                 reg1019,
                 reg1015,
                 reg1012,
                 reg1010,
                 reg1007,
                 reg1006,
                 reg1004,
                 forvar1003,
                 forvar1001,
                 reg995,
                 reg993,
                 forvar992,
                 reg991,
                 reg987,
                 reg1000,
                 reg999,
                 reg996,
                 forvar995,
                 forvar993,
                 forvar991,
                 reg990,
                 forvar987,
                 reg985,
                 forvar983,
                 reg982,
                 reg980,
                 reg978,
                 forvar973,
                 reg972,
                 reg970,
                 forvar969,
                 reg966,
                 reg964,
                 forvar956,
                 reg953,
                 reg959,
                 reg958,
                 reg954,
                 forvar953,
                 reg951,
                 reg946,
                 reg944,
                 reg943,
                 forvar939,
                 reg937,
                 reg942,
                 reg940,
                 reg939,
                 reg938,
                 forvar937,
                 reg934,
                 forvar930,
                 reg928,
                 forvar921,
                 reg920,
                 reg925,
                 reg923,
                 forvar920,
                 reg919,
                 reg917,
                 reg913,
                 forvar909,
                 reg908,
                 reg907,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg907 = (&(&(~wire902)));
      reg908 = wire902;
    end
  always
    @(posedge clk) begin
      for (forvar909 = (1'h0); (forvar909 < (2'h3)); forvar909 = (forvar909 + (1'h1)))
        begin
          if ((~&(|$unsigned($unsigned((wire902 ? forvar909 : (8'ha3)))))))
            begin
              reg910 <= $unsigned((wire904[(4'hb):(4'h9)] || (~|$signed(wire906))));
            end
          else
            begin
              reg910 <= $unsigned(wire903);
              reg911 <= $unsigned($unsigned((~$signed(wire904))));
              reg912 <= (-(^~(~(~|wire906))));
              reg913 = (8'hb1);
            end
        end
      reg914 <= $signed((-reg913[(3'h4):(3'h4)]));
      reg915 <= reg913;
      reg916 <= reg912[(3'h6):(3'h4)];
      if ($signed((wire902[(1'h1):(1'h0)] > {((reg912 ? reg916 : reg912) ?
              ((8'hbe) <<< reg915) : $signed(wire903)),
          $unsigned($unsigned(wire904))})))
        begin
          if ($unsigned($signed({$signed((reg916 == reg915))})))
            begin
              reg917 = (~&$signed(((|$signed(reg910)) <= wire902[(1'h0):(1'h0)])));
              reg918 <= reg916[(4'hf):(2'h2)];
            end
          else
            begin
              reg918 <= $signed((forvar909[(3'h6):(1'h1)] <<< ($unsigned(reg913) ?
                  ((&wire902) >= $signed(reg913)) : (reg915[(1'h0):(1'h0)] ?
                      $signed(reg915) : wire905[(3'h7):(3'h6)]))));
              reg919 = ($signed({$signed(reg914)}) ?
                  ($signed($unsigned($signed((8'hbc)))) ?
                      (~|reg913[(1'h0):(1'h0)]) : ((-forvar909) ?
                          $signed({reg912}) : (^$signed(reg912)))) : $unsigned(({(reg912 + wire904)} <<< {reg916[(4'hf):(1'h1)]})));
            end
          for (forvar920 = (1'h0); (forvar920 < (2'h3)); forvar920 = (forvar920 + (1'h1)))
            begin
              reg921 <= (~(^~$signed((reg910 - $signed(forvar909)))));
              reg922 <= $unsigned(forvar909);
              reg923 = reg912[(1'h1):(1'h1)];
              reg924 <= $signed($unsigned((~^(-$signed((8'hb4))))));
              reg925 = $unsigned($signed($signed({reg912,
                  reg916[(5'h11):(3'h4)]})));
            end
        end
      else
        begin
          reg917 = {((($signed(reg917) ? reg910 : $unsigned(reg923)) ?
                      (~&(&wire904)) : reg911) ?
                  (+$unsigned((|reg923))) : wire903)};
          reg919 = (|$signed($unsigned({$signed(forvar909),
              $unsigned(reg912)})));
          reg920 = ({(wire903[(4'ha):(3'h6)] ?
                  reg923 : $unsigned((reg922 ? reg921 : wire905))),
              $signed(reg913[(4'h9):(4'h9)])} << (~|reg919[(3'h4):(3'h4)]));
          for (forvar921 = (1'h0); (forvar921 < (1'h1)); forvar921 = (forvar921 + (1'h1)))
            begin
              reg923 = reg912[(2'h3):(1'h0)];
              reg925 = $unsigned({reg917,
                  ($unsigned(forvar921) ?
                      reg912 : ({wire905, reg919} ?
                          {reg914} : (reg923 ? reg911 : wire903)))});
              reg926 <= $unsigned($signed(($signed((8'h9d)) ?
                  reg919[(1'h1):(1'h0)] : ($signed((7'h46)) >>> reg913))));
              reg927 <= forvar909[(1'h0):(1'h0)];
              reg928 = $signed((forvar920[(3'h7):(2'h3)] ?
                  (^(&forvar909)) : $unsigned({(^~reg918),
                      $unsigned(reg925)})));
            end
        end
    end
  assign wire929 = wire904;
  always
    @(posedge clk) begin
      if ($signed({(-(~^(wire906 ? reg914 : reg924))),
          ($signed($signed(reg924)) | reg910[(3'h6):(3'h4)])}))
        begin
          for (forvar930 = (1'h0); (forvar930 < (2'h3)); forvar930 = (forvar930 + (1'h1)))
            begin
              reg931 <= (~|$signed((((~|reg915) ?
                  $unsigned(reg918) : {reg910}) <<< $signed($unsigned(wire905)))));
              reg932 <= reg912;
              reg933 <= {(|(|(-$unsigned(reg910))))};
              reg934 = ($signed(($signed((~^wire904)) ?
                  reg932 : reg931[(3'h4):(1'h0)])) < $unsigned(reg914[(4'h8):(3'h5)]));
              reg935 <= $signed((8'ha5));
            end
          reg936 <= {(&(~^((reg926 ? reg933 : reg926) <= {reg918}))),
              (&{$signed((forvar930 + reg910))})};
          for (forvar937 = (1'h0); (forvar937 < (2'h2)); forvar937 = (forvar937 + (1'h1)))
            begin
              reg938 = $signed((wire904[(3'h5):(3'h4)] | ($unsigned((reg921 ?
                  (8'ha5) : reg927)) || {(forvar937 ? wire929 : reg921),
                  (~&reg921)})));
              reg939 = $signed($signed((&(~^wire903))));
              reg940 = wire905[(1'h0):(1'h0)];
              reg941 <= $unsigned(((({reg934} ?
                      (~^(8'ha4)) : (^~reg912)) >> $signed((reg915 ?
                      reg918 : wire905))) ?
                  $signed((|(reg922 ?
                      reg934 : reg934))) : $signed(($unsigned(reg915) << reg915[(1'h0):(1'h0)]))));
            end
          reg942 = ($unsigned((((wire904 > (8'ha1)) >= $unsigned(wire906)) < $unsigned((7'h40)))) ?
              (reg910[(3'h7):(1'h1)] != $signed($signed(reg914[(1'h0):(1'h0)]))) : $signed((wire906 ?
                  $signed((reg935 ?
                      reg914 : reg935)) : reg927[(1'h1):(1'h0)])));
        end
      else
        begin
          if ((-reg932[(2'h2):(1'h0)]))
            begin
              reg930 <= (((((reg934 * reg934) ?
                      $signed(reg918) : (reg911 ~^ reg938)) + $unsigned($signed(wire905))) ?
                  (8'haf) : reg916[(5'h10):(4'he)]) < (|(($unsigned(reg914) ?
                      $unsigned(reg921) : ((8'hb2) ? forvar937 : reg942)) ?
                  (reg922[(1'h0):(1'h0)] ?
                      (wire906 > reg915) : reg912[(4'he):(4'hb)]) : ((wire903 | reg936) ?
                      $unsigned(reg936) : $signed(reg933)))));
              reg934 = wire902;
              reg937 = wire906[(4'h8):(3'h6)];
              reg938 = (~&{reg942});
            end
          else
            begin
              reg930 <= (7'h48);
              reg931 <= $unsigned((7'h45));
              reg932 <= $signed($signed((wire902[(1'h1):(1'h0)] ?
                  ((reg912 ^ reg912) ?
                      reg934 : {reg916,
                          wire906}) : ($unsigned((8'hae)) > {reg938}))));
              reg934 = ((+($unsigned(reg924) < reg934)) - (^(~|((reg937 ?
                      wire929 : wire903) ?
                  (8'haa) : {reg934, reg941}))));
              reg937 = {wire905, $signed((+$signed(((8'hba) ^~ reg916))))};
            end
          for (forvar939 = (1'h0); (forvar939 < (2'h2)); forvar939 = (forvar939 + (1'h1)))
            begin
              reg940 = reg912[(4'h8):(3'h5)];
              reg942 = $signed(reg936);
            end
          reg943 = $unsigned(reg910[(2'h3):(1'h0)]);
          reg944 = $unsigned($unsigned($signed((^~reg918))));
          reg945 <= {(($unsigned($unsigned(wire906)) >> $unsigned(reg938[(4'h9):(3'h7)])) ?
                  {reg942[(3'h7):(2'h2)],
                      (forvar939[(1'h1):(1'h0)] <= reg910)} : $signed({forvar930[(1'h0):(1'h0)],
                      {reg937, reg934}}))};
        end
      if ((~reg924))
        begin
          reg946 = ((~&$unsigned(($unsigned(forvar937) ?
                  (reg939 ? reg935 : wire904) : $unsigned(reg921)))) ?
              (8'hb6) : $unsigned((-($unsigned(reg930) ?
                  (7'h48) : wire904[(1'h0):(1'h0)]))));
        end
      else
        begin
          reg947 <= wire903[(4'hc):(4'h9)];
          if ($signed($unsigned((($unsigned((7'h43)) ? reg935 : (^~reg912)) ?
              $unsigned($signed(reg943)) : (8'ha7)))))
            begin
              reg948 <= {(^~(~|$unsigned(reg935[(5'h12):(3'h5)]))),
                  reg918[(4'ha):(3'h5)]};
              reg949 <= $signed(($unsigned(reg916[(4'hb):(4'h8)]) ?
                  $signed((-reg927)) : reg940[(5'h13):(2'h3)]));
              reg950 <= wire929[(4'hb):(3'h6)];
              reg951 = $signed(((reg939 ?
                  (^$unsigned(wire929)) : reg921[(1'h1):(1'h1)]) != (~&(~|reg933))));
            end
          else
            begin
              reg951 = (|{($signed(wire905) || $signed((reg926 << wire903))),
                  $unsigned($signed(reg914))});
              reg952 <= reg942;
            end
        end
      if ((~&(((reg940 ?
              $unsigned(forvar937) : reg910[(1'h1):(1'h1)]) | reg939) ?
          reg911[(1'h1):(1'h0)] : (reg914 >> reg926[(4'h8):(3'h5)]))))
        begin
          for (forvar953 = (1'h0); (forvar953 < (1'h1)); forvar953 = (forvar953 + (1'h1)))
            begin
              reg954 = ($signed(forvar930) << ($signed((reg948 != {forvar939})) ?
                  ((^$signed(forvar939)) ^ (^(reg935 ?
                      reg949 : (7'h45)))) : (&$signed({wire904}))));
              reg955 <= reg932[(1'h0):(1'h0)];
            end
          if ((($signed(reg911) ?
              $signed(((reg947 ? reg922 : (8'hb3)) != (reg951 ?
                  reg934 : reg930))) : {$signed(reg910),
                  reg910[(1'h0):(1'h0)]}) + ((reg934 ^ $unsigned((forvar953 ?
                  (8'haa) : reg938))) ?
              ((+$unsigned(reg952)) ?
                  $unsigned((forvar953 ?
                      reg946 : reg948)) : ((+reg921) + reg943[(4'h8):(2'h2)])) : ((^~(-wire904)) ?
                  reg946[(5'h14):(1'h1)] : ({reg921, reg931} ?
                      (8'ha5) : (~^(8'hb9)))))))
            begin
              reg956 <= reg910[(3'h5):(2'h2)];
              reg957 <= reg951;
            end
          else
            begin
              reg958 = $signed(wire906[(3'h7):(3'h5)]);
            end
          reg959 = (&$unsigned($signed($signed((^~wire903)))));
          reg960 <= ({$unsigned(((|reg956) ?
                      $signed(reg914) : reg926[(4'hf):(1'h0)])),
                  wire904[(4'h9):(4'h8)]} ?
              $unsigned(reg927[(2'h2):(2'h2)]) : (reg934 != (8'hb6)));
        end
      else
        begin
          reg953 = $unsigned({{((reg931 || reg936) ?
                      $signed(wire902) : (reg956 ? reg942 : reg952)),
                  ($unsigned(reg918) ? (-reg936) : wire906[(3'h4):(3'h4)])}});
          reg955 <= (reg947[(1'h1):(1'h1)] ?
              $unsigned($signed((~&$unsigned(reg910)))) : $signed($unsigned($signed((reg921 ?
                  reg932 : reg946)))));
          for (forvar956 = (1'h0); (forvar956 < (2'h3)); forvar956 = (forvar956 + (1'h1)))
            begin
              reg957 <= forvar953;
              reg958 = $signed($signed(reg924));
              reg960 <= ((($unsigned($unsigned(reg960)) > $unsigned(reg931)) ^ ((~$unsigned(forvar956)) - ($signed(reg950) ?
                  $signed((8'ha2)) : {reg935}))) * (|(reg949[(4'ha):(4'h9)] ?
                  $signed((!reg939)) : reg949)));
              reg961 <= $signed((^((&(|(8'ha4))) + reg926)));
            end
          if ((wire903[(4'hb):(1'h0)] ?
              reg939[(4'he):(2'h2)] : ((reg961[(1'h0):(1'h0)] & $unsigned((reg915 ?
                      (7'h46) : wire906))) ?
                  (^$unsigned(forvar939)) : $signed($signed({reg935})))))
            begin
              reg962 <= (8'ha5);
              reg963 <= ($unsigned((7'h43)) ? reg916 : reg962);
            end
          else
            begin
              reg964 = reg955;
              reg965 <= ($unsigned((({reg945,
                  reg933} & wire903[(3'h6):(1'h0)]) - reg932[(1'h0):(1'h0)])) | reg964[(1'h0):(1'h0)]);
              reg966 = $signed(reg942);
              reg967 <= reg966[(4'he):(2'h3)];
            end
        end
      reg968 <= $signed((((7'h4a) * $unsigned((reg918 ^~ reg964))) ?
          reg953 : reg924));
      for (forvar969 = (1'h0); (forvar969 < (3'h4)); forvar969 = (forvar969 + (1'h1)))
        begin
          if (((&(~&(8'hb5))) >= {$signed((reg965[(3'h4):(1'h1)] ?
                  reg943 : (reg934 ? reg937 : reg935))),
              reg965[(3'h5):(2'h3)]}))
            begin
              reg970 = reg933[(1'h0):(1'h0)];
              reg971 <= (~|reg964[(1'h0):(1'h0)]);
              reg972 = $signed((~(8'hae)));
            end
          else
            begin
              reg970 = (+reg940[(5'h18):(1'h1)]);
            end
          for (forvar973 = (1'h0); (forvar973 < (1'h1)); forvar973 = (forvar973 + (1'h1)))
            begin
              reg974 <= ((!($unsigned($signed((8'hb6))) ?
                      {(reg942 ? (8'ha2) : reg934),
                          $unsigned(wire929)} : (~&{reg961}))) ?
                  ($signed(((reg941 & reg910) ~^ $signed(reg948))) ?
                      (-forvar939) : reg927) : reg964);
              reg975 <= wire906;
            end
          if ($signed((&$signed($signed(reg948)))))
            begin
              reg976 <= ($signed((&reg967)) ?
                  (&$signed(reg941[(2'h2):(1'h0)])) : reg955);
              reg977 <= $signed(forvar930);
              reg978 = reg921[(1'h1):(1'h0)];
              reg979 <= $signed(($signed(($unsigned(reg950) ?
                      (reg978 && forvar969) : $signed(reg940))) ?
                  $signed((~^reg953[(4'he):(3'h4)])) : $signed(reg960)));
              reg980 = reg951;
            end
          else
            begin
              reg978 = ((7'h41) ?
                  (reg942 ?
                      ({((8'ha7) ? reg940 : (8'ha4)),
                          (+forvar973)} * ((&reg950) ?
                          $unsigned(reg945) : ((7'h45) ?
                              (8'hba) : forvar953))) : $signed(reg912)) : (~&$signed($unsigned(forvar956[(4'hd):(3'h7)]))));
              reg980 = wire902[(2'h2):(2'h2)];
              reg981 <= $unsigned($unsigned(reg918[(2'h2):(2'h2)]));
              reg982 = (((((&reg965) >>> {reg981,
                      (8'hac)}) || {((8'hab) != reg915)}) && ({{wire905,
                          (8'hbe)},
                      $signed((8'haf))} >>> (8'h9c))) ?
                  (reg942 ?
                      reg932 : (reg924[(5'h12):(5'h12)] ~^ ({reg981, reg952} ?
                          (~&reg937) : reg940[(3'h6):(1'h0)]))) : (((~&$signed(reg972)) ?
                          $unsigned((reg967 ?
                              reg960 : wire904)) : reg927[(1'h0):(1'h0)]) ?
                      reg912[(4'hd):(2'h2)] : (!({reg938, (7'h48)} ?
                          reg967 : (reg911 ? reg965 : reg930)))));
            end
          for (forvar983 = (1'h0); (forvar983 < (2'h2)); forvar983 = (forvar983 + (1'h1)))
            begin
              reg984 <= reg943[(4'h8):(3'h4)];
            end
          reg985 = $signed(($signed((reg914 & (reg980 ?
              reg918 : wire904))) < $unsigned((~&(reg942 ?
              (8'h9f) : reg936)))));
        end
    end
  assign wire986 = $unsigned(({$unsigned(reg956[(2'h2):(1'h0)]),
                           reg933[(2'h3):(2'h3)]} ?
                       $signed((((8'ha6) ?
                           reg932 : (8'hae)) & wire929[(4'h9):(3'h6)])) : reg914[(4'ha):(3'h6)]));
  always
    @(posedge clk) begin
      if ((&reg911[(5'h12):(2'h2)]))
        begin
          for (forvar987 = (1'h0); (forvar987 < (3'h4)); forvar987 = (forvar987 + (1'h1)))
            begin
              reg988 <= reg949[(4'h8):(1'h1)];
              reg989 <= $signed(wire902[(1'h1):(1'h1)]);
              reg990 = {$unsigned((reg936 >> (8'hb5)))};
            end
          for (forvar991 = (1'h0); (forvar991 < (1'h0)); forvar991 = (forvar991 + (1'h1)))
            begin
              reg992 <= (8'hb9);
            end
          for (forvar993 = (1'h0); (forvar993 < (3'h4)); forvar993 = (forvar993 + (1'h1)))
            begin
              reg994 <= {(((~^(reg961 ? reg947 : reg963)) + {reg976}) ?
                      (reg933 ?
                          ($signed(reg950) ?
                              $unsigned(reg988) : (reg977 != reg968)) : $unsigned($signed(reg967))) : ($signed((reg936 ?
                              reg936 : wire902)) ?
                          ($signed((8'h9d)) ?
                              {reg952} : $unsigned(reg922)) : reg956[(5'h12):(3'h5)])),
                  reg992};
            end
          for (forvar995 = (1'h0); (forvar995 < (1'h1)); forvar995 = (forvar995 + (1'h1)))
            begin
              reg996 = $signed((({(~|reg965)} ~^ (-(^reg926))) ?
                  ({reg961[(5'h14):(4'hf)]} ^~ reg914[(4'h8):(2'h2)]) : $signed(($unsigned(reg948) <= (reg915 ?
                      (8'hb6) : (8'hbf))))));
              reg997 <= wire906[(1'h0):(1'h0)];
              reg998 <= {(^~reg950[(1'h1):(1'h1)]),
                  (-$unsigned((~&(reg971 == reg976))))};
              reg999 = reg962[(3'h4):(1'h1)];
              reg1000 = {$unsigned(wire904[(4'hc):(4'hb)])};
            end
        end
      else
        begin
          reg987 = {(!($signed((reg947 - reg999)) <<< (&wire929[(4'h8):(3'h7)])))};
          reg988 <= ($unsigned($unsigned((reg979 - (~&reg949)))) ?
              (reg922 + (&forvar987)) : {{{$signed(reg932),
                          reg932[(1'h0):(1'h0)]},
                      reg921[(2'h2):(1'h0)]},
                  $signed(reg924[(4'he):(3'h4)])});
          if (((wire905 ?
                  $unsigned($unsigned($signed(forvar991))) : {$unsigned(reg950)}) ?
              $signed((reg912[(2'h3):(1'h0)] + $unsigned(reg987[(5'h13):(4'hf)]))) : $unsigned(reg930[(2'h3):(2'h2)])))
            begin
              reg990 = $unsigned({(reg914[(3'h4):(1'h0)] ?
                      reg971[(4'h9):(3'h6)] : $unsigned((!wire986)))});
              reg991 = wire906;
            end
          else
            begin
              reg990 = ($unsigned((reg955[(4'hb):(1'h1)] && $signed($unsigned(reg988)))) ^ ($unsigned(((reg926 << reg945) & (reg961 ?
                  wire986 : reg947))) >>> $unsigned(((reg927 >= reg930) ?
                  reg918[(4'h8):(2'h2)] : forvar995[(2'h2):(2'h2)]))));
            end
          for (forvar992 = (1'h0); (forvar992 < (1'h0)); forvar992 = (forvar992 + (1'h1)))
            begin
              reg993 = $unsigned((reg956[(3'h6):(3'h6)] ?
                  ($signed((~&(8'hae))) ?
                      $signed((|reg999)) : forvar992[(3'h6):(3'h6)]) : ({forvar991} ?
                      $signed((&reg947)) : (wire929[(1'h0):(1'h0)] ^ ((8'hb9) ?
                          reg998 : reg963)))));
              reg995 = (7'h43);
              reg996 = ((wire905[(5'h14):(4'h9)] >> $unsigned($unsigned($signed((8'ha3))))) < $unsigned({$unsigned((8'hb3))}));
              reg999 = {(|($signed(reg911[(4'h9):(1'h1)]) ?
                      reg915 : ((reg963 + reg926) ^ (reg945 + reg988)))),
                  (($signed({reg960}) ?
                          wire929[(3'h4):(1'h1)] : $signed($signed(wire929))) ?
                      $signed(reg989) : (8'haa))};
              reg1000 = (!$unsigned({wire903[(4'h9):(3'h7)]}));
            end
        end
      for (forvar1001 = (1'h0); (forvar1001 < (1'h1)); forvar1001 = (forvar1001 + (1'h1)))
        begin
          reg1002 <= $signed($signed($unsigned($unsigned(reg991[(1'h0):(1'h0)]))));
          for (forvar1003 = (1'h0); (forvar1003 < (2'h2)); forvar1003 = (forvar1003 + (1'h1)))
            begin
              reg1004 = reg968;
            end
          reg1005 <= $unsigned(($signed($unsigned((reg994 ?
              reg987 : reg922))) << $signed(($signed(reg957) ?
              reg927[(2'h2):(1'h1)] : reg967))));
          if ($signed((+$unsigned((7'h43)))))
            begin
              reg1006 = ((^~($signed(reg933[(3'h6):(2'h3)]) ?
                      (reg974[(4'h9):(1'h1)] << {(8'had)}) : {$signed(reg971)})) ?
                  $signed((8'ha4)) : (forvar992 | $unsigned($signed(reg922))));
              reg1007 = $unsigned((~{($unsigned(reg922) * $unsigned(reg922))}));
              reg1008 <= {reg948[(2'h3):(2'h3)]};
              reg1009 <= {$unsigned((($unsigned((8'had)) < (~reg945)) > {(^~reg999),
                      (wire903 >>> (8'hbd))})),
                  (reg999[(1'h0):(1'h0)] || $unsigned(((+reg996) ?
                      (~reg947) : (forvar995 ^ (8'hb3)))))};
              reg1010 = reg994;
            end
          else
            begin
              reg1008 <= reg974[(3'h5):(2'h3)];
              reg1009 <= (reg948[(2'h3):(2'h3)] <<< ($signed(reg926) <= reg1005[(3'h6):(3'h4)]));
              reg1011 <= reg996[(1'h1):(1'h0)];
              reg1012 = ((reg950 || ({$unsigned(reg936)} ?
                  reg1007[(3'h7):(1'h0)] : {reg993})) != (~^$unsigned(({wire905,
                  reg931} <<< (reg984 ? reg960 : reg935)))));
              reg1013 <= ((({(+reg965)} <<< reg999[(1'h0):(1'h0)]) ?
                      (($signed((8'hbe)) >= (reg997 ? reg910 : reg1008)) ?
                          ($unsigned((7'h47)) ?
                              $unsigned(reg926) : (reg979 ?
                                  reg1010 : reg922)) : (^(reg998 ?
                              reg1008 : reg911))) : $signed(reg967)) ?
                  $signed((7'h44)) : {forvar992[(4'hd):(1'h1)],
                      $signed(wire906[(2'h2):(1'h1)])});
            end
          reg1014 <= reg990[(2'h3):(1'h0)];
        end
      if ((+$unsigned($signed((8'hab)))))
        begin
          if ($signed($signed(({reg933[(3'h4):(1'h1)], (8'hba)} ?
              $unsigned((reg977 || (8'hbb))) : reg927))))
            begin
              reg1015 = $unsigned((-($signed(wire906) <= reg1008)));
              reg1016 <= $signed(reg999[(4'h9):(2'h2)]);
              reg1017 <= wire902;
              reg1018 <= $signed(($signed((((8'ha5) * reg922) > (reg993 | reg993))) << (-(&(-forvar992)))));
              reg1019 = (|(($unsigned(reg975) ? forvar987 : (8'h9c)) ?
                  (8'h9c) : $signed($signed($signed((8'hac))))));
            end
          else
            begin
              reg1016 <= $signed($signed({(!(reg989 ? reg1017 : forvar1001)),
                  reg1008[(3'h4):(2'h2)]}));
              reg1019 = $signed($unsigned(forvar995));
            end
        end
      else
        begin
          reg1016 <= (^$signed(reg1010[(1'h0):(1'h0)]));
          if ({reg926[(1'h1):(1'h0)]})
            begin
              reg1019 = $unsigned((8'h9f));
              reg1020 <= (7'h42);
              reg1021 = $unsigned($unsigned((&$unsigned((reg1010 >= reg931)))));
              reg1022 <= reg930;
            end
          else
            begin
              reg1019 = ({reg952[(5'h10):(4'hd)]} << (~&{$unsigned((~reg977))}));
              reg1020 <= ($unsigned(((7'h47) ~^ $signed(wire903[(4'ha):(2'h2)]))) ?
                  (^$unsigned($signed((forvar987 ?
                      reg968 : forvar992)))) : $unsigned(($unsigned((8'h9c)) - reg912)));
              reg1022 <= ((~^(((-reg992) ?
                      (forvar995 ?
                          (8'h9e) : reg996) : $signed(reg1012)) ^ wire929[(3'h4):(2'h3)])) ?
                  (^~reg941) : forvar993[(1'h1):(1'h0)]);
              reg1023 = $unsigned((-$unsigned((((8'hbf) & reg979) >> reg990))));
              reg1024 <= $signed($signed((reg1002[(4'h9):(2'h3)] < reg1014)));
            end
          reg1025 = ((-$signed((reg941 != reg1023))) + (~|(8'hb8)));
        end
    end
  always
    @(posedge clk) begin
      if ($signed(reg931[(2'h3):(1'h1)]))
        begin
          reg1026 = (($signed($signed(((7'h45) == reg1008))) ?
                  reg997 : (&({reg949, (8'hb3)} == {(7'h45)}))) ?
              ({(reg935[(4'hb):(1'h1)] ?
                      (reg971 <= reg926) : reg948[(3'h4):(1'h1)]),
                  {(reg1011 || reg914)}} | $signed($signed(reg1016))) : reg1024[(3'h6):(3'h6)]);
        end
      else
        begin
          for (forvar1026 = (1'h0); (forvar1026 < (1'h1)); forvar1026 = (forvar1026 + (1'h1)))
            begin
              reg1027 <= reg960;
            end
          reg1028 <= reg961[(4'h9):(2'h3)];
          if ($signed(($unsigned(((reg921 ? (7'h44) : reg915) ?
                  reg941 : reg912[(5'h14):(4'h9)])) ?
              reg912[(3'h4):(2'h2)] : reg979[(3'h7):(3'h5)])))
            begin
              reg1029 = {(reg933[(3'h6):(2'h3)] | $unsigned((~^(reg956 ?
                      reg968 : reg933))))};
              reg1030 <= ($unsigned($unsigned((|(~|reg988)))) <= reg1020[(4'h8):(3'h5)]);
              reg1031 <= $signed((reg998 ?
                  (reg968[(2'h2):(1'h0)] ^~ {$signed(reg961),
                      reg984[(3'h6):(1'h0)]}) : (-$unsigned($unsigned(reg1020)))));
              reg1032 = ($unsigned(((reg1022 ?
                          reg1020[(3'h7):(2'h2)] : $unsigned(reg1029)) ?
                      (~&$unsigned(reg1014)) : ($unsigned(reg981) ?
                          (-reg1026) : (!reg931)))) ?
                  reg931[(4'hd):(4'ha)] : reg931[(3'h7):(1'h0)]);
              reg1033 <= wire906[(1'h1):(1'h1)];
            end
          else
            begin
              reg1030 <= $signed(reg1009[(3'h4):(1'h0)]);
              reg1032 = reg1017;
            end
          reg1034 = ((((-reg924[(2'h3):(1'h0)]) >= (-(reg998 & reg977))) < $signed((reg967[(3'h5):(2'h2)] ?
                  $signed(reg968) : reg926[(4'h8):(2'h2)]))) ?
              $signed((-$signed((|wire903)))) : (-$signed({(reg911 * (8'ha0))})));
        end
      for (forvar1035 = (1'h0); (forvar1035 < (3'h4)); forvar1035 = (forvar1035 + (1'h1)))
        begin
          reg1036 <= {($signed($signed($signed(reg976))) < ((8'hae) != $signed(wire986)))};
          reg1037 = $signed(((reg1005 ?
              (~^reg984[(3'h4):(1'h0)]) : reg956) ^~ (!(|reg1034[(4'hc):(4'h8)]))));
          for (forvar1038 = (1'h0); (forvar1038 < (2'h3)); forvar1038 = (forvar1038 + (1'h1)))
            begin
              reg1039 <= (8'ha3);
            end
          if ({reg981[(3'h5):(2'h2)]})
            begin
              reg1040 <= (^reg1032[(2'h3):(1'h0)]);
              reg1041 <= $signed(reg971[(3'h7):(3'h4)]);
              reg1042 = $signed($signed($signed((&wire929[(2'h2):(2'h2)]))));
            end
          else
            begin
              reg1040 <= reg1013[(4'hc):(4'ha)];
              reg1041 <= $signed({$signed((7'h48))});
              reg1042 = (((reg1005 ?
                  $unsigned((&reg1013)) : $unsigned((|reg1024))) - ((^reg1037[(1'h0):(1'h0)]) ?
                  wire903 : $signed((reg1037 ?
                      reg916 : reg949)))) || forvar1038[(3'h6):(2'h2)]);
            end
        end
      for (forvar1043 = (1'h0); (forvar1043 < (2'h2)); forvar1043 = (forvar1043 + (1'h1)))
        begin
          reg1044 <= ((|($signed($unsigned(reg962)) ?
              $unsigned((~&reg916)) : ($unsigned(wire904) ?
                  (reg1029 > reg956) : reg989[(1'h0):(1'h0)]))) ^~ ((~^{$unsigned(reg960)}) ?
              (~|(~&$unsigned((7'h40)))) : reg1032[(4'hb):(4'h8)]));
          if ((((reg1016[(2'h2):(2'h2)] ?
              {(reg1011 ? (8'had) : reg1030), $signed(reg1022)} : ((~^reg1026) ?
                  (reg1033 ^ reg916) : $signed(reg1029))) >> (~&((reg957 ?
              reg945 : reg1014) * {reg932}))) & $unsigned({((~|reg1034) >> reg992[(3'h7):(3'h4)])})))
            begin
              reg1045 <= (8'hb5);
              reg1046 = $signed($unsigned(reg927[(1'h0):(1'h0)]));
              reg1047 <= reg975;
            end
          else
            begin
              reg1046 = ({{((reg924 <= (8'hb1)) < $signed((8'h9f)))},
                  $signed({(reg994 || reg950),
                      wire903[(2'h3):(1'h1)]})} * (reg960 - $unsigned(($unsigned(reg936) ?
                  reg912[(4'h9):(2'h2)] : {reg955}))));
              reg1048 = (^($signed(((reg974 ?
                      (8'had) : reg918) ^ ((8'hae) > (7'h42)))) ?
                  ({$signed(reg979), (~reg998)} ?
                      ($signed(reg976) <<< $signed(wire929)) : reg910) : $signed(((^reg918) & {reg1018,
                      reg1029}))));
              reg1049 = {(reg924[(5'h12):(4'hb)] ?
                      {(reg952 ? $unsigned(reg1013) : reg1047[(3'h7):(1'h1)]),
                          reg1026} : ($unsigned($signed(reg994)) ?
                          {(reg965 >= (8'h9f)),
                              reg935[(2'h2):(2'h2)]} : ((8'hbc) ?
                              ((8'hb7) <= reg1002) : (&reg924)))),
                  ((($signed(reg967) < reg1031[(1'h0):(1'h0)]) ?
                      reg1008[(5'h13):(3'h5)] : $unsigned($signed(reg1002))) & (|$signed(reg977[(4'h8):(3'h5)])))};
              reg1050 <= $signed($signed(reg1022[(4'h8):(4'h8)]));
            end
          if (({$unsigned((+(|reg916)))} == reg912))
            begin
              reg1051 = ($signed((^~$unsigned($unsigned(wire929)))) || $unsigned((-((reg962 ?
                  (8'ha1) : reg1036) * (-reg977)))));
              reg1052 = $signed($signed(($unsigned(reg949[(4'h9):(2'h3)]) ?
                  wire903[(4'h8):(3'h4)] : ($signed((8'hb2)) - (reg1028 ^~ reg1018)))));
              reg1053 <= ($unsigned(reg1040[(3'h4):(2'h2)]) ?
                  {((-reg971) >= reg955)} : wire902);
            end
          else
            begin
              reg1051 = reg1036[(1'h1):(1'h1)];
              reg1052 = ($signed((8'hbc)) ?
                  ((~&($signed(reg997) ?
                      (^reg912) : reg1041[(4'hd):(4'ha)])) <<< (~&((~&reg998) ?
                      (wire986 || (8'h9d)) : (reg1008 | reg977)))) : (^~(forvar1035 ?
                      $unsigned((reg912 >> reg1052)) : ((^~reg1041) ?
                          $unsigned(reg994) : $signed(reg1037)))));
              reg1053 <= $unsigned(reg997);
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned($signed($signed(((reg1017 ? reg977 : reg1036) | (8'hb3))))))
        begin
          reg1054 <= reg1040;
          reg1055 = (^~{$signed($unsigned((8'hb9)))});
          for (forvar1056 = (1'h0); (forvar1056 < (1'h0)); forvar1056 = (forvar1056 + (1'h1)))
            begin
              reg1057 <= {((($unsigned(reg1011) && {reg1024}) + reg976) | reg998),
                  reg932[(2'h3):(1'h0)]};
              reg1058 <= (((wire906[(2'h3):(1'h0)] ?
                          (~&(7'h44)) : $signed(reg930[(1'h1):(1'h0)])) ?
                      reg968[(1'h1):(1'h1)] : reg1047[(4'ha):(1'h0)]) ?
                  $unsigned($unsigned(reg933[(1'h0):(1'h0)])) : (&(reg955[(4'h9):(3'h7)] | $signed({reg911}))));
              reg1059 <= $signed((reg941 & {$unsigned((~^wire904))}));
              reg1060 = reg1058;
              reg1061 <= (~|(~&(|$unsigned(((7'h45) ? (7'h42) : reg935)))));
            end
          reg1062 = (&{{$unsigned(((8'ha0) ? reg1017 : reg947))}});
          for (forvar1063 = (1'h0); (forvar1063 < (1'h0)); forvar1063 = (forvar1063 + (1'h1)))
            begin
              reg1064 <= wire903[(1'h1):(1'h0)];
              reg1065 <= ($signed(wire903) ?
                  (reg971 ?
                      reg933 : (~&($unsigned((8'hb4)) ?
                          (reg1017 ?
                              reg1016 : reg998) : reg1040))) : (reg1060[(5'h11):(4'ha)] ?
                      ($unsigned((reg1054 ^~ (8'ha3))) ?
                          $signed((7'h46)) : $unsigned((reg965 + reg916))) : reg1060));
              reg1066 = reg984[(3'h5):(1'h0)];
            end
        end
      else
        begin
          reg1054 <= {((((reg988 ? (8'hb6) : reg1013) ?
                          $signed(reg945) : (!reg992)) ?
                      (^(&reg961)) : (reg975[(1'h1):(1'h0)] & {reg1064})) ?
                  (reg933 >> (|reg1031)) : $signed((~|(reg1014 == reg952)))),
              (((reg1005 ^~ $unsigned((7'h43))) ?
                  reg1005 : ($signed(reg1064) ?
                      ((8'hb8) ?
                          reg979 : reg1033) : reg1009[(3'h5):(1'h0)])) == $signed((|(&wire902))))};
          if (reg960)
            begin
              reg1055 = {$signed(reg998[(3'h6):(3'h4)]),
                  forvar1056[(3'h7):(3'h5)]};
              reg1056 <= (~|(~$signed(reg975)));
              reg1060 = {(reg1053[(2'h3):(2'h2)] * $unsigned(((reg926 ?
                          reg1044 : wire929) ?
                      reg1040 : (reg1030 ? reg1064 : reg968)))),
                  {(wire902 ? (+(reg922 & reg931)) : {(+reg1062)})}};
              reg1061 <= ($signed($unsigned($signed(reg956[(3'h7):(3'h4)]))) * (~&$signed((^(reg1055 ?
                  reg930 : reg1016)))));
              reg1063 <= ((~&(-{reg979[(2'h3):(2'h2)]})) ?
                  (~|reg962[(2'h3):(2'h3)]) : (-((&(reg1054 ?
                          (8'ha1) : reg1017)) ?
                      (~|reg1027) : ($unsigned(wire986) ?
                          (reg1009 != (8'ha4)) : (^reg926)))));
            end
          else
            begin
              reg1056 <= {$unsigned($unsigned(((reg977 >> forvar1063) ?
                      $unsigned(reg936) : {reg952, reg1062})))};
              reg1057 <= $unsigned(reg1057);
              reg1060 = reg1053;
              reg1062 = (!((8'hac) >>> (reg927 <= $signed((wire929 * reg916)))));
            end
          reg1064 <= {(~|(reg976[(3'h7):(3'h5)] | $unsigned({reg960})))};
          for (forvar1065 = (1'h0); (forvar1065 < (3'h4)); forvar1065 = (forvar1065 + (1'h1)))
            begin
              reg1066 = reg950[(1'h1):(1'h0)];
              reg1067 = (^~$signed(reg1002));
            end
          if (reg989[(2'h2):(1'h0)])
            begin
              reg1068 = $unsigned(((((~|reg960) & $unsigned(reg936)) >= $unsigned(reg976[(4'h9):(3'h6)])) ?
                  (reg1020 == (8'hb9)) : $signed(((reg1056 | reg948) ?
                      (reg988 ? (8'ha0) : reg916) : $signed(reg981)))));
              reg1069 <= ($signed((|(~^(reg965 ^~ reg1020)))) ?
                  ((((reg1005 != (7'h48)) >= $signed(forvar1065)) <<< $signed($signed(reg968))) ?
                      (!reg968) : (~|(!(~(7'h47))))) : $signed(reg956));
            end
          else
            begin
              reg1068 = {$unsigned($unsigned(($signed(reg1055) * (reg927 ?
                      reg1045 : reg956))))};
              reg1070 = reg1054[(3'h7):(3'h4)];
              reg1071 <= ($signed($signed((~&(reg1028 << reg1016)))) ?
                  reg1033 : (+($unsigned((reg1068 ? reg1069 : reg971)) ?
                      $unsigned(reg1030[(3'h5):(2'h2)]) : ((reg952 ?
                          reg992 : reg962) + (reg915 ? reg1063 : reg1059)))));
            end
        end
      if (reg1028)
        begin
          for (forvar1072 = (1'h0); (forvar1072 < (2'h2)); forvar1072 = (forvar1072 + (1'h1)))
            begin
              reg1073 <= (~|reg1036[(3'h6):(2'h3)]);
              reg1074 = $signed((reg918[(3'h5):(1'h1)] ?
                  wire902 : (((^~reg997) <= (wire905 ?
                      reg976 : (7'h45))) == (!(|wire929)))));
              reg1075 <= (8'ha8);
              reg1076 = $unsigned($unsigned(reg955));
            end
          if ((~($signed(({(8'ha6), reg1063} & reg918[(1'h0):(1'h0)])) ?
              reg948[(3'h4):(1'h0)] : reg979)))
            begin
              reg1077 = ((8'hbc) ?
                  (~^$signed($unsigned((reg1008 + (8'hb6))))) : ((^~(8'hba)) << (({reg1017,
                          reg1067} ?
                      $unsigned(reg1063) : {reg1009}) <= reg988[(2'h3):(1'h1)])));
              reg1078 = reg974;
              reg1079 <= {(|reg949[(4'h9):(4'h9)]),
                  (($signed((^~reg947)) ?
                      (~(reg952 ? reg927 : reg931)) : ((reg930 ?
                              reg960 : reg1011) ?
                          $signed(reg968) : ((8'h9d) ?
                              reg933 : (8'hbe)))) == (reg1071[(3'h5):(3'h4)] ?
                      {(reg912 ^~ reg1005)} : (^~((8'hbd) ?
                          reg1024 : wire904))))};
            end
          else
            begin
              reg1077 = $signed(reg916[(5'h13):(1'h0)]);
              reg1078 = reg967[(2'h3):(2'h3)];
              reg1079 <= reg924[(4'h8):(1'h0)];
            end
          reg1080 <= ((|(reg1075[(4'h8):(1'h1)] ?
              reg1064 : ($signed(reg941) ?
                  (reg910 ~^ reg988) : {reg1074}))) <= (($unsigned(reg1022[(4'hf):(2'h2)]) < ((!reg1040) ?
              reg1078[(4'h9):(2'h3)] : ((7'h46) & reg962))) > $unsigned($unsigned((reg965 ?
              reg930 : reg1058)))));
          for (forvar1081 = (1'h0); (forvar1081 < (3'h4)); forvar1081 = (forvar1081 + (1'h1)))
            begin
              reg1082 = (wire906[(4'h9):(3'h7)] ?
                  (|reg1075[(2'h2):(2'h2)]) : (8'hb1));
              reg1083 = reg962;
              reg1084 = {((^~reg955[(1'h1):(1'h0)]) - (($unsigned(reg918) != reg984) << (reg914[(3'h5):(3'h5)] ^ {(8'hb0)})))};
              reg1085 = reg933[(2'h2):(2'h2)];
              reg1086 = {$signed($signed(({reg975} ?
                      $unsigned(reg965) : ((8'hbf) ? reg1030 : forvar1081)))),
                  reg1078[(2'h3):(2'h2)]};
            end
          if (((reg981 != $signed(((reg1059 ? reg950 : (8'h9e)) ?
              {(8'h9f)} : $unsigned(reg1027)))) > $signed((reg1066 & reg968[(2'h2):(1'h0)]))))
            begin
              reg1087 <= reg1078;
              reg1088 = (forvar1063[(4'hd):(3'h4)] || $signed((^({reg1058} >= reg922[(3'h6):(1'h1)]))));
              reg1089 = $signed((reg926[(4'hd):(4'h9)] ?
                  {($unsigned(reg1075) ^ reg955[(1'h0):(1'h0)])} : {$signed((~&reg1016))}));
            end
          else
            begin
              reg1087 <= (~$signed((^~$unsigned(((8'ha6) ~^ (8'ha5))))));
              reg1090 <= ((!(~|reg988[(3'h6):(2'h3)])) >> reg1070[(3'h5):(2'h3)]);
            end
        end
      else
        begin
          if ($signed(((-$unsigned(reg922[(2'h3):(2'h3)])) ?
              {$signed((wire929 && reg1064)),
                  $signed((+reg1076))} : ($unsigned((!reg1040)) != (reg1030 ?
                  $unsigned(reg1055) : (!reg979))))))
            begin
              reg1072 = reg947[(1'h0):(1'h0)];
              reg1073 <= $unsigned(reg1031);
              reg1075 <= ({reg957} > reg1039);
            end
          else
            begin
              reg1073 <= {$unsigned((reg962[(1'h0):(1'h0)] > ((~|wire929) < $unsigned(reg955))))};
              reg1074 = (&$unsigned(reg975[(1'h0):(1'h0)]));
              reg1076 = (~&$signed(reg1069));
              reg1077 = $unsigned((~&{$signed((&reg911))}));
            end
          reg1078 = ({$unsigned(reg1068),
              reg998[(1'h1):(1'h0)]} ^~ (^(~&$signed((reg1028 >= reg1072)))));
          reg1081 = reg916[(1'h0):(1'h0)];
        end
      for (forvar1091 = (1'h0); (forvar1091 < (3'h4)); forvar1091 = (forvar1091 + (1'h1)))
        begin
          reg1092 = reg1002;
          if (reg1073)
            begin
              reg1093 <= (^~($unsigned($signed(reg956[(2'h2):(1'h0)])) || ($signed((~^reg941)) ^ (reg927[(2'h2):(1'h1)] ?
                  ((8'hbc) && reg962) : (^(8'hb3))))));
              reg1094 <= {{$signed(reg1040[(4'he):(4'h9)])}};
            end
          else
            begin
              reg1095 = ($signed($signed(reg955[(3'h4):(1'h0)])) ?
                  $signed((reg994 & (reg949 >>> (!(8'ha8))))) : $unsigned($unsigned((reg1060[(5'h12):(4'hd)] >> (&reg1055)))));
              reg1096 <= reg1061;
              reg1097 <= $unsigned(($unsigned((~&$unsigned(reg924))) ?
                  wire906[(4'h9):(4'h8)] : reg994[(4'hd):(3'h7)]));
              reg1098 = $signed(reg1058);
              reg1099 <= (~^$signed(reg947));
            end
        end
    end
  assign wire1100 = ($signed($signed((reg1058[(3'h7):(3'h6)] ?
                            wire906[(2'h2):(1'h0)] : (reg1030 >>> reg1014)))) ?
                        ($signed(({reg979} != (!(7'h47)))) ?
                            (({reg924, reg1071} <= reg1030) ?
                                reg932[(2'h3):(2'h2)] : (|reg981[(3'h4):(1'h0)])) : ($unsigned($unsigned(reg967)) ?
                                ($unsigned((8'ha6)) ?
                                    (reg960 ^~ wire986) : (reg933 ?
                                        reg914 : reg945)) : (8'ha1))) : (((8'haf) ^ reg927) * (reg1097[(3'h5):(3'h4)] ?
                            ($signed(reg1069) <= (reg1065 ?
                                (8'hb0) : reg998)) : $unsigned($signed(reg965)))));
  assign wire1101 = (8'h9c);
  assign wire1102 = (~($unsigned($signed((wire902 > reg933))) ?
                        $unsigned(((~^reg984) ?
                            (reg956 != wire1100) : $signed(reg1005))) : ($unsigned((&reg998)) >= reg1087)));
  assign wire1103 = reg981[(1'h1):(1'h0)];
  assign wire1104 = reg971;
  always
    @(posedge clk) begin
      if (({reg988} < (^~(reg1028 ? (8'h9d) : $signed($unsigned(reg974))))))
        begin
          reg1105 <= ($signed((($signed(reg1013) ~^ (reg1087 & reg914)) ?
              $unsigned({reg988,
                  reg1030}) : $unsigned((reg1097 >= reg971)))) - ({reg1065[(4'hb):(3'h5)]} ?
              {reg1033,
                  ($unsigned(reg998) ~^ ((8'ha2) ~^ reg1041))} : reg945[(3'h6):(3'h6)]));
          reg1106 = (~reg963[(4'hd):(2'h2)]);
        end
      else
        begin
          reg1106 = $unsigned(reg921[(1'h0):(1'h0)]);
          for (forvar1107 = (1'h0); (forvar1107 < (2'h2)); forvar1107 = (forvar1107 + (1'h1)))
            begin
              reg1108 = (~&$signed(reg930[(1'h1):(1'h0)]));
              reg1109 <= $signed(reg927);
              reg1110 = $signed({$signed(($signed(reg962) ?
                      $unsigned(reg1079) : $signed(wire1100))),
                  reg1071[(3'h4):(1'h0)]});
              reg1111 <= (&($unsigned((reg1056[(2'h3):(1'h0)] < $unsigned(wire903))) ?
                  (8'h9d) : (8'hbf)));
            end
          reg1112 = wire905;
          if ((^~reg1073[(4'hb):(2'h2)]))
            begin
              reg1113 <= $signed(reg1073[(5'h11):(3'h5)]);
              reg1114 = (&reg1008[(4'h9):(4'h9)]);
            end
          else
            begin
              reg1113 <= {((-(^~reg992)) ?
                      $unsigned({reg926, reg1014}) : reg956[(4'he):(4'h9)]),
                  (~reg948[(2'h2):(2'h2)])};
            end
        end
      for (forvar1115 = (1'h0); (forvar1115 < (3'h4)); forvar1115 = (forvar1115 + (1'h1)))
        begin
          reg1116 <= reg1069;
          reg1117 = reg1041[(4'hd):(4'hc)];
          if (reg1071)
            begin
              reg1118 = $unsigned((&reg1013[(2'h2):(1'h0)]));
            end
          else
            begin
              reg1119 <= $unsigned($signed(reg1053));
              reg1120 = ((($signed((reg960 ?
                      wire1104 : reg1053)) >>> reg1105) == (!$signed((reg1045 ?
                      wire1101 : forvar1115)))) ?
                  $signed($unsigned((-$unsigned(reg1016)))) : reg1045[(3'h4):(2'h2)]);
              reg1121 = $signed(wire1101[(1'h1):(1'h0)]);
              reg1122 <= reg1039;
            end
          if (((8'h9e) * (8'h9e)))
            begin
              reg1123 = (~|reg1120);
              reg1124 <= reg1118[(2'h3):(2'h3)];
            end
          else
            begin
              reg1124 <= {$unsigned($signed(($signed(reg1058) > reg1028)))};
            end
          if (((~($unsigned({reg998}) != (7'h46))) <= reg998))
            begin
              reg1125 = $unsigned({((^{reg965}) != $signed($signed(reg1094)))});
              reg1126 = reg974;
              reg1127 = reg1075[(1'h0):(1'h0)];
              reg1128 = reg968[(1'h0):(1'h0)];
            end
          else
            begin
              reg1129 <= {(&($unsigned($signed(reg910)) ?
                      reg1039 : (~^reg1013[(3'h4):(3'h4)]))),
                  (-reg1039[(2'h2):(1'h1)])};
              reg1130 <= (7'h42);
            end
        end
      if ($signed($signed((~&reg1061))))
        begin
          reg1131 = $unsigned(reg1108[(4'hd):(1'h0)]);
          if (reg1036[(2'h3):(1'h1)])
            begin
              reg1132 <= reg1128[(2'h2):(1'h1)];
              reg1133 <= reg1036[(3'h4):(2'h2)];
              reg1134 = reg952[(4'h8):(2'h3)];
              reg1135 = $unsigned($signed({reg949,
                  (reg1105 ? reg1030[(3'h6):(3'h5)] : (wire1103 < (7'h43)))}));
            end
          else
            begin
              reg1134 = ($signed(reg1016) ^ reg924);
              reg1136 <= (^$signed(reg976[(1'h1):(1'h1)]));
              reg1137 <= $unsigned(reg1125);
              reg1138 = reg1099;
              reg1139 <= reg1133;
            end
          reg1140 = wire905;
          reg1141 <= $unsigned((^~reg1053[(4'hc):(2'h3)]));
        end
      else
        begin
          for (forvar1131 = (1'h0); (forvar1131 < (1'h0)); forvar1131 = (forvar1131 + (1'h1)))
            begin
              reg1132 <= (((wire1103[(1'h1):(1'h0)] - $unsigned($unsigned(wire904))) >>> (^~(^(+reg1047)))) > ($signed((8'hb7)) ?
                  ($unsigned((!reg961)) == reg927[(1'h0):(1'h0)]) : (reg1127[(1'h0):(1'h0)] < reg971[(4'hd):(1'h0)])));
              reg1133 <= wire904[(4'hc):(2'h3)];
            end
          for (forvar1134 = (1'h0); (forvar1134 < (1'h0)); forvar1134 = (forvar1134 + (1'h1)))
            begin
              reg1135 = $unsigned($signed((forvar1107 ?
                  reg1022[(5'h10):(4'hb)] : reg1093)));
              reg1136 <= {forvar1134[(5'h18):(1'h1)]};
              reg1137 <= $signed((~|(&(reg1121 ?
                  $signed((8'ha5)) : (~reg1031)))));
              reg1139 <= $unsigned((($unsigned(reg1024[(4'hd):(4'hd)]) ~^ reg1093) >> (($unsigned(reg1059) ?
                      (reg1124 ? reg971 : reg1063) : (reg914 > (8'had))) ?
                  reg1123[(4'hb):(3'h5)] : $unsigned($signed(wire902)))));
              reg1141 <= ((reg1047 ?
                  $unsigned(((reg1129 ? reg967 : reg1045) ?
                      $signed(reg1045) : $unsigned(reg1045))) : {($signed(reg1127) == reg1117),
                      (~^(reg1116 == reg1008))}) != {reg1005, (7'h46)});
            end
          reg1142 = wire906;
        end
      for (forvar1143 = (1'h0); (forvar1143 < (1'h0)); forvar1143 = (forvar1143 + (1'h1)))
        begin
          reg1144 <= (reg918[(3'h4):(1'h0)] && ($signed($unsigned((~^reg1011))) ?
              $unsigned({$unsigned((8'hbc))}) : wire1101));
          for (forvar1145 = (1'h0); (forvar1145 < (1'h0)); forvar1145 = (forvar1145 + (1'h1)))
            begin
              reg1146 <= {$signed((|$signed(((7'h46) + (7'h40))))),
                  ((~^(~^(reg1069 ?
                      reg992 : reg974))) >= {$unsigned($signed((7'h41))),
                      reg1045[(4'h8):(1'h1)]})};
              reg1147 = $unsigned({wire1104[(1'h1):(1'h0)],
                  $unsigned($unsigned($unsigned(forvar1115)))});
              reg1148 = $unsigned({(&reg1094[(3'h5):(2'h2)]),
                  (reg1020[(4'h9):(1'h1)] && {((8'h9d) ^~ reg945)})});
            end
          for (forvar1149 = (1'h0); (forvar1149 < (3'h4)); forvar1149 = (forvar1149 + (1'h1)))
            begin
              reg1150 = {reg981[(2'h3):(1'h0)],
                  ($unsigned((reg1119 ? {reg1014} : (8'h9f))) ?
                      reg957 : (($unsigned(reg948) ^ $signed(reg1136)) + reg1028))};
              reg1151 <= ($signed({((reg1124 ? reg1014 : reg1013) >>> (reg1125 ?
                          reg1079 : reg1058))}) ?
                  reg989 : $signed(reg1017));
            end
          if (reg962)
            begin
              reg1152 <= (($signed({$signed((7'h42)), wire929}) ?
                      reg926 : ((reg1036 ~^ (reg1138 ? (8'haf) : reg1114)) ?
                          {reg1080[(1'h0):(1'h0)]} : (&(7'h43)))) ?
                  (reg1016 ~^ (^(~|(|reg1146)))) : (~|($signed(reg1018[(4'he):(3'h5)]) ?
                      ((^reg1016) ?
                          ((8'ha5) ?
                              forvar1107 : reg1017) : (reg988 <= reg1079)) : $unsigned(reg1135))));
            end
          else
            begin
              reg1152 <= reg1141;
            end
        end
    end
  assign wire1153 = reg997;
  always
    @(posedge clk) begin
      if ((^~(~|({reg984[(3'h4):(2'h3)]} ?
          ((reg1099 && reg989) ^ $signed(wire1101)) : reg977[(3'h7):(3'h5)]))))
        begin
          reg1154 <= (~reg1059[(5'h18):(4'h8)]);
          if ($unsigned($unsigned($signed(($unsigned(reg968) ~^ (reg1050 ?
              reg927 : reg989))))))
            begin
              reg1155 <= $unsigned($signed(reg1099[(1'h1):(1'h0)]));
              reg1156 = $unsigned($unsigned($signed((reg921[(1'h0):(1'h0)] ?
                  reg1119 : (reg918 ? reg1105 : (8'ha6))))));
              reg1157 = $unsigned($signed(wire1104));
            end
          else
            begin
              reg1156 = (&(reg1017 <<< $unsigned($signed(reg921[(1'h1):(1'h0)]))));
              reg1157 = reg1039[(2'h3):(2'h3)];
            end
          reg1158 = {{$signed((reg1156[(1'h0):(1'h0)] - {(7'h41)}))},
              $signed($signed($signed({(7'h44), reg1146})))};
          if (reg1154)
            begin
              reg1159 = reg912[(3'h4):(1'h0)];
              reg1160 = reg1031[(1'h0):(1'h0)];
              reg1161 <= $unsigned((~^$signed(($signed(reg1105) ?
                  (reg1022 ? reg1152 : reg1158) : (reg1047 ?
                      reg945 : reg1017)))));
              reg1162 = reg915[(1'h0):(1'h0)];
              reg1163 <= $unsigned(reg1022);
            end
          else
            begin
              reg1161 <= (wire1100 ?
                  $unsigned($unsigned((^~$unsigned(reg910)))) : (~reg1050));
              reg1163 <= $unsigned((reg1156[(3'h5):(1'h1)] >= reg1139[(3'h5):(3'h4)]));
              reg1164 <= (((reg1017 ?
                      $signed(reg1017) : (~$unsigned(reg1161))) ?
                  $signed(reg1157) : ((wire1101[(2'h3):(1'h1)] ?
                          (reg1018 ? reg1156 : reg931) : {reg968, (8'ha9)}) ?
                      {{reg1013, reg1073},
                          $signed(reg950)} : $unsigned((|reg915)))) >>> ((^(reg989[(1'h0):(1'h0)] ?
                  (~&reg1005) : $unsigned(reg1028))) * wire906));
              reg1165 <= reg1041[(1'h0):(1'h0)];
              reg1166 <= {reg947};
            end
        end
      else
        begin
          reg1154 <= (reg981 ?
              $signed(reg1116) : (reg968[(1'h1):(1'h1)] & ($unsigned($signed(reg965)) ?
                  reg922[(1'h0):(1'h0)] : {$signed((7'h43))})));
          if (((!{{(reg977 ? (8'hba) : reg936), (reg949 & reg955)},
                  reg977[(2'h2):(1'h0)]}) ?
              (&(($unsigned((8'hbd)) ?
                      (reg930 ? reg1113 : (8'ha4)) : reg1045[(2'h3):(2'h2)]) ?
                  $unsigned(reg1061) : $unsigned({reg992}))) : $signed($signed(reg960))))
            begin
              reg1155 <= reg1030[(1'h1):(1'h0)];
              reg1156 = reg1090[(5'h11):(4'he)];
              reg1161 <= reg1122;
              reg1163 <= reg1040[(4'hc):(2'h3)];
            end
          else
            begin
              reg1155 <= {reg981, (8'hbd)};
              reg1161 <= (~|reg949[(1'h0):(1'h0)]);
              reg1163 <= reg941;
              reg1167 = (~^($signed((^$signed((7'h48)))) ?
                  (~reg918[(4'h9):(4'h8)]) : $unsigned(((reg1087 ?
                      reg1020 : reg915) << reg952))));
              reg1168 <= reg948[(1'h0):(1'h0)];
            end
          reg1169 = ($unsigned({$signed((8'hbc)),
              (~(reg1163 ? reg911 : reg1124))}) >>> reg963);
          reg1170 <= (-$unsigned(((((8'ha5) ?
                  (8'hbd) : (7'h44)) * $unsigned(reg931)) ?
              reg955 : (((8'hb1) <= reg955) ?
                  reg1130[(1'h0):(1'h0)] : (~reg945)))));
          reg1171 = (^(!reg1141[(4'h9):(3'h5)]));
        end
      if ((reg971[(4'hc):(1'h1)] ? reg1132 : (&(+$unsigned({reg1093})))))
        begin
          reg1172 = reg997[(1'h1):(1'h0)];
          reg1173 <= reg949;
        end
      else
        begin
          reg1173 <= (-(($signed($unsigned((8'haa))) <<< $unsigned((reg1167 ?
                  reg1028 : reg1031))) ?
              $signed(($signed(wire929) & (8'h9f))) : $signed(((reg1069 ^ reg1111) <<< $unsigned(reg1028)))));
          reg1174 = wire1103[(3'h7):(3'h6)];
          reg1175 = reg988[(1'h0):(1'h0)];
        end
      reg1176 = (reg1054 ?
          ((reg1137[(1'h1):(1'h0)] != (!$signed(reg1175))) ^ ($unsigned((reg1154 - reg1061)) ?
              (|$signed(reg1159)) : (8'hb0))) : $signed((reg1122[(4'hc):(4'h8)] ?
              $signed(((8'ha0) <= (8'ha6))) : ($signed(reg926) >= reg949))));
    end
  assign wire1177 = ($signed((~reg921[(2'h2):(1'h1)])) & ($unsigned(reg997[(4'h9):(4'h8)]) ?
                        wire1103[(3'h6):(2'h3)] : (^~($unsigned(reg1053) ?
                            $unsigned(reg960) : (reg1053 >>> reg948)))));
  assign wire1178 = (-(8'had));
  assign wire1179 = reg914;
  assign wire1180 = $signed((~|((~|reg1094[(4'hd):(2'h3)]) ~^ $unsigned(reg1020[(1'h1):(1'h0)]))));
  assign wire1181 = $unsigned(reg1033[(3'h6):(3'h5)]);
  assign wire1182 = reg1005[(3'h4):(3'h4)];
  always
    @(posedge clk) begin
      for (forvar1183 = (1'h0); (forvar1183 < (1'h1)); forvar1183 = (forvar1183 + (1'h1)))
        begin
          for (forvar1184 = (1'h0); (forvar1184 < (1'h0)); forvar1184 = (forvar1184 + (1'h1)))
            begin
              reg1185 <= ((reg1075[(2'h2):(1'h0)] ^ (((reg1099 ^ reg931) ^ ((8'h9d) ?
                  reg957 : reg1047)) & (reg947[(3'h4):(1'h0)] + reg1094))) >>> $unsigned(reg922));
            end
        end
      reg1186 <= {(({{reg1124},
              {reg1094}} > reg1041) || ($signed(reg1105[(1'h1):(1'h1)]) ?
              wire902 : ((reg1059 ~^ (8'hbe)) >>> reg916[(5'h15):(3'h5)])))};
      reg1187 = reg948;
      reg1188 <= (7'h49);
    end
  always
    @(posedge clk) begin
      for (forvar1189 = (1'h0); (forvar1189 < (3'h4)); forvar1189 = (forvar1189 + (1'h1)))
        begin
          for (forvar1190 = (1'h0); (forvar1190 < (3'h4)); forvar1190 = (forvar1190 + (1'h1)))
            begin
              reg1191 = $signed(reg1137[(2'h3):(2'h2)]);
              reg1192 <= ((~^{(!reg1008),
                      (((7'h42) ? wire1177 : reg1063) <= $unsigned(reg1094))}) ?
                  (!((~&$unsigned(reg1018)) | $unsigned((reg1191 && reg1018)))) : $unsigned((((wire1177 && reg988) && {reg933,
                          reg979}) ?
                      reg1185[(3'h6):(3'h4)] : {$signed(reg1053)})));
              reg1193 = $signed($unsigned(((-reg957[(3'h7):(2'h2)]) ?
                  ((reg1116 ?
                      reg1163 : wire1100) >>> reg1017) : $signed((&reg1011)))));
              reg1194 <= $unsigned($unsigned(reg952[(2'h2):(1'h0)]));
            end
          for (forvar1195 = (1'h0); (forvar1195 < (1'h0)); forvar1195 = (forvar1195 + (1'h1)))
            begin
              reg1196 <= reg960;
            end
          reg1197 = reg1009[(3'h5):(3'h4)];
          reg1198 = reg931[(2'h3):(1'h1)];
        end
      reg1199 = wire929;
      reg1200 <= (-$signed({($unsigned(reg1130) ?
              (reg1130 > reg1005) : $unsigned(wire1104)),
          $unsigned({reg1005, reg1165})}));
      for (forvar1201 = (1'h0); (forvar1201 < (2'h2)); forvar1201 = (forvar1201 + (1'h1)))
        begin
          if ($unsigned((reg1047[(3'h5):(3'h4)] + wire929[(2'h2):(2'h2)])))
            begin
              reg1202 <= ((+$unsigned($signed(reg1040[(4'ha):(4'h8)]))) ?
                  $unsigned($signed((~|(-reg955)))) : (wire1178 < {(+(7'h47))}));
              reg1203 = $unsigned($signed(reg1027[(3'h5):(1'h0)]));
            end
          else
            begin
              reg1202 <= $signed((reg1185 + $unsigned(reg992[(3'h5):(2'h3)])));
            end
          reg1204 = ($signed({$unsigned((reg1020 | reg1008)),
              reg911[(4'he):(4'h9)]}) << (($signed(reg984) ?
              $signed(reg916[(4'ha):(4'h8)]) : reg963[(4'hd):(2'h3)]) - $signed(reg1122[(4'hc):(4'ha)])));
          reg1205 <= reg1022[(4'he):(4'he)];
          for (forvar1206 = (1'h0); (forvar1206 < (1'h0)); forvar1206 = (forvar1206 + (1'h1)))
            begin
              reg1207 = reg1040[(4'ha):(4'h8)];
            end
          reg1208 <= reg1027;
        end
      for (forvar1209 = (1'h0); (forvar1209 < (1'h0)); forvar1209 = (forvar1209 + (1'h1)))
        begin
          for (forvar1210 = (1'h0); (forvar1210 < (3'h4)); forvar1210 = (forvar1210 + (1'h1)))
            begin
              reg1211 <= $unsigned(reg967);
              reg1212 <= {((reg1165[(4'hd):(4'h8)] & $signed((reg1202 >= reg1020))) == $signed($unsigned((7'h48))))};
              reg1213 = reg1075;
              reg1214 <= $signed(reg1022[(3'h5):(2'h2)]);
            end
          if ($unsigned(reg1130[(3'h6):(1'h1)]))
            begin
              reg1215 = (~|$unsigned($signed($unsigned({reg1130}))));
              reg1216 <= reg1073;
              reg1217 = reg1161[(4'hc):(4'ha)];
            end
          else
            begin
              reg1216 <= {(((reg1166[(4'hb):(3'h6)] >= reg947) ?
                          $signed(reg1109) : {(wire1181 ~^ reg1016),
                              $unsigned(forvar1209)}) ?
                      ((reg977[(4'hd):(2'h3)] ?
                          (reg914 ?
                              (7'h40) : reg1056) : ((8'hb4) | reg1009)) <<< ((wire1102 || reg1065) ?
                          reg967[(1'h1):(1'h1)] : reg1208)) : $unsigned(reg1028[(1'h1):(1'h0)])),
                  (reg1093[(1'h1):(1'h1)] ?
                      ((~$signed(reg1031)) > reg1056) : $signed(reg1130[(4'h9):(1'h1)]))};
              reg1217 = ($unsigned((+$signed(reg921[(2'h2):(1'h0)]))) ?
                  {reg915,
                      (reg1056[(3'h6):(3'h6)] ?
                          reg994[(3'h5):(1'h0)] : $unsigned((8'h9e)))} : reg955[(3'h6):(1'h1)]);
              reg1218 <= ({$signed(($signed(reg1139) <<< (+reg1020))),
                      ($signed((reg1144 - reg911)) ?
                          $unsigned($unsigned(reg1063)) : reg1170)} ?
                  {($signed($signed(reg918)) ?
                          ($signed(reg1031) <<< (forvar1206 ?
                              wire903 : (7'h48))) : reg1011),
                      (~^$signed($signed(reg1073)))} : ((reg1031 & $unsigned({reg1018})) - $unsigned({(wire1101 | reg1105),
                      (reg975 + reg915)})));
              reg1219 <= reg1002[(2'h2):(1'h1)];
            end
        end
    end
  assign wire1220 = (^reg1163[(2'h3):(2'h2)]);
  always
    @(posedge clk) begin
      for (forvar1221 = (1'h0); (forvar1221 < (3'h4)); forvar1221 = (forvar1221 + (1'h1)))
        begin
          if (reg1170)
            begin
              reg1222 <= reg1056;
              reg1223 = $unsigned((!(-reg1033[(1'h1):(1'h1)])));
              reg1224 <= (reg941[(3'h4):(1'h0)] ?
                  (^~$unsigned((8'hb0))) : reg1166[(5'h10):(2'h2)]);
              reg1225 = {(~|(reg952[(4'hc):(4'hc)] ?
                      (&reg1122[(3'h6):(3'h6)]) : $signed((reg1040 & reg1165))))};
            end
          else
            begin
              reg1222 <= $signed($unsigned((reg1061 <<< reg1211[(5'h10):(4'hd)])));
              reg1224 <= reg994[(4'hb):(1'h0)];
              reg1226 <= {(reg1113[(3'h5):(3'h5)] <= (+$signed(reg1152[(5'h11):(3'h5)])))};
              reg1227 = ($signed((^~{reg1008[(3'h7):(3'h4)]})) ^~ $unsigned($unsigned((reg1016[(3'h5):(1'h0)] ^ $unsigned((8'hb8))))));
              reg1228 <= reg956[(2'h3):(2'h3)];
            end
          for (forvar1229 = (1'h0); (forvar1229 < (2'h2)); forvar1229 = (forvar1229 + (1'h1)))
            begin
              reg1230 <= $signed(reg960);
              reg1231 = ($signed(((reg1219[(4'h8):(3'h7)] ?
                      (8'hb9) : reg1054[(4'h9):(2'h2)]) ?
                  ((reg947 ^ reg910) ?
                      (~reg1069) : reg976) : reg921)) ^ reg1069[(5'h13):(5'h12)]);
              reg1232 <= {reg950, $unsigned($signed(reg1230))};
              reg1233 = (^$unsigned({((reg1044 ? wire1220 : reg1119) ?
                      wire986 : (wire1101 != reg1018))}));
              reg1234 <= reg1057;
            end
          if (reg1096)
            begin
              reg1235 = (8'ha8);
            end
          else
            begin
              reg1235 = reg1058;
              reg1236 <= (7'h47);
              reg1237 <= ($signed(($signed({reg1200}) ?
                      reg1033 : {$signed((8'ha1))})) ?
                  (+(!(!$signed(reg1233)))) : reg931[(5'h10):(5'h10)]);
              reg1238 <= $signed((8'hba));
            end
        end
      reg1239 = reg1017[(3'h5):(2'h3)];
      reg1240 <= (&$unsigned((+$signed(reg988[(3'h5):(2'h3)]))));
      reg1241 = ($signed($signed($signed(reg992[(3'h6):(3'h5)]))) ?
          $signed((~|reg1238)) : $unsigned(reg918[(1'h1):(1'h0)]));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module619
#(parameter param784 = ((~&{(((8'hbd) || (8'h9c)) >> ((8'hbd) ? (8'haa) : (8'ha4))), ((~|(8'hb9)) ? ((8'hbc) <<< (7'h4a)) : {(8'ha4), (7'h4a)})}) ? {((-((7'h46) * (8'hb0))) ? (^(|(8'hbb))) : (~(8'ha8))), (~|((&(8'h9d)) ~^ (+(8'hb8))))} : (&(~^((|(8'h9f)) < (^(7'h49)))))), 
parameter param785 = param784)
(y, clk, wire624, wire623, wire622, wire621, wire620);
  output wire [(32'h840):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire624;
  input wire [(2'h2):(1'h0)] wire623;
  input wire signed [(3'h5):(1'h0)] wire622;
  input wire signed [(5'h12):(1'h0)] wire621;
  input wire [(5'h13):(1'h0)] wire620;
  wire signed [(2'h2):(1'h0)] wire783;
  wire signed [(4'hb):(1'h0)] wire782;
  wire [(4'hd):(1'h0)] wire766;
  wire signed [(4'hb):(1'h0)] wire765;
  wire signed [(4'hb):(1'h0)] wire632;
  wire [(5'h14):(1'h0)] wire631;
  wire signed [(2'h3):(1'h0)] wire630;
  reg signed [(4'he):(1'h0)] reg781 = (1'h0);
  reg [(4'h8):(1'h0)] reg780 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg779 = (1'h0);
  reg [(3'h4):(1'h0)] reg776 = (1'h0);
  reg [(2'h2):(1'h0)] reg773 = (1'h0);
  reg [(4'hb):(1'h0)] reg771 = (1'h0);
  reg [(5'h14):(1'h0)] reg770 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg764 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg763 = (1'h0);
  reg [(4'he):(1'h0)] reg762 = (1'h0);
  reg [(5'h16):(1'h0)] reg758 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg756 = (1'h0);
  reg [(4'he):(1'h0)] reg755 = (1'h0);
  reg [(4'he):(1'h0)] reg754 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg752 = (1'h0);
  reg signed [(4'he):(1'h0)] reg749 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg745 = (1'h0);
  reg [(3'h6):(1'h0)] reg744 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg742 = (1'h0);
  reg [(4'hb):(1'h0)] reg741 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg739 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg735 = (1'h0);
  reg [(5'h14):(1'h0)] reg733 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg731 = (1'h0);
  reg [(4'hf):(1'h0)] reg729 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg727 = (1'h0);
  reg [(4'he):(1'h0)] reg726 = (1'h0);
  reg [(5'h15):(1'h0)] reg725 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg722 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg719 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg716 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg713 = (1'h0);
  reg [(5'h11):(1'h0)] reg712 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg709 = (1'h0);
  reg [(5'h12):(1'h0)] reg705 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg704 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg701 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg700 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg699 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg697 = (1'h0);
  reg [(3'h4):(1'h0)] reg691 = (1'h0);
  reg [(4'ha):(1'h0)] reg689 = (1'h0);
  reg [(4'hd):(1'h0)] reg686 = (1'h0);
  reg [(4'hc):(1'h0)] reg682 = (1'h0);
  reg [(4'h8):(1'h0)] reg681 = (1'h0);
  reg [(5'h11):(1'h0)] reg677 = (1'h0);
  reg [(3'h4):(1'h0)] reg673 = (1'h0);
  reg [(4'ha):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg669 = (1'h0);
  reg [(3'h7):(1'h0)] reg666 = (1'h0);
  reg [(4'h8):(1'h0)] reg664 = (1'h0);
  reg [(5'h17):(1'h0)] reg663 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg657 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg655 = (1'h0);
  reg signed [(4'he):(1'h0)] reg654 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg650 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg649 = (1'h0);
  reg [(5'h12):(1'h0)] reg648 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg647 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg645 = (1'h0);
  reg [(5'h18):(1'h0)] reg643 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg642 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg641 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg639 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg636 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg633 = (1'h0);
  reg [(5'h11):(1'h0)] reg629 = (1'h0);
  reg [(4'h9):(1'h0)] reg628 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg627 = (1'h0);
  reg [(5'h16):(1'h0)] reg626 = (1'h0);
  reg [(3'h6):(1'h0)] reg778 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar777 = (1'h0);
  reg [(3'h6):(1'h0)] reg775 = (1'h0);
  reg [(4'hb):(1'h0)] reg774 = (1'h0);
  reg [(4'hc):(1'h0)] reg772 = (1'h0);
  reg [(4'hb):(1'h0)] reg767 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg769 = (1'h0);
  reg signed [(4'he):(1'h0)] reg768 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar767 = (1'h0);
  reg [(5'h18):(1'h0)] reg761 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar760 = (1'h0);
  reg [(2'h3):(1'h0)] reg759 = (1'h0);
  reg [(5'h16):(1'h0)] reg757 = (1'h0);
  reg [(5'h10):(1'h0)] reg753 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg751 = (1'h0);
  reg [(4'hd):(1'h0)] reg750 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg748 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg747 = (1'h0);
  reg [(5'h10):(1'h0)] reg746 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg743 = (1'h0);
  reg [(3'h6):(1'h0)] forvar740 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar738 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg737 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg736 = (1'h0);
  reg [(4'hb):(1'h0)] reg734 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg732 = (1'h0);
  reg [(5'h18):(1'h0)] forvar730 = (1'h0);
  reg signed [(4'he):(1'h0)] reg728 = (1'h0);
  reg [(5'h18):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg723 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg721 = (1'h0);
  reg [(4'hd):(1'h0)] reg720 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar718 = (1'h0);
  reg [(5'h16):(1'h0)] reg717 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg715 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg714 = (1'h0);
  reg [(2'h2):(1'h0)] reg711 = (1'h0);
  reg [(3'h5):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg708 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg707 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg706 = (1'h0);
  reg [(3'h4):(1'h0)] reg703 = (1'h0);
  reg signed [(4'he):(1'h0)] reg702 = (1'h0);
  reg [(5'h10):(1'h0)] reg696 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg695 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg694 = (1'h0);
  reg [(5'h11):(1'h0)] reg693 = (1'h0);
  reg [(4'h9):(1'h0)] reg692 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg690 = (1'h0);
  reg [(3'h5):(1'h0)] reg688 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg687 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg685 = (1'h0);
  reg [(3'h7):(1'h0)] forvar684 = (1'h0);
  reg [(5'h18):(1'h0)] reg683 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg680 = (1'h0);
  reg [(5'h11):(1'h0)] reg679 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar678 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg676 = (1'h0);
  reg [(5'h12):(1'h0)] reg675 = (1'h0);
  reg [(5'h17):(1'h0)] reg674 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar672 = (1'h0);
  reg [(5'h17):(1'h0)] forvar671 = (1'h0);
  reg [(3'h7):(1'h0)] reg668 = (1'h0);
  reg [(4'he):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg665 = (1'h0);
  reg [(3'h6):(1'h0)] reg662 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar660 = (1'h0);
  reg [(5'h11):(1'h0)] reg652 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg660 = (1'h0);
  reg [(2'h3):(1'h0)] reg658 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg656 = (1'h0);
  reg [(3'h7):(1'h0)] reg653 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar652 = (1'h0);
  reg [(5'h12):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg646 = (1'h0);
  reg [(4'hc):(1'h0)] reg644 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar641 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg634 = (1'h0);
  reg [(3'h4):(1'h0)] reg640 = (1'h0);
  reg [(5'h11):(1'h0)] reg638 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg637 = (1'h0);
  reg [(2'h2):(1'h0)] reg635 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar634 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar625 = (1'h0);
  assign y = {wire783,
                 wire782,
                 wire766,
                 wire765,
                 wire632,
                 wire631,
                 wire630,
                 reg781,
                 reg780,
                 reg779,
                 reg776,
                 reg773,
                 reg771,
                 reg770,
                 reg764,
                 reg763,
                 reg762,
                 reg758,
                 reg756,
                 reg755,
                 reg754,
                 reg752,
                 reg749,
                 reg745,
                 reg744,
                 reg742,
                 reg741,
                 reg739,
                 reg735,
                 reg733,
                 reg731,
                 reg729,
                 reg727,
                 reg726,
                 reg725,
                 reg722,
                 reg719,
                 reg716,
                 reg713,
                 reg712,
                 reg709,
                 reg705,
                 reg704,
                 reg701,
                 reg700,
                 reg699,
                 reg698,
                 reg697,
                 reg691,
                 reg689,
                 reg686,
                 reg682,
                 reg681,
                 reg677,
                 reg673,
                 reg670,
                 reg669,
                 reg666,
                 reg664,
                 reg663,
                 reg659,
                 reg657,
                 reg655,
                 reg654,
                 reg650,
                 reg649,
                 reg648,
                 reg647,
                 reg645,
                 reg643,
                 reg642,
                 reg641,
                 reg639,
                 reg636,
                 reg633,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg778,
                 forvar777,
                 reg775,
                 reg774,
                 reg772,
                 reg767,
                 reg769,
                 reg768,
                 forvar767,
                 reg761,
                 forvar760,
                 reg759,
                 reg757,
                 reg753,
                 reg751,
                 reg750,
                 reg748,
                 reg747,
                 reg746,
                 reg743,
                 forvar740,
                 forvar738,
                 reg737,
                 reg736,
                 reg734,
                 reg732,
                 forvar730,
                 reg728,
                 reg724,
                 reg723,
                 reg721,
                 reg720,
                 forvar718,
                 reg717,
                 reg715,
                 reg714,
                 reg711,
                 reg710,
                 reg708,
                 reg707,
                 reg706,
                 reg703,
                 reg702,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg690,
                 reg688,
                 reg687,
                 reg685,
                 forvar684,
                 reg683,
                 reg680,
                 reg679,
                 forvar678,
                 reg676,
                 reg675,
                 reg674,
                 forvar672,
                 forvar671,
                 reg668,
                 reg667,
                 reg665,
                 reg662,
                 reg661,
                 forvar660,
                 reg652,
                 reg660,
                 reg658,
                 reg656,
                 reg653,
                 forvar652,
                 reg651,
                 reg646,
                 reg644,
                 forvar641,
                 reg634,
                 reg640,
                 reg638,
                 reg637,
                 reg635,
                 forvar634,
                 forvar625,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar625 = (1'h0); (forvar625 < (1'h0)); forvar625 = (forvar625 + (1'h1)))
        begin
          reg626 <= $unsigned({{$signed($unsigned(wire622))}});
          reg627 <= wire621[(1'h1):(1'h0)];
          reg628 <= ($unsigned(reg627) ?
              $signed((wire624[(3'h7):(1'h0)] ^~ {(wire622 ? reg626 : reg627),
                  (|(7'h46))})) : (^~($unsigned($unsigned(wire621)) << (wire622[(2'h2):(2'h2)] || reg627))));
        end
      reg629 <= ((~&((~&reg628) * $unsigned((8'hb9)))) ?
          wire623[(2'h2):(2'h2)] : wire623);
    end
  assign wire630 = (|((reg627 ?
                           $unsigned((~^(8'hb0))) : ((~wire622) ^ (reg628 ?
                               (8'ha1) : reg629))) ?
                       wire620[(4'hc):(1'h1)] : (reg627 ?
                           ((wire623 && (7'h49)) ?
                               (reg626 ?
                                   reg627 : wire623) : wire622[(1'h0):(1'h0)]) : ($signed(reg626) & $unsigned((8'ha3))))));
  assign wire631 = ((!wire623) ?
                       ($signed(((wire624 ? reg627 : wire630) ?
                           ((7'h49) ? wire621 : reg626) : (wire630 ?
                               wire624 : reg626))) != {(reg627 ?
                               (reg627 ?
                                   wire624 : wire620) : $unsigned((8'hb3)))}) : $unsigned((reg627[(3'h4):(1'h1)] ?
                           $signed({wire624, wire621}) : wire620)));
  assign wire632 = $unsigned(reg629[(3'h6):(2'h3)]);
  always
    @(posedge clk) begin
      if ((-{reg629, (8'hb7)}))
        begin
          reg633 <= (~^$unsigned($unsigned(wire620[(4'hc):(4'ha)])));
          for (forvar634 = (1'h0); (forvar634 < (2'h3)); forvar634 = (forvar634 + (1'h1)))
            begin
              reg635 = (reg628[(3'h5):(3'h4)] ?
                  $unsigned((~(((8'hbc) ? wire630 : wire621) ?
                      (~^wire631) : wire621[(4'hd):(4'ha)]))) : ((wire624[(3'h7):(3'h4)] ?
                          $signed(reg627) : (8'hb5)) ?
                      (({(7'h47)} || (reg629 != wire631)) ?
                          ({wire623} ?
                              (&(8'ha3)) : wire623[(1'h0):(1'h0)]) : $signed($signed(wire624))) : (!(wire623[(1'h1):(1'h1)] ?
                          $unsigned(wire630) : $signed(wire623)))));
              reg636 <= $unsigned(wire620[(4'ha):(2'h3)]);
            end
          if (wire624[(4'hc):(1'h0)])
            begin
              reg637 = reg627[(1'h0):(1'h0)];
              reg638 = $unsigned(($unsigned($unsigned({wire621})) ^ $unsigned(($unsigned((8'haa)) ?
                  (wire620 * reg628) : $unsigned(reg636)))));
              reg639 <= {(reg636[(4'h8):(1'h1)] ?
                      (~^($signed((7'h41)) - $signed((8'ha1)))) : (((reg633 ?
                                  (8'hae) : wire630) ?
                              (&reg628) : (&reg628)) ?
                          ($unsigned(wire630) ^ $signed(reg627)) : (~(~^reg637)))),
                  (($unsigned((forvar634 < reg637)) > (^~((8'hb1) >= (7'h40)))) ?
                      (wire622 << ({reg638} ?
                          (wire630 ?
                              reg626 : wire623) : (^~wire631))) : $unsigned(((~&reg629) * {(8'ha0)})))};
              reg640 = wire632[(3'h4):(1'h0)];
              reg641 <= (reg628 || ((!wire630[(1'h1):(1'h0)]) ^~ reg627));
            end
          else
            begin
              reg637 = forvar634[(1'h1):(1'h0)];
              reg639 <= ($signed((reg628 ?
                      (-forvar634[(2'h2):(2'h2)]) : (reg637[(3'h5):(1'h1)] ^ (~^(8'hb8))))) ?
                  reg638[(3'h7):(1'h0)] : ({wire623[(1'h0):(1'h0)]} ~^ reg636[(1'h0):(1'h0)]));
              reg640 = (reg635[(2'h2):(1'h1)] * $unsigned((~|($unsigned((8'hbf)) ~^ (!reg640)))));
            end
        end
      else
        begin
          reg634 = (((8'hba) ?
                  ((8'hbf) ?
                      wire624[(4'ha):(3'h7)] : ($signed((8'haf)) ?
                          (wire632 <<< (8'hb8)) : $unsigned(wire632))) : reg640) ?
              $unsigned(reg629) : ($unsigned(($signed(wire621) ?
                      (wire620 <<< reg627) : $signed(wire630))) ?
                  ({$signed((7'h44)),
                      $signed(wire624)} ^ wire630[(1'h0):(1'h0)]) : (({(8'hb2),
                      reg626} >>> reg635) & $signed((&wire630)))));
          reg636 <= $unsigned((8'hba));
          if ($unsigned(((8'h9e) ?
              ((wire620[(4'hc):(2'h3)] ?
                  $unsigned(reg634) : reg627) | (-(reg639 << wire630))) : (($signed(wire624) ?
                  {wire631} : reg635[(1'h1):(1'h0)]) * $signed({reg641})))))
            begin
              reg639 <= ($signed($signed(((reg641 ? reg628 : reg637) ?
                  reg635[(1'h0):(1'h0)] : $unsigned(forvar634)))) + wire632);
              reg640 = {reg637};
            end
          else
            begin
              reg637 = reg638[(4'he):(3'h7)];
              reg638 = {$unsigned($signed(($signed(reg636) ?
                      $signed(wire624) : $unsigned(reg629)))),
                  $unsigned(wire621[(1'h1):(1'h1)])};
              reg639 <= (wire623[(1'h0):(1'h0)] <= (((!(wire624 < wire630)) - (~^(~&(8'ha2)))) <<< (+reg634)));
              reg640 = (reg635[(2'h2):(1'h0)] ?
                  reg636 : (^~wire620[(4'hd):(4'hc)]));
            end
          for (forvar641 = (1'h0); (forvar641 < (3'h4)); forvar641 = (forvar641 + (1'h1)))
            begin
              reg642 <= {reg635[(1'h0):(1'h0)], reg639[(4'hb):(4'hb)]};
              reg643 <= ((~|$signed(wire621[(1'h0):(1'h0)])) ?
                  $unsigned(reg635) : (((reg633[(1'h1):(1'h1)] ?
                          $unsigned(wire624) : {(7'h41)}) & reg633) ?
                      ((forvar634 == $unsigned(wire621)) ?
                          (^~{reg627,
                              wire623}) : $signed($signed(reg640))) : (((reg637 ?
                              (8'ha9) : reg629) ?
                          reg634 : (~^forvar641)) ^ wire630[(2'h2):(2'h2)])));
            end
          reg644 = (~&forvar634);
        end
    end
  always
    @(posedge clk) begin
      if ((&reg643))
        begin
          reg645 <= (reg627[(2'h3):(2'h3)] * (&$unsigned((reg626[(3'h7):(3'h5)] <= (wire632 ~^ reg643)))));
        end
      else
        begin
          reg645 <= $unsigned(((|(+(reg642 ~^ reg633))) < ($unsigned({reg627,
                  reg636}) ?
              ($signed((8'h9d)) ^ (reg639 ?
                  reg628 : (7'h49))) : (~^reg628[(2'h2):(1'h0)]))));
          if ((8'hb3))
            begin
              reg646 = (8'h9d);
              reg647 <= ((+(wire623[(1'h1):(1'h0)] ?
                  $unsigned((+wire632)) : ((~^reg642) >>> $unsigned(wire622)))) <<< $unsigned((+((reg646 ?
                  wire622 : (8'hbb)) < (|(7'h48))))));
              reg648 <= ($unsigned($signed({$signed((7'h45))})) ^~ $signed(((wire623 * reg643[(5'h15):(4'h8)]) >> $unsigned((wire621 ?
                  (8'hbc) : wire622)))));
            end
          else
            begin
              reg646 = ((((wire622 > (~&wire630)) ?
                      wire630[(2'h3):(1'h0)] : $signed($signed(wire624))) ?
                  $unsigned((~|(reg646 - reg645))) : {(wire622 != (reg628 ?
                          (8'h9d) : reg647)),
                      (~|{wire623})}) ^~ reg627);
            end
        end
      reg649 <= reg639[(5'h10):(4'hd)];
      reg650 <= reg646[(4'h8):(3'h6)];
      if ($signed({$unsigned({$signed(wire624)})}))
        begin
          reg651 = reg633[(3'h6):(3'h4)];
          for (forvar652 = (1'h0); (forvar652 < (1'h0)); forvar652 = (forvar652 + (1'h1)))
            begin
              reg653 = reg626;
              reg654 <= $unsigned(wire624[(5'h10):(4'hf)]);
              reg655 <= (($signed(reg629) ?
                      $unsigned((-$signed(reg645))) : (reg653[(3'h5):(1'h0)] ?
                          (~&{(7'h49), reg650}) : (reg626 < $signed(reg648)))) ?
                  $unsigned(($signed($signed(reg642)) ?
                      ((wire620 ? (8'h9f) : reg627) ?
                          $unsigned((8'hb1)) : (^~reg629)) : $signed({reg643}))) : $unsigned($unsigned((reg654[(4'hd):(3'h7)] && (~^(8'hb8))))));
            end
          reg656 = (reg655 ?
              ($signed((~|(~forvar652))) ?
                  $signed(wire623[(1'h1):(1'h1)]) : (^~$unsigned((^(8'hbd))))) : $unsigned($unsigned(wire632)));
          reg657 <= $signed(wire622[(3'h5):(2'h2)]);
          if ((reg655 ?
              (&$unsigned(((&reg650) | (reg645 - reg643)))) : $signed((^$signed({reg654,
                  reg656})))))
            begin
              reg658 = ($unsigned((reg650 - (reg639[(1'h0):(1'h0)] ^~ $signed(wire622)))) ?
                  wire630 : {$unsigned($unsigned((~&(8'hb8))))});
            end
          else
            begin
              reg658 = ({(^~{(reg649 ? reg649 : wire623)}),
                  (|$unsigned(reg658))} != reg633[(2'h3):(1'h0)]);
              reg659 <= reg655;
              reg660 = ((wire624[(4'ha):(2'h3)] - (&$unsigned(((7'h40) ?
                  wire630 : reg627)))) == $signed((wire632 ?
                  $unsigned((wire621 != (8'hb8))) : $signed((!reg633)))));
            end
        end
      else
        begin
          if ($unsigned((reg659 ?
              $unsigned({(+reg651), reg636[(1'h0):(1'h0)]}) : (+(((8'hb2) ?
                      wire621 : wire621) ?
                  {forvar652} : (reg636 ~^ reg646))))))
            begin
              reg651 = $unsigned((reg629 ?
                  wire623 : (~wire623[(1'h0):(1'h0)])));
              reg652 = $signed($unsigned(reg646[(4'hc):(3'h5)]));
              reg653 = reg651[(5'h12):(3'h4)];
              reg656 = (8'ha0);
              reg658 = $signed((8'haf));
            end
          else
            begin
              reg651 = wire620;
              reg654 <= reg659[(4'ha):(2'h2)];
              reg655 <= (reg639[(4'h8):(3'h5)] ?
                  $signed(reg650[(2'h3):(2'h2)]) : wire621[(5'h11):(1'h0)]);
              reg656 = $signed($signed((((reg628 << reg655) ?
                      reg656[(3'h4):(3'h4)] : $unsigned(reg642)) ?
                  (&(wire624 <<< reg639)) : ($unsigned(reg629) ?
                      (8'hb5) : reg636))));
            end
          reg659 <= (reg639[(4'ha):(3'h6)] ^~ (^$signed(reg654[(3'h7):(3'h5)])));
          for (forvar660 = (1'h0); (forvar660 < (2'h2)); forvar660 = (forvar660 + (1'h1)))
            begin
              reg661 = ($unsigned(((8'hae) != (reg651 <= (reg629 || forvar652)))) < $signed($unsigned((~|forvar652))));
              reg662 = (^(({(wire631 ? reg636 : reg661)} ?
                  ({reg627} * $unsigned((7'h49))) : (~&wire631)) + reg655[(2'h3):(1'h0)]));
              reg663 <= (+(((reg633[(4'h8):(2'h3)] ?
                      reg657 : $unsigned(reg653)) ?
                  ({reg651,
                      reg658} & (wire624 == wire622)) : {wire632}) ^~ {(~(!(8'ha5)))}));
              reg664 <= (((reg655 ?
                          wire620 : ($signed(reg646) ~^ $signed(forvar660))) ?
                      $signed((~|$unsigned(reg652))) : {($signed(reg648) ^~ $signed(reg649)),
                          ($unsigned(reg633) * reg642[(3'h6):(1'h0)])}) ?
                  $unsigned($unsigned((~|(reg661 ?
                      (7'h41) : reg662)))) : reg639[(2'h2):(1'h1)]);
            end
          reg665 = (~^(wire620 << (~{(reg652 << wire622)})));
          if ((^$unsigned(((+(~^reg657)) ?
              ((8'h9f) != (~reg649)) : (wire624[(3'h7):(1'h1)] ?
                  $signed(reg659) : (wire622 ? reg628 : reg663))))))
            begin
              reg666 <= forvar652[(3'h6):(2'h3)];
              reg667 = $unsigned(((($signed(reg654) || (^reg627)) * $unsigned((&reg665))) ?
                  $unsigned({reg649[(4'hb):(2'h3)]}) : $unsigned(((^wire623) | wire631[(5'h12):(3'h6)]))));
              reg668 = $unsigned($signed((reg626[(5'h13):(2'h2)] ?
                  ($signed(reg629) ?
                      (-reg645) : reg650[(4'he):(4'hc)]) : reg643)));
              reg669 <= ((&($signed($signed((8'ha6))) + ($unsigned(reg653) ?
                  (reg626 == reg649) : (wire624 ?
                      reg626 : reg657)))) << $unsigned(reg664[(1'h0):(1'h0)]));
              reg670 <= $signed(wire624);
            end
          else
            begin
              reg666 <= (((((reg641 ? wire631 : reg664) ?
                          {reg649} : {reg641, forvar652}) ?
                      ((~reg664) ?
                          (reg646 ~^ reg654) : forvar660) : $signed({wire620})) || (!((~&reg659) - (reg636 ?
                      (8'h9d) : reg641)))) ?
                  reg651[(3'h6):(2'h2)] : ($unsigned(wire620) ?
                      (reg626 - ($signed(wire620) ?
                          {reg668} : reg670)) : $signed(reg629[(1'h1):(1'h0)])));
              reg669 <= ((~^($unsigned($unsigned(reg668)) ?
                  $signed($unsigned(reg649)) : $unsigned(reg662))) >> wire624);
              reg670 <= (8'hb3);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar671 = (1'h0); (forvar671 < (2'h3)); forvar671 = (forvar671 + (1'h1)))
        begin
          for (forvar672 = (1'h0); (forvar672 < (2'h2)); forvar672 = (forvar672 + (1'h1)))
            begin
              reg673 <= (7'h47);
              reg674 = ($unsigned((~&({wire620} <= $unsigned(reg655)))) - forvar672);
              reg675 = (reg666[(1'h1):(1'h0)] <= (^~reg655));
            end
          reg676 = $signed($signed({(^reg659)}));
          reg677 <= ((reg663 ?
              (reg636 + (^reg639)) : (8'hb2)) * $unsigned((reg664 && reg670[(4'ha):(4'ha)])));
          for (forvar678 = (1'h0); (forvar678 < (2'h2)); forvar678 = (forvar678 + (1'h1)))
            begin
              reg679 = forvar678[(1'h0):(1'h0)];
              reg680 = (~|reg641[(2'h2):(1'h1)]);
              reg681 <= $signed((~^$signed(reg645[(1'h1):(1'h0)])));
              reg682 <= ({{($signed((8'ha2)) ?
                          (reg639 ?
                              reg666 : reg639) : wire624[(3'h6):(3'h5)])}} <= reg643[(4'hc):(4'hc)]);
              reg683 = $unsigned($signed(reg666));
            end
        end
      for (forvar684 = (1'h0); (forvar684 < (2'h2)); forvar684 = (forvar684 + (1'h1)))
        begin
          reg685 = ((reg676 ?
                  wire632 : {(~$signed(reg627)),
                      $unsigned(reg674[(5'h15):(4'hb)])}) ?
              {forvar672[(4'ha):(4'ha)]} : $unsigned(({$unsigned(reg659)} ?
                  reg682 : (+$signed(reg643)))));
          reg686 <= reg633;
          if (((reg681[(1'h0):(1'h0)] > $signed({reg686[(4'h8):(3'h5)]})) ?
              (reg629 ?
                  (reg675 ?
                      (reg683 + {reg673,
                          (8'hbc)}) : ($unsigned((8'h9c)) | reg669)) : reg673[(3'h4):(3'h4)]) : $signed(reg655[(1'h0):(1'h0)])))
            begin
              reg687 = $signed(reg675);
              reg688 = ({(($signed((8'h9d)) ?
                      reg647[(1'h1):(1'h1)] : reg664[(4'h8):(4'h8)]) ^~ $signed((&reg686)))} ^ $unsigned($unsigned((^reg686))));
              reg689 <= {reg685[(4'h9):(3'h5)], reg626};
              reg690 = {reg664};
            end
          else
            begin
              reg689 <= reg657[(3'h6):(2'h3)];
              reg691 <= $unsigned(wire632);
              reg692 = reg629[(3'h7):(3'h6)];
              reg693 = (!(+(7'h44)));
              reg694 = {reg647[(2'h3):(1'h0)]};
            end
          reg695 = (reg628 ? (7'h41) : (&$unsigned(reg649)));
        end
    end
  always
    @(posedge clk) begin
      if (reg641)
        begin
          reg696 = reg689[(1'h0):(1'h0)];
        end
      else
        begin
          reg697 <= $signed((wire620 ?
              ($signed($signed(reg650)) ?
                  wire632 : reg629[(4'ha):(3'h7)]) : (|$signed((reg639 == wire623)))));
          if (reg682)
            begin
              reg698 <= reg655;
              reg699 <= $unsigned(reg636[(3'h6):(2'h2)]);
              reg700 <= ($unsigned((wire621[(2'h2):(2'h2)] > (8'ha6))) ?
                  (~&reg697[(4'h9):(3'h6)]) : (!reg628));
              reg701 <= wire632[(1'h0):(1'h0)];
            end
          else
            begin
              reg702 = (($signed((reg641 ?
                      (+reg682) : (wire630 ?
                          (8'ha8) : wire624))) || $signed(reg664)) ?
                  $signed((({reg626} ?
                          $signed((8'ha1)) : (wire632 ? reg677 : reg628)) ?
                      $signed((reg682 ? reg641 : reg666)) : {reg648,
                          (!(8'hb2))})) : $unsigned(($unsigned((reg663 - wire630)) || ((|reg626) ?
                      ((8'ha0) | (7'h49)) : (^wire624)))));
              reg703 = (^reg628[(4'h8):(3'h6)]);
            end
          if (reg682)
            begin
              reg704 <= ((~{{{(8'hbd)}, (reg669 ~^ reg657)},
                      $unsigned((reg657 ? reg641 : reg659))}) ?
                  reg627 : reg702);
              reg705 <= $unsigned(reg703[(2'h2):(2'h2)]);
            end
          else
            begin
              reg706 = ((reg700 ?
                  (~|$unsigned((reg666 ?
                      wire631 : (8'hbb)))) : (8'hb9)) ^~ (&reg626));
              reg707 = {(~($unsigned((-reg696)) ?
                      $unsigned((+reg659)) : {$unsigned(reg639)})),
                  reg706[(3'h6):(3'h6)]};
              reg708 = ((($signed(wire623) ?
                          $unsigned((reg628 ?
                              (8'ha5) : (8'h9d))) : $signed((~|reg703))) ?
                      ((reg643 ? $signed(reg654) : $unsigned(reg669)) ?
                          $signed((~^reg701)) : wire624) : reg706) ?
                  (~^$unsigned(reg628)) : {(^$unsigned($unsigned(reg673)))});
              reg709 <= (~&{((((8'hb7) | reg682) <<< (8'h9f)) || (!reg673))});
              reg710 = (8'hba);
            end
          if (($unsigned((&(^{reg700, (8'hab)}))) ?
              $unsigned($signed((8'hab))) : ({wire630,
                  (-(~&(7'h45)))} + $unsigned(reg655[(3'h5):(2'h3)]))))
            begin
              reg711 = (reg654 || $unsigned(({(^(8'hb9))} ?
                  (reg628 >> reg689[(4'h9):(2'h3)]) : reg704)));
              reg712 <= $signed(reg708);
              reg713 <= $signed($unsigned(($unsigned({reg628}) ?
                  $unsigned(reg657) : reg673)));
              reg714 = ($signed((!{$signed(reg706),
                  reg649})) < $signed(reg691));
              reg715 = (8'h9d);
            end
          else
            begin
              reg711 = (^~reg697);
              reg714 = reg703;
              reg715 = reg650[(4'hc):(4'h8)];
              reg716 <= reg641[(1'h1):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg717 = $signed(($unsigned($signed((~reg689))) + (reg705[(3'h6):(3'h5)] ?
          {$signed(wire631), reg716[(4'hd):(3'h6)]} : (7'h41))));
      for (forvar718 = (1'h0); (forvar718 < (1'h1)); forvar718 = (forvar718 + (1'h1)))
        begin
          reg719 <= (reg641 * wire624);
          reg720 = (&(~(((reg704 * reg642) ^~ $signed((8'h9c))) << wire630[(1'h1):(1'h0)])));
          reg721 = $signed(($unsigned($signed((reg670 ? reg663 : reg643))) ?
              (8'hb5) : reg713));
          if (((-(~&$signed((-(8'h9f))))) && $signed(reg628)))
            begin
              reg722 <= reg654;
            end
          else
            begin
              reg722 <= (~(reg717 || (wire622[(3'h4):(1'h1)] ?
                  reg704 : reg643[(4'hc):(3'h5)])));
              reg723 = {$signed((reg670[(3'h5):(2'h2)] >= reg689[(2'h3):(2'h3)]))};
            end
          if ($unsigned($unsigned(reg647[(1'h1):(1'h0)])))
            begin
              reg724 = (((~(reg639[(4'hd):(4'h9)] ?
                          $signed(reg691) : (~&reg677))) ?
                      $signed(reg682[(1'h0):(1'h0)]) : (~^{(reg717 ^~ wire631)})) ?
                  (|(reg701[(4'he):(1'h0)] == $signed(wire623[(1'h1):(1'h0)]))) : (!$signed($signed($signed(reg641)))));
              reg725 <= $unsigned($unsigned((|{reg673[(1'h1):(1'h0)]})));
              reg726 <= $unsigned(reg663[(3'h7):(1'h1)]);
              reg727 <= (wire632 ?
                  ((reg659 ?
                          $unsigned(reg670[(3'h6):(2'h3)]) : reg627[(2'h3):(1'h0)]) ?
                      $unsigned(reg724) : (|(reg712 + reg659))) : $signed((($unsigned(reg666) ?
                          (reg697 == reg642) : $signed((8'ha4))) ?
                      $unsigned(((8'haf) ?
                          reg689 : reg721)) : {(reg701 >> (7'h42))})));
              reg728 = ($unsigned(({(^~wire620)} ?
                  ((reg663 >>> wire630) ? {reg716} : reg719) : ((7'h4a) ?
                      $unsigned(reg670) : (reg627 - wire622)))) + (reg636 + reg636[(2'h3):(1'h1)]));
            end
          else
            begin
              reg725 <= $signed(forvar718);
              reg726 <= reg677;
              reg727 <= $unsigned($signed($unsigned((8'hbe))));
              reg728 = $unsigned(($unsigned(({(8'hb2)} ? (!reg629) : reg712)) ?
                  reg698 : (8'hb8)));
              reg729 <= $unsigned(((((reg697 <= reg673) <<< $signed(reg709)) >= $signed((8'hac))) && $signed(($unsigned(reg705) < reg670[(3'h4):(1'h1)]))));
            end
        end
      for (forvar730 = (1'h0); (forvar730 < (2'h2)); forvar730 = (forvar730 + (1'h1)))
        begin
          if ((wire630[(1'h1):(1'h1)] ?
              ($unsigned({(wire624 ? reg717 : reg727),
                  wire621}) >>> ($unsigned((forvar730 ~^ reg691)) ?
                  reg673[(1'h0):(1'h0)] : (reg633[(3'h7):(3'h5)] | $signed(reg669)))) : $unsigned(reg670)))
            begin
              reg731 <= wire623[(1'h0):(1'h0)];
              reg732 = reg700;
              reg733 <= $signed(((^~reg626) ?
                  $signed({reg705[(1'h1):(1'h0)]}) : (&reg650)));
            end
          else
            begin
              reg731 <= $signed(($signed(reg713) ?
                  $signed(($unsigned((8'hac)) ?
                      reg698 : reg642)) : ($signed($unsigned(reg673)) == $unsigned((reg627 & forvar730)))));
              reg732 = wire630[(2'h3):(1'h0)];
              reg734 = (!({reg666, reg717[(5'h12):(1'h1)]} ?
                  $signed(reg725) : $signed((~(~&reg686)))));
              reg735 <= ((reg669 ?
                      reg689[(2'h2):(2'h2)] : ($unsigned((~^(8'hbc))) ?
                          reg713 : ((reg719 ^~ (8'haa)) <<< {reg677}))) ?
                  reg686[(3'h7):(3'h5)] : (^~reg713));
              reg736 = reg726;
            end
          reg737 = wire631;
        end
      for (forvar738 = (1'h0); (forvar738 < (3'h4)); forvar738 = (forvar738 + (1'h1)))
        begin
          reg739 <= reg691;
          for (forvar740 = (1'h0); (forvar740 < (2'h3)); forvar740 = (forvar740 + (1'h1)))
            begin
              reg741 <= (|reg736);
              reg742 <= $unsigned($signed(reg659));
              reg743 = ($signed($unsigned(((~wire622) - reg739))) ?
                  $signed(((^$unsigned((8'hb5))) >> reg717[(5'h11):(4'hb)])) : (~^(((+(8'hb4)) ~^ {(8'hba),
                      forvar740}) <<< forvar730)));
              reg744 <= (~|(reg643 ?
                  reg732 : $signed($signed($unsigned((8'hb2))))));
            end
          reg745 <= ($unsigned(reg699[(3'h6):(3'h5)]) ?
              $unsigned(((~^reg670[(3'h7):(2'h2)]) ?
                  $signed(reg716[(4'hb):(3'h6)]) : reg677[(4'hd):(3'h4)])) : (reg732[(4'he):(4'h8)] >> (8'hba)));
        end
      if (((~&(wire621[(4'h8):(2'h2)] ?
              $unsigned((~(8'ha4))) : ((reg697 <= reg628) - reg726))) ?
          $unsigned($unsigned($signed(((8'hb3) ? reg717 : reg626)))) : wire632))
        begin
          if ((~^((|(&reg681)) ?
              ($signed(reg628[(3'h7):(3'h5)]) ^ ((reg720 ?
                  reg659 : (7'h40)) <<< (reg726 ?
                  reg666 : wire631))) : $signed($signed({(8'h9f)})))))
            begin
              reg746 = $signed(reg719);
              reg747 = reg627;
              reg748 = ($signed(($unsigned((~&wire624)) ?
                      reg689[(2'h2):(1'h0)] : ((~|reg699) & (reg726 ~^ reg725)))) ?
                  $signed(reg720) : reg736[(1'h1):(1'h1)]);
              reg749 <= ((^(+$unsigned($signed(reg746)))) < (reg737[(4'ha):(4'h8)] ?
                  ({reg723[(5'h11):(4'he)],
                      (reg729 ?
                          reg726 : reg664)} & ($unsigned((8'hbb)) == reg663)) : (-reg657)));
            end
          else
            begin
              reg749 <= reg699[(3'h5):(2'h3)];
              reg750 = ($signed($unsigned(reg726)) << $unsigned({(7'h43)}));
              reg751 = ($signed((8'hab)) ?
                  $unsigned({$signed((~reg669)),
                      reg698[(2'h2):(2'h2)]}) : (reg663[(1'h1):(1'h1)] <<< reg734));
              reg752 <= ($unsigned(reg748) >= (~reg737));
            end
          reg753 = {$unsigned(reg689), (wire621 == {reg682})};
          reg754 <= ((reg739[(3'h6):(2'h2)] | $signed($signed({reg716,
                  reg716}))) ?
              forvar730[(4'he):(4'hc)] : $unsigned(reg743[(4'hd):(1'h0)]));
          if ((|($signed(((reg724 ? reg735 : (7'h47)) * {reg734})) ?
              ({reg699[(3'h5):(1'h0)]} >> reg633) : $signed($unsigned((reg657 ?
                  reg720 : reg750))))))
            begin
              reg755 <= (~^($signed(reg726[(2'h3):(1'h1)]) ?
                  forvar738 : (8'h9f)));
              reg756 <= $signed($signed((8'ha8)));
              reg757 = (~|$unsigned(reg669));
            end
          else
            begin
              reg755 <= wire623;
              reg757 = $unsigned(forvar718[(4'hd):(4'hc)]);
              reg758 <= ($unsigned(($unsigned((reg689 ? (8'ha5) : (7'h46))) ?
                      (((7'h49) ? wire622 : reg633) ?
                          (reg670 ?
                              (8'ha7) : reg664) : (~|reg722)) : (!(^~reg743)))) ?
                  (+$unsigned($signed(reg709))) : $unsigned(reg673[(2'h3):(2'h2)]));
            end
        end
      else
        begin
          reg749 <= (8'hbe);
          if ($unsigned(((((forvar730 ?
                  (8'ha6) : reg659) == $unsigned((7'h46))) && wire624) ?
              (8'h9d) : $signed(($unsigned(reg734) ?
                  $signed(reg744) : {reg721})))))
            begin
              reg750 = ((({$signed(reg732), $signed(forvar738)} ?
                      reg691[(1'h1):(1'h1)] : ((8'ha8) ^~ $signed(reg757))) < $signed(reg681)) ?
                  $signed(((!{wire621}) != reg709)) : $unsigned($unsigned((|$signed(wire632)))));
              reg752 <= reg722[(3'h4):(1'h0)];
              reg754 <= (^(~^(-(!reg754[(4'hb):(4'h9)]))));
            end
          else
            begin
              reg752 <= reg745;
              reg753 = $unsigned($unsigned({(^reg704[(1'h1):(1'h1)])}));
              reg754 <= ((wire620 ?
                      $signed((!((8'hbe) ? (8'hb1) : reg689))) : reg682) ?
                  $unsigned(((-{reg756}) ?
                      reg722 : ($signed(reg735) == (reg754 >= reg720)))) : $signed(($signed($unsigned(reg729)) >>> reg701[(4'h9):(2'h2)])));
              reg757 = ($unsigned(forvar718) ?
                  ($signed(forvar738) != $signed(reg741)) : (~^(~$unsigned(reg723[(2'h3):(2'h3)]))));
            end
          reg759 = (reg758 ?
              reg734 : $signed((((|reg736) ?
                  {reg641,
                      (8'ha4)} : reg757[(3'h5):(3'h5)]) & ($unsigned(wire631) || (reg712 >>> reg628)))));
          for (forvar760 = (1'h0); (forvar760 < (2'h3)); forvar760 = (forvar760 + (1'h1)))
            begin
              reg761 = reg691[(1'h0):(1'h0)];
              reg762 <= ((~&$unsigned(reg732)) + (reg727 ?
                  ($unsigned((^(8'h9c))) >= (reg648[(4'he):(4'ha)] ?
                      ((7'h43) ? reg719 : reg720) : (reg629 ?
                          reg657 : reg721))) : $unsigned($unsigned(((7'h44) && forvar718)))));
              reg763 <= {{(~$unsigned($signed(reg698)))},
                  (!(reg753 & $signed((reg761 ? wire622 : reg759))))};
              reg764 <= (reg755[(1'h1):(1'h0)] && ($signed((+$unsigned(reg689))) ?
                  (((reg650 ?
                      reg682 : reg754) > $unsigned(wire630)) <<< reg756) : (reg666 < $signed(wire623))));
            end
        end
    end
  assign wire765 = (^~$signed((({reg729, reg705} >= (reg639 ?
                       reg641 : (8'hb6))) || $unsigned((reg643 ?
                       reg628 : reg689)))));
  assign wire766 = ($unsigned(($unsigned((reg650 * (8'hbc))) <<< $signed(reg756[(3'h4):(1'h1)]))) ?
                       $unsigned(({{reg744, reg686}} ^~ {reg655,
                           (^(8'hb7))})) : ((((^~reg727) >= $signed((8'had))) ?
                           $unsigned($unsigned(wire620)) : $unsigned(reg756[(4'hf):(4'hc)])) ~^ reg698));
  always
    @(posedge clk) begin
      if (wire630[(1'h1):(1'h0)])
        begin
          for (forvar767 = (1'h0); (forvar767 < (1'h0)); forvar767 = (forvar767 + (1'h1)))
            begin
              reg768 = (reg739[(2'h3):(2'h2)] * ((7'h4a) >> {($unsigned(reg716) ?
                      (-reg626) : ((7'h4a) ? reg691 : wire766)),
                  $signed(reg691[(1'h0):(1'h0)])}));
              reg769 = (~&((-$signed({wire620})) > reg719[(5'h12):(3'h5)]));
            end
          if (wire621[(2'h2):(2'h2)])
            begin
              reg770 <= reg677;
              reg771 <= (wire766 <= reg762);
            end
          else
            begin
              reg770 <= wire624[(4'hb):(4'hb)];
              reg771 <= $signed($unsigned($unsigned((8'hb4))));
            end
        end
      else
        begin
          reg767 = $signed(reg655);
          reg770 <= ($signed($signed($signed(reg699))) >>> reg770);
          if ($unsigned($signed(reg628[(1'h1):(1'h0)])))
            begin
              reg772 = wire620[(4'h9):(2'h2)];
              reg773 <= reg673;
              reg774 = (($unsigned({reg713[(3'h6):(2'h3)],
                  (reg649 ? wire623 : reg741)}) >>> {(~&reg666)}) == reg756);
              reg775 = (8'ha0);
            end
          else
            begin
              reg772 = reg712;
              reg774 = reg775;
              reg775 = ($signed($signed((~&{reg727}))) ?
                  (^(~&reg627)) : (!$signed(((-reg762) ?
                      ((7'h47) ? reg664 : reg725) : reg627))));
              reg776 <= (!$signed($signed(wire622)));
            end
          for (forvar777 = (1'h0); (forvar777 < (2'h2)); forvar777 = (forvar777 + (1'h1)))
            begin
              reg778 = {((8'ha8) << (({reg639, reg731} ?
                          (-wire620) : (reg769 ? reg754 : reg713)) ?
                      reg645 : reg686))};
              reg779 <= ($signed(reg629) != (reg659[(1'h1):(1'h0)] && ($signed((8'ha7)) ?
                  ((reg647 <<< reg722) >> ((8'hb2) ?
                      reg691 : reg745)) : {((8'hbc) ~^ reg626)})));
            end
        end
      reg780 <= ((~$unsigned(((reg677 ? reg762 : reg681) ?
              reg698 : reg769[(3'h7):(2'h2)]))) ?
          (&reg745) : {$signed(($unsigned(reg741) ?
                  (~^wire765) : (reg739 == reg770))),
              $signed($unsigned(((8'had) != reg733)))});
      reg781 <= wire630[(1'h1):(1'h1)];
    end
  assign wire782 = $signed((($signed($unsigned(reg666)) * $unsigned((^reg697))) && {reg764,
                       (reg657 ~^ (reg726 << (7'h42)))}));
  assign wire783 = reg713[(3'h4):(3'h4)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module255
#(parameter param615 = {{{((~|(8'haa)) & (^(8'hb5))), (((8'had) < (8'haa)) ~^ {(8'hbd)})}, (+((&(8'h9f)) ? (-(7'h4a)) : ((8'hb6) ? (8'hb8) : (8'ha3))))}})
(y, clk, wire259, wire258, wire257, wire256);
  output wire [(32'h1265):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h18):(1'h0)] wire259;
  input wire [(3'h6):(1'h0)] wire258;
  input wire signed [(4'hb):(1'h0)] wire257;
  input wire [(3'h4):(1'h0)] wire256;
  wire [(5'h12):(1'h0)] wire614;
  wire [(4'he):(1'h0)] wire613;
  wire signed [(4'h9):(1'h0)] wire612;
  wire [(2'h2):(1'h0)] wire583;
  wire signed [(3'h7):(1'h0)] wire542;
  wire signed [(4'hd):(1'h0)] wire541;
  wire signed [(4'hb):(1'h0)] wire457;
  wire signed [(5'h11):(1'h0)] wire436;
  wire signed [(4'h8):(1'h0)] wire435;
  wire signed [(4'hd):(1'h0)] wire370;
  wire signed [(5'h11):(1'h0)] wire342;
  reg [(4'hc):(1'h0)] reg609 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg607 = (1'h0);
  reg [(5'h14):(1'h0)] reg604 = (1'h0);
  reg [(5'h18):(1'h0)] reg601 = (1'h0);
  reg [(4'hc):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg598 = (1'h0);
  reg [(4'hd):(1'h0)] reg595 = (1'h0);
  reg [(3'h4):(1'h0)] reg593 = (1'h0);
  reg [(5'h15):(1'h0)] reg591 = (1'h0);
  reg [(3'h5):(1'h0)] reg590 = (1'h0);
  reg [(5'h11):(1'h0)] reg585 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg584 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg582 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg579 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg578 = (1'h0);
  reg [(3'h4):(1'h0)] reg576 = (1'h0);
  reg [(3'h5):(1'h0)] reg574 = (1'h0);
  reg [(3'h7):(1'h0)] reg573 = (1'h0);
  reg [(4'ha):(1'h0)] reg572 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg569 = (1'h0);
  reg [(2'h2):(1'h0)] reg567 = (1'h0);
  reg [(4'hb):(1'h0)] reg566 = (1'h0);
  reg [(5'h14):(1'h0)] reg565 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg560 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg558 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg553 = (1'h0);
  reg [(3'h4):(1'h0)] reg544 = (1'h0);
  reg [(4'hf):(1'h0)] reg551 = (1'h0);
  reg [(5'h13):(1'h0)] reg549 = (1'h0);
  reg [(3'h5):(1'h0)] reg546 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg545 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg543 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg539 = (1'h0);
  reg [(5'h16):(1'h0)] reg537 = (1'h0);
  reg [(4'hd):(1'h0)] reg536 = (1'h0);
  reg [(2'h2):(1'h0)] reg531 = (1'h0);
  reg [(4'h8):(1'h0)] reg526 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg520 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg528 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg517 = (1'h0);
  reg [(5'h10):(1'h0)] reg516 = (1'h0);
  reg [(2'h2):(1'h0)] reg514 = (1'h0);
  reg [(2'h3):(1'h0)] reg512 = (1'h0);
  reg [(5'h12):(1'h0)] reg510 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg508 = (1'h0);
  reg signed [(4'he):(1'h0)] reg504 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg503 = (1'h0);
  reg signed [(4'he):(1'h0)] reg502 = (1'h0);
  reg [(5'h10):(1'h0)] reg501 = (1'h0);
  reg [(3'h6):(1'h0)] reg500 = (1'h0);
  reg [(4'ha):(1'h0)] reg496 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg494 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg489 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg485 = (1'h0);
  reg [(5'h15):(1'h0)] reg481 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg478 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg476 = (1'h0);
  reg [(3'h7):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg469 = (1'h0);
  reg [(4'hc):(1'h0)] reg463 = (1'h0);
  reg [(4'hb):(1'h0)] reg465 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg461 = (1'h0);
  reg [(5'h13):(1'h0)] reg459 = (1'h0);
  reg [(5'h12):(1'h0)] reg455 = (1'h0);
  reg [(5'h18):(1'h0)] reg454 = (1'h0);
  reg [(3'h5):(1'h0)] reg452 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg450 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg444 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg441 = (1'h0);
  reg [(4'ha):(1'h0)] reg440 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg437 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg431 = (1'h0);
  reg [(5'h11):(1'h0)] reg433 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg429 = (1'h0);
  reg [(4'hf):(1'h0)] reg427 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg426 = (1'h0);
  reg [(5'h17):(1'h0)] reg423 = (1'h0);
  reg [(4'h9):(1'h0)] reg420 = (1'h0);
  reg [(3'h7):(1'h0)] reg418 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg415 = (1'h0);
  reg [(4'h8):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg409 = (1'h0);
  reg [(3'h4):(1'h0)] reg408 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg399 = (1'h0);
  reg [(5'h16):(1'h0)] reg397 = (1'h0);
  reg [(2'h3):(1'h0)] reg392 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg389 = (1'h0);
  reg [(3'h5):(1'h0)] reg388 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg385 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg384 = (1'h0);
  reg [(4'ha):(1'h0)] reg379 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg374 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg373 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg369 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg368 = (1'h0);
  reg [(5'h11):(1'h0)] reg367 = (1'h0);
  reg [(3'h4):(1'h0)] reg366 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg364 = (1'h0);
  reg [(4'hb):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg356 = (1'h0);
  reg [(2'h3):(1'h0)] reg355 = (1'h0);
  reg [(4'he):(1'h0)] reg350 = (1'h0);
  reg [(5'h14):(1'h0)] reg348 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg345 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg344 = (1'h0);
  reg [(4'ha):(1'h0)] reg343 = (1'h0);
  reg [(4'h8):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg339 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg334 = (1'h0);
  reg [(5'h15):(1'h0)] reg332 = (1'h0);
  reg [(3'h7):(1'h0)] reg330 = (1'h0);
  reg [(5'h16):(1'h0)] reg329 = (1'h0);
  reg [(5'h14):(1'h0)] reg328 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg327 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg325 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg322 = (1'h0);
  reg [(5'h10):(1'h0)] reg320 = (1'h0);
  reg [(4'ha):(1'h0)] reg319 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg318 = (1'h0);
  reg [(5'h17):(1'h0)] reg317 = (1'h0);
  reg [(4'h8):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg314 = (1'h0);
  reg [(4'h8):(1'h0)] reg313 = (1'h0);
  reg [(4'hc):(1'h0)] reg311 = (1'h0);
  reg [(3'h7):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg309 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg305 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg297 = (1'h0);
  reg [(5'h14):(1'h0)] reg301 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg300 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg299 = (1'h0);
  reg [(4'hc):(1'h0)] reg298 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg289 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg292 = (1'h0);
  reg [(5'h16):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg290 = (1'h0);
  reg [(2'h2):(1'h0)] reg287 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg285 = (1'h0);
  reg [(3'h5):(1'h0)] reg282 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg278 = (1'h0);
  reg [(3'h7):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg273 = (1'h0);
  reg [(3'h5):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg269 = (1'h0);
  reg [(3'h7):(1'h0)] reg266 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar605 = (1'h0);
  reg [(4'hc):(1'h0)] reg611 = (1'h0);
  reg [(4'h9):(1'h0)] reg610 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg608 = (1'h0);
  reg [(5'h17):(1'h0)] reg606 = (1'h0);
  reg [(4'hd):(1'h0)] reg605 = (1'h0);
  reg [(5'h13):(1'h0)] reg603 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg602 = (1'h0);
  reg [(3'h7):(1'h0)] reg599 = (1'h0);
  reg [(4'hf):(1'h0)] reg597 = (1'h0);
  reg [(4'hc):(1'h0)] reg596 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar593 = (1'h0);
  reg [(5'h11):(1'h0)] reg594 = (1'h0);
  reg [(4'he):(1'h0)] reg592 = (1'h0);
  reg [(2'h2):(1'h0)] reg589 = (1'h0);
  reg [(4'hb):(1'h0)] reg588 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg587 = (1'h0);
  reg [(4'h8):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar581 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg580 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar577 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg575 = (1'h0);
  reg signed [(4'he):(1'h0)] reg571 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg568 = (1'h0);
  reg [(5'h14):(1'h0)] forvar564 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg561 = (1'h0);
  reg [(5'h10):(1'h0)] reg559 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg557 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg556 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg555 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg554 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar552 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg548 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg550 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar548 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg547 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar544 = (1'h0);
  reg [(3'h4):(1'h0)] reg540 = (1'h0);
  reg [(4'h8):(1'h0)] forvar538 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg535 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg534 = (1'h0);
  reg [(5'h12):(1'h0)] forvar533 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg530 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar516 = (1'h0);
  reg [(4'hd):(1'h0)] reg527 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar526 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg525 = (1'h0);
  reg [(5'h14):(1'h0)] reg524 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg523 = (1'h0);
  reg [(3'h6):(1'h0)] reg522 = (1'h0);
  reg [(5'h14):(1'h0)] reg521 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar520 = (1'h0);
  reg signed [(4'he):(1'h0)] reg519 = (1'h0);
  reg [(5'h13):(1'h0)] reg518 = (1'h0);
  reg [(4'h8):(1'h0)] reg515 = (1'h0);
  reg [(5'h17):(1'h0)] forvar513 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg511 = (1'h0);
  reg [(5'h18):(1'h0)] reg509 = (1'h0);
  reg [(4'h9):(1'h0)] reg507 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar506 = (1'h0);
  reg [(5'h18):(1'h0)] reg505 = (1'h0);
  reg [(4'hc):(1'h0)] reg499 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg498 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar497 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg495 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg493 = (1'h0);
  reg [(4'hc):(1'h0)] forvar492 = (1'h0);
  reg [(4'h9):(1'h0)] reg491 = (1'h0);
  reg [(4'hc):(1'h0)] reg490 = (1'h0);
  reg [(2'h2):(1'h0)] reg488 = (1'h0);
  reg [(5'h11):(1'h0)] reg487 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar486 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg484 = (1'h0);
  reg [(4'h9):(1'h0)] reg483 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg482 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg480 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg479 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar477 = (1'h0);
  reg [(5'h10):(1'h0)] forvar475 = (1'h0);
  reg [(5'h13):(1'h0)] reg474 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar473 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg471 = (1'h0);
  reg [(5'h10):(1'h0)] forvar470 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg460 = (1'h0);
  reg [(5'h12):(1'h0)] reg468 = (1'h0);
  reg [(5'h14):(1'h0)] reg467 = (1'h0);
  reg [(3'h4):(1'h0)] reg466 = (1'h0);
  reg [(2'h3):(1'h0)] reg464 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar463 = (1'h0);
  reg [(4'he):(1'h0)] reg462 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar460 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg458 = (1'h0);
  reg [(4'hd):(1'h0)] reg456 = (1'h0);
  reg [(5'h15):(1'h0)] reg453 = (1'h0);
  reg [(4'h9):(1'h0)] reg451 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg447 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar446 = (1'h0);
  reg [(3'h6):(1'h0)] reg445 = (1'h0);
  reg [(2'h3):(1'h0)] reg443 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg439 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar438 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg434 = (1'h0);
  reg [(5'h17):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar431 = (1'h0);
  reg [(5'h12):(1'h0)] reg430 = (1'h0);
  reg [(5'h10):(1'h0)] reg428 = (1'h0);
  reg [(2'h2):(1'h0)] reg425 = (1'h0);
  reg [(5'h18):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar422 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg421 = (1'h0);
  reg [(4'hd):(1'h0)] forvar419 = (1'h0);
  reg [(5'h17):(1'h0)] reg417 = (1'h0);
  reg [(4'he):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg412 = (1'h0);
  reg [(4'he):(1'h0)] reg411 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg410 = (1'h0);
  reg [(2'h2):(1'h0)] forvar399 = (1'h0);
  reg [(4'hf):(1'h0)] reg407 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg404 = (1'h0);
  reg [(4'hb):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg402 = (1'h0);
  reg [(5'h15):(1'h0)] reg401 = (1'h0);
  reg signed [(4'he):(1'h0)] reg400 = (1'h0);
  reg [(5'h14):(1'h0)] reg398 = (1'h0);
  reg [(5'h16):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg395 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg394 = (1'h0);
  reg [(4'h9):(1'h0)] reg393 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg391 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg387 = (1'h0);
  reg [(5'h11):(1'h0)] forvar386 = (1'h0);
  reg [(3'h5):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar380 = (1'h0);
  reg [(4'hd):(1'h0)] reg378 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg377 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg376 = (1'h0);
  reg [(4'hb):(1'h0)] reg375 = (1'h0);
  reg [(4'hf):(1'h0)] forvar372 = (1'h0);
  reg signed [(4'he):(1'h0)] reg371 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg365 = (1'h0);
  reg [(4'h8):(1'h0)] reg361 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg360 = (1'h0);
  reg [(4'h8):(1'h0)] reg359 = (1'h0);
  reg [(4'h9):(1'h0)] reg358 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg354 = (1'h0);
  reg [(3'h4):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar352 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar351 = (1'h0);
  reg [(4'hc):(1'h0)] reg349 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg347 = (1'h0);
  reg [(2'h2):(1'h0)] forvar346 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg340 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg338 = (1'h0);
  reg [(4'hf):(1'h0)] reg337 = (1'h0);
  reg [(4'h9):(1'h0)] forvar336 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar335 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar333 = (1'h0);
  reg [(4'h8):(1'h0)] forvar318 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg331 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg326 = (1'h0);
  reg [(3'h4):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg321 = (1'h0);
  reg [(4'hb):(1'h0)] reg316 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg312 = (1'h0);
  reg [(5'h11):(1'h0)] reg308 = (1'h0);
  reg [(5'h10):(1'h0)] reg306 = (1'h0);
  reg [(4'hd):(1'h0)] forvar303 = (1'h0);
  reg [(4'h8):(1'h0)] forvar295 = (1'h0);
  reg [(3'h5):(1'h0)] reg304 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg303 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg302 = (1'h0);
  reg [(4'he):(1'h0)] forvar297 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg296 = (1'h0);
  reg [(4'hf):(1'h0)] reg295 = (1'h0);
  reg [(4'hd):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar288 = (1'h0);
  reg [(3'h6):(1'h0)] reg293 = (1'h0);
  reg [(5'h14):(1'h0)] forvar289 = (1'h0);
  reg [(5'h13):(1'h0)] reg288 = (1'h0);
  reg [(4'he):(1'h0)] reg286 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg284 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar283 = (1'h0);
  reg [(5'h11):(1'h0)] reg281 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg280 = (1'h0);
  reg [(4'ha):(1'h0)] reg279 = (1'h0);
  reg [(4'h9):(1'h0)] reg277 = (1'h0);
  reg signed [(4'he):(1'h0)] reg276 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg274 = (1'h0);
  reg [(4'ha):(1'h0)] reg272 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar271 = (1'h0);
  reg [(5'h14):(1'h0)] reg268 = (1'h0);
  reg [(5'h12):(1'h0)] reg267 = (1'h0);
  reg [(3'h5):(1'h0)] reg265 = (1'h0);
  reg [(5'h10):(1'h0)] forvar262 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg261 = (1'h0);
  reg [(5'h16):(1'h0)] reg260 = (1'h0);
  assign y = {wire614,
                 wire613,
                 wire612,
                 wire583,
                 wire542,
                 wire541,
                 wire457,
                 wire436,
                 wire435,
                 wire370,
                 wire342,
                 reg609,
                 reg607,
                 reg604,
                 reg601,
                 reg600,
                 reg598,
                 reg595,
                 reg593,
                 reg591,
                 reg590,
                 reg585,
                 reg584,
                 reg582,
                 reg579,
                 reg578,
                 reg576,
                 reg574,
                 reg573,
                 reg572,
                 reg570,
                 reg569,
                 reg567,
                 reg566,
                 reg565,
                 reg563,
                 reg562,
                 reg560,
                 reg558,
                 reg553,
                 reg544,
                 reg551,
                 reg549,
                 reg546,
                 reg545,
                 reg543,
                 reg539,
                 reg537,
                 reg536,
                 reg531,
                 reg526,
                 reg520,
                 reg529,
                 reg528,
                 reg517,
                 reg516,
                 reg514,
                 reg512,
                 reg510,
                 reg508,
                 reg504,
                 reg503,
                 reg502,
                 reg501,
                 reg500,
                 reg496,
                 reg494,
                 reg489,
                 reg485,
                 reg481,
                 reg478,
                 reg476,
                 reg472,
                 reg469,
                 reg463,
                 reg465,
                 reg461,
                 reg459,
                 reg455,
                 reg454,
                 reg452,
                 reg450,
                 reg449,
                 reg444,
                 reg441,
                 reg440,
                 reg437,
                 reg431,
                 reg433,
                 reg429,
                 reg427,
                 reg426,
                 reg423,
                 reg420,
                 reg418,
                 reg416,
                 reg415,
                 reg414,
                 reg409,
                 reg408,
                 reg406,
                 reg405,
                 reg399,
                 reg397,
                 reg392,
                 reg389,
                 reg388,
                 reg385,
                 reg384,
                 reg379,
                 reg374,
                 reg373,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg364,
                 reg363,
                 reg362,
                 reg357,
                 reg356,
                 reg355,
                 reg350,
                 reg348,
                 reg345,
                 reg344,
                 reg343,
                 reg341,
                 reg339,
                 reg334,
                 reg332,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg325,
                 reg322,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg315,
                 reg314,
                 reg313,
                 reg311,
                 reg310,
                 reg309,
                 reg307,
                 reg305,
                 reg297,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg289,
                 reg292,
                 reg291,
                 reg290,
                 reg287,
                 reg285,
                 reg282,
                 reg278,
                 reg275,
                 reg273,
                 reg270,
                 reg269,
                 reg266,
                 reg264,
                 reg263,
                 forvar605,
                 reg611,
                 reg610,
                 reg608,
                 reg606,
                 reg605,
                 reg603,
                 reg602,
                 reg599,
                 reg597,
                 reg596,
                 forvar593,
                 reg594,
                 reg592,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 forvar581,
                 reg580,
                 forvar577,
                 reg575,
                 reg571,
                 reg568,
                 forvar564,
                 reg561,
                 reg559,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 forvar552,
                 reg548,
                 reg550,
                 forvar548,
                 reg547,
                 forvar544,
                 reg540,
                 forvar538,
                 reg535,
                 reg534,
                 forvar533,
                 reg532,
                 reg530,
                 forvar516,
                 reg527,
                 forvar526,
                 reg525,
                 reg524,
                 reg523,
                 reg522,
                 reg521,
                 forvar520,
                 reg519,
                 reg518,
                 reg515,
                 forvar513,
                 reg511,
                 reg509,
                 reg507,
                 forvar506,
                 reg505,
                 reg499,
                 reg498,
                 forvar497,
                 reg495,
                 reg493,
                 forvar492,
                 reg491,
                 reg490,
                 reg488,
                 reg487,
                 forvar486,
                 reg484,
                 reg483,
                 reg482,
                 reg480,
                 reg479,
                 forvar477,
                 forvar475,
                 reg474,
                 forvar473,
                 reg471,
                 forvar470,
                 reg460,
                 reg468,
                 reg467,
                 reg466,
                 reg464,
                 forvar463,
                 reg462,
                 forvar460,
                 reg458,
                 reg456,
                 reg453,
                 reg451,
                 reg448,
                 reg447,
                 forvar446,
                 reg445,
                 reg443,
                 reg442,
                 reg439,
                 forvar438,
                 reg434,
                 reg432,
                 forvar431,
                 reg430,
                 reg428,
                 reg425,
                 reg424,
                 forvar422,
                 reg421,
                 forvar419,
                 reg417,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 forvar399,
                 reg407,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg398,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg391,
                 reg390,
                 reg387,
                 forvar386,
                 reg383,
                 reg382,
                 reg381,
                 forvar380,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 forvar372,
                 reg371,
                 reg365,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 reg354,
                 reg353,
                 forvar352,
                 forvar351,
                 reg349,
                 reg347,
                 forvar346,
                 reg340,
                 reg338,
                 reg337,
                 forvar336,
                 forvar335,
                 forvar333,
                 forvar318,
                 reg331,
                 reg326,
                 reg324,
                 reg323,
                 reg321,
                 reg316,
                 reg312,
                 reg308,
                 reg306,
                 forvar303,
                 forvar295,
                 reg304,
                 reg303,
                 reg302,
                 forvar297,
                 reg296,
                 reg295,
                 reg294,
                 forvar288,
                 reg293,
                 forvar289,
                 reg288,
                 reg286,
                 reg284,
                 forvar283,
                 reg281,
                 reg280,
                 reg279,
                 reg277,
                 reg276,
                 reg274,
                 reg272,
                 forvar271,
                 reg268,
                 reg267,
                 reg265,
                 forvar262,
                 reg261,
                 reg260,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg260 = wire258;
      reg261 = (reg260 ?
          ((wire256 & (~reg260[(4'hb):(3'h5)])) ?
              reg260[(5'h15):(5'h11)] : $signed($signed((+wire258)))) : $signed({wire258[(1'h1):(1'h1)]}));
      for (forvar262 = (1'h0); (forvar262 < (1'h0)); forvar262 = (forvar262 + (1'h1)))
        begin
          reg263 <= ((^reg260) > ($signed(reg261[(3'h4):(2'h2)]) ?
              $unsigned($signed(reg260)) : (((forvar262 <= forvar262) ?
                      reg261 : (reg260 == (7'h40))) ?
                  ($signed(wire259) + $unsigned(reg260)) : wire256)));
          if ($unsigned(($signed((~|$signed(wire256))) > $signed($signed({wire256})))))
            begin
              reg264 <= reg260[(2'h2):(1'h0)];
              reg265 = {{(~^$signed($signed(reg263)))},
                  $signed((!wire259[(3'h5):(2'h2)]))};
              reg266 <= (!reg260);
              reg267 = $signed((wire258 ?
                  $unsigned(({reg265} & (wire256 ?
                      wire258 : reg263))) : wire259[(1'h0):(1'h0)]));
              reg268 = $unsigned($signed($unsigned(reg260)));
            end
          else
            begin
              reg265 = ($signed($unsigned({(reg261 || wire259)})) ?
                  ((((reg264 ?
                          reg267 : reg261) & forvar262[(4'hd):(2'h3)]) ^ {reg260[(5'h12):(4'h8)],
                          (|(8'ha4))}) ?
                      {$unsigned($unsigned(wire259)),
                          $unsigned((!(8'haf)))} : {(+$signed(reg263)),
                          ($unsigned((8'ha2)) ?
                              reg260 : (^wire258))}) : (reg266[(3'h5):(2'h2)] + (reg268[(4'hf):(3'h6)] == $unsigned((wire257 ?
                      reg264 : reg261)))));
              reg266 <= $unsigned((~(!($unsigned(reg263) + $unsigned((8'had))))));
              reg269 <= ((($signed((~|wire259)) ?
                      reg264[(4'h8):(3'h5)] : wire256) ?
                  $signed($unsigned($unsigned(forvar262))) : (^~$unsigned((reg263 - reg260)))) <= reg267);
              reg270 <= reg269[(4'hc):(1'h0)];
            end
          for (forvar271 = (1'h0); (forvar271 < (2'h2)); forvar271 = (forvar271 + (1'h1)))
            begin
              reg272 = $signed($unsigned(wire256[(1'h0):(1'h0)]));
              reg273 <= forvar271[(4'hb):(4'ha)];
              reg274 = $unsigned(reg270[(2'h2):(1'h0)]);
              reg275 <= ($unsigned((((!reg270) ?
                  reg267[(2'h2):(1'h0)] : $unsigned(forvar271)) != $signed($unsigned(reg261)))) ^ {forvar271,
                  (~|((&reg260) ? (reg272 == reg264) : reg261))});
              reg276 = (~^$signed(reg261));
            end
          if ($unsigned($signed(reg274)))
            begin
              reg277 = $unsigned(reg264);
              reg278 <= reg261[(2'h3):(1'h0)];
              reg279 = (!$signed((wire257[(4'ha):(1'h1)] ?
                  (8'h9f) : $signed((|reg267)))));
            end
          else
            begin
              reg277 = ((~&{forvar271, {(~&reg267), reg266[(1'h0):(1'h0)]}}) ?
                  ($unsigned((reg265 != {reg261,
                      reg279})) & reg260[(5'h11):(4'hd)]) : (reg276 != ($unsigned((reg267 ?
                      (8'hae) : (8'hb7))) & $signed({(8'hbe)}))));
              reg279 = ($unsigned(reg265) >= $signed(($signed($signed((8'ha6))) ?
                  (^{reg274}) : reg261[(1'h1):(1'h1)])));
              reg280 = $unsigned((~|reg260));
              reg281 = (~&reg269[(5'h10):(5'h10)]);
              reg282 <= reg279;
            end
          for (forvar283 = (1'h0); (forvar283 < (2'h3)); forvar283 = (forvar283 + (1'h1)))
            begin
              reg284 = $unsigned(reg279);
              reg285 <= $signed((((^~$signed(forvar283)) ?
                  $signed($unsigned(reg263)) : $unsigned(((8'ha2) >>> forvar262))) - (^$unsigned((|(8'hb8))))));
              reg286 = (!(forvar262[(4'ha):(3'h6)] <<< (~|reg282)));
              reg287 <= ((^((-$unsigned(reg270)) - reg281)) ?
                  (^(7'h43)) : $unsigned($unsigned($unsigned($unsigned(reg274)))));
            end
        end
      if (reg284)
        begin
          reg288 = reg274[(1'h0):(1'h0)];
          for (forvar289 = (1'h0); (forvar289 < (1'h0)); forvar289 = (forvar289 + (1'h1)))
            begin
              reg290 <= $signed((~^$signed((reg278[(3'h6):(2'h3)] ?
                  $signed(reg278) : $unsigned(wire257)))));
              reg291 <= (wire259 <<< reg266[(3'h5):(3'h5)]);
            end
          reg292 <= {({reg284[(1'h1):(1'h1)]} ?
                  reg286 : $unsigned($signed((reg273 ? reg286 : reg281))))};
          reg293 = reg291[(5'h10):(4'hd)];
        end
      else
        begin
          for (forvar288 = (1'h0); (forvar288 < (2'h2)); forvar288 = (forvar288 + (1'h1)))
            begin
              reg289 <= $unsigned((~^(reg292[(4'h8):(1'h1)] ?
                  reg274 : (reg273 >= reg279))));
              reg290 <= (~^($unsigned($signed(reg272[(4'h8):(1'h0)])) ?
                  ((((8'ha2) ?
                      reg281 : reg287) & (forvar289 ^ reg264)) ^ (reg280[(1'h1):(1'h0)] == $signed(forvar271))) : wire259));
              reg291 <= $signed(wire257);
              reg293 = reg269[(1'h1):(1'h1)];
              reg294 = (reg270 ?
                  (~|(!$unsigned((reg278 ? (8'hb2) : reg273)))) : (&(8'hbc)));
            end
        end
      if ($unsigned($signed((reg266 || reg266[(3'h6):(3'h5)]))))
        begin
          reg295 = $signed((8'ha9));
          reg296 = $signed($signed($signed(((forvar271 ? wire256 : (7'h44)) ?
              {reg284} : $unsigned(reg284)))));
          for (forvar297 = (1'h0); (forvar297 < (3'h4)); forvar297 = (forvar297 + (1'h1)))
            begin
              reg298 <= $signed(((!forvar262[(3'h7):(3'h7)]) ?
                  $unsigned(reg290[(4'h9):(3'h7)]) : forvar283[(1'h1):(1'h1)]));
              reg299 <= reg278[(3'h6):(2'h3)];
              reg300 <= $unsigned($unsigned((reg260 > $signed($unsigned(forvar297)))));
              reg301 <= {reg276,
                  ($signed(($signed(reg272) ?
                      $signed(reg300) : (+reg279))) ^~ (7'h40))};
              reg302 = (&($unsigned(((reg299 ^~ reg277) ^~ reg300)) ?
                  reg285[(2'h3):(1'h0)] : ((~^(reg269 ?
                      reg278 : forvar271)) ^ $signed($unsigned(forvar262)))));
            end
          reg303 = (((|reg260) ?
                  reg267 : ((&reg270[(3'h4):(1'h1)]) ?
                      reg285 : $signed({wire257, reg299}))) ?
              $signed($unsigned(reg268[(3'h7):(2'h2)])) : ($unsigned(((reg296 ?
                      reg278 : (8'hbf)) ^ ((8'hb4) ~^ reg266))) ?
                  {reg299[(1'h1):(1'h0)]} : (+(8'hac))));
          reg304 = (8'hb7);
        end
      else
        begin
          for (forvar295 = (1'h0); (forvar295 < (1'h1)); forvar295 = (forvar295 + (1'h1)))
            begin
              reg297 <= $unsigned(wire259[(2'h3):(2'h2)]);
              reg298 <= $unsigned(((reg292[(5'h11):(1'h0)] ^ {(~^reg288)}) ?
                  ((^~reg270) * ((!reg279) <= (^reg300))) : (($signed(reg297) ?
                      reg261 : (forvar271 ? (8'hb2) : reg289)) || ({reg286,
                          reg287} ?
                      $unsigned(forvar283) : (reg295 <= reg279)))));
              reg299 <= reg284[(2'h3):(1'h0)];
              reg302 = (reg279[(4'h9):(3'h6)] & reg299);
            end
          for (forvar303 = (1'h0); (forvar303 < (1'h1)); forvar303 = (forvar303 + (1'h1)))
            begin
              reg305 <= $signed($unsigned($signed($signed((!forvar262)))));
              reg306 = $signed(reg288);
              reg307 <= ($unsigned(($unsigned((reg269 ? (8'h9e) : (8'hb7))) ?
                  $signed($signed(reg292)) : $unsigned((-reg284)))) || reg272[(4'h8):(3'h4)]);
              reg308 = (reg282[(3'h5):(1'h1)] ?
                  (|{reg295[(4'hd):(2'h2)],
                      reg281[(4'he):(4'h8)]}) : ($unsigned((^$unsigned(reg304))) >= $unsigned({$unsigned(reg276)})));
              reg309 <= (reg298 - ($signed(reg290) ?
                  $unsigned(reg272[(3'h4):(1'h1)]) : $signed($unsigned((reg278 ?
                      reg278 : reg278)))));
            end
          reg310 <= (forvar295 ?
              $signed(reg294[(4'hd):(2'h3)]) : (((-(&reg285)) << (reg279 ?
                      (|reg279) : {reg302, forvar303})) ?
                  {forvar283,
                      $signed((reg275 > wire259))} : (^($signed((8'had)) ?
                      $signed(wire259) : reg282[(3'h5):(2'h3)]))));
          if ((&reg299))
            begin
              reg311 <= ($unsigned((-(+{reg303}))) ?
                  (~$signed(($unsigned(reg282) > (8'h9c)))) : reg269[(3'h6):(3'h6)]);
              reg312 = (((((|forvar283) ?
                  (reg280 + reg299) : $unsigned(reg282)) | (reg287[(2'h2):(1'h1)] != wire259[(4'ha):(3'h6)])) ^~ $unsigned(reg274[(4'h9):(1'h1)])) + ((|$unsigned((reg268 ?
                  reg282 : reg266))) << (reg268[(5'h12):(4'hc)] ?
                  reg288 : reg273)));
              reg313 <= forvar295[(2'h3):(1'h0)];
              reg314 <= reg274[(2'h2):(2'h2)];
              reg315 <= (reg280 | $signed({(~&(reg290 ? reg286 : reg293)),
                  ((!forvar297) >> $signed(reg275))}));
            end
          else
            begin
              reg312 = reg293[(2'h2):(1'h1)];
              reg313 <= (reg286[(1'h1):(1'h0)] <<< (!(reg297[(3'h7):(3'h5)] ?
                  (7'h43) : $unsigned({reg272, (8'hb2)}))));
              reg314 <= $unsigned($signed({((reg300 >= wire259) ?
                      (forvar289 ? reg282 : reg268) : $signed(reg267)),
                  ($signed(forvar289) ? $signed(reg309) : (8'hb5))}));
              reg315 <= $unsigned(({((reg279 ^~ (8'hbb)) ?
                      $unsigned((7'h45)) : reg286[(4'h9):(3'h5)]),
                  ((reg269 ? reg314 : reg301) ?
                      $unsigned(reg278) : $signed(reg266))} + $signed(reg272)));
            end
        end
    end
  always
    @(posedge clk) begin
      if (wire258[(3'h5):(1'h1)])
        begin
          if ($unsigned((~&(wire258[(1'h0):(1'h0)] ?
              $signed($signed(reg298)) : (|reg300[(1'h1):(1'h0)])))))
            begin
              reg316 = reg311[(1'h0):(1'h0)];
              reg317 <= $signed(($unsigned($unsigned(((8'ha8) | reg278))) <= reg264[(3'h6):(3'h4)]));
            end
          else
            begin
              reg316 = ({reg299,
                  ({(~&(8'hab)),
                      reg311} | ((reg301 + (8'hbe)) == reg263))} << reg297[(3'h4):(3'h4)]);
              reg317 <= (reg269[(3'h5):(2'h3)] ^~ (wire258 >>> $signed({$signed(reg282),
                  (^reg292)})));
              reg318 <= ((|(-((^~(8'ha0)) >>> (reg285 ?
                  (7'h40) : reg298)))) <= $unsigned((((reg315 ?
                  reg287 : reg309) || (reg301 ? reg273 : reg305)) ~^ (((7'h48) ?
                  reg317 : reg313) > $signed((7'h42))))));
              reg319 <= ($unsigned(($unsigned(reg298) ~^ reg266[(2'h3):(1'h1)])) << $unsigned(reg269));
              reg320 <= reg266[(2'h3):(2'h3)];
            end
          if ((({(reg299 >= (reg317 ?
                      reg298 : reg299))} >= {$unsigned(reg275)}) ?
              $signed(((-(-(8'ha5))) ?
                  (~(reg285 == reg317)) : $unsigned($unsigned(reg320)))) : $unsigned((!reg310[(3'h5):(3'h5)]))))
            begin
              reg321 = reg291;
              reg322 <= $unsigned(reg263);
            end
          else
            begin
              reg321 = (($unsigned(reg290[(3'h4):(1'h1)]) - {reg285,
                  ($unsigned(reg311) || (reg316 ?
                      reg307 : reg300))}) >= $unsigned(reg315[(2'h3):(2'h2)]));
              reg323 = reg311[(3'h6):(1'h1)];
            end
          reg324 = $unsigned($signed((8'h9f)));
          reg325 <= $unsigned($signed((($signed(reg318) & reg275) >> reg315[(2'h3):(2'h3)])));
          if ({{(~&reg319), reg298[(3'h5):(3'h5)]},
              ((wire258[(3'h4):(1'h0)] ?
                  reg290[(4'hd):(3'h5)] : $signed(reg287)) * reg292[(1'h1):(1'h0)])})
            begin
              reg326 = {(&$signed($signed(reg323)))};
            end
          else
            begin
              reg327 <= $signed(($unsigned($unsigned($signed(reg323))) ?
                  reg318[(1'h1):(1'h1)] : wire257[(1'h0):(1'h0)]));
              reg328 <= ($unsigned(reg315) + $unsigned($unsigned({$unsigned(reg323)})));
              reg329 <= {(&(reg321 || reg313))};
              reg330 <= ({reg297[(2'h3):(2'h2)]} ?
                  $unsigned((^~reg264)) : ({reg287[(1'h0):(1'h0)], (8'h9d)} ?
                      ((reg310[(3'h7):(1'h0)] ?
                          ((8'ha2) <= wire259) : (reg275 ?
                              reg324 : reg324)) - {(reg297 < (7'h46))}) : reg305));
              reg331 = ((!$unsigned($signed((reg322 - reg273)))) || (8'hbc));
            end
        end
      else
        begin
          reg317 <= wire259[(4'he):(4'hc)];
          for (forvar318 = (1'h0); (forvar318 < (2'h2)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg319 <= reg320[(1'h1):(1'h1)];
              reg320 <= reg275;
            end
          if (((~^reg330) ?
              forvar318 : (|(reg320 ?
                  reg324 : $unsigned(reg292[(3'h6):(2'h2)])))))
            begin
              reg322 <= ((7'h43) ?
                  (($signed((reg292 == reg297)) - reg282) ?
                      reg278 : ((~&(reg309 >= reg282)) >= reg320)) : ((+((|reg324) ?
                          (8'hbc) : (reg289 ? reg324 : (8'hb3)))) ?
                      ((~$unsigned(reg263)) * reg310[(2'h3):(1'h1)]) : (|reg299)));
              reg323 = ($signed(reg309) ?
                  $signed(reg323[(4'he):(4'he)]) : reg270[(1'h0):(1'h0)]);
              reg325 <= ($signed({$unsigned((reg325 ? reg270 : reg328))}) ?
                  $signed(($unsigned($unsigned(reg318)) ?
                      (reg313[(3'h7):(2'h2)] ?
                          $unsigned(reg327) : ((8'haf) ?
                              reg273 : reg331)) : (reg326 == $signed((8'hb3))))) : reg314);
              reg327 <= $unsigned(reg317[(4'hd):(1'h1)]);
            end
          else
            begin
              reg322 <= $signed(reg314[(3'h6):(3'h6)]);
              reg323 = (reg318 ?
                  (reg314[(3'h4):(1'h0)] ?
                      $signed((^(-reg310))) : (8'ha2)) : $signed((&(forvar318 ?
                      (~reg311) : (reg311 ? reg301 : wire257)))));
              reg325 <= (reg285 >= (~&{((&reg263) ?
                      (^reg326) : wire256[(2'h3):(1'h0)])}));
              reg327 <= {$unsigned(($unsigned((reg291 ? reg273 : reg305)) ?
                      $unsigned((~|(7'h46))) : ({reg270, reg309} ?
                          reg315[(3'h5):(3'h4)] : (!reg317))))};
            end
        end
      reg332 <= (~|reg325[(3'h6):(1'h1)]);
      for (forvar333 = (1'h0); (forvar333 < (1'h1)); forvar333 = (forvar333 + (1'h1)))
        begin
          reg334 <= (8'hb1);
        end
      for (forvar335 = (1'h0); (forvar335 < (1'h0)); forvar335 = (forvar335 + (1'h1)))
        begin
          for (forvar336 = (1'h0); (forvar336 < (2'h2)); forvar336 = (forvar336 + (1'h1)))
            begin
              reg337 = $unsigned((^reg315[(4'h8):(3'h5)]));
              reg338 = $unsigned($signed($unsigned($unsigned(reg334))));
              reg339 <= (~&(reg269[(4'hf):(4'ha)] & $signed($signed($unsigned(reg309)))));
              reg340 = $unsigned((^reg314));
            end
          reg341 <= $unsigned({{$signed((|wire258))}, $signed(forvar318)});
        end
    end
  assign wire342 = reg275;
  always
    @(posedge clk) begin
      if ($unsigned(reg285))
        begin
          reg343 <= ($unsigned($signed(({reg299} != $unsigned(reg291)))) ?
              reg310 : $unsigned($unsigned(($signed((8'h9f)) <= (8'hab)))));
          reg344 <= (reg320[(4'hf):(1'h0)] >= $unsigned(($signed((reg266 ?
                  reg273 : wire257)) ?
              {reg305[(2'h2):(1'h0)], (~&wire258)} : (~&$unsigned(reg317)))));
          reg345 <= (^$signed($unsigned((+$unsigned((8'hb8))))));
          for (forvar346 = (1'h0); (forvar346 < (1'h1)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 = reg314[(3'h5):(2'h2)];
              reg348 <= (~|(^{(((8'hb5) ?
                      reg305 : reg264) >>> $signed(reg328))}));
              reg349 = reg305[(4'he):(2'h3)];
              reg350 <= (-$signed($unsigned(((+reg275) & reg322[(4'hb):(3'h6)]))));
            end
        end
      else
        begin
          reg343 <= (reg350[(4'h9):(3'h6)] << (~|reg314));
          reg344 <= reg290[(2'h3):(1'h0)];
        end
      for (forvar351 = (1'h0); (forvar351 < (1'h0)); forvar351 = (forvar351 + (1'h1)))
        begin
          for (forvar352 = (1'h0); (forvar352 < (1'h1)); forvar352 = (forvar352 + (1'h1)))
            begin
              reg353 = reg343[(1'h0):(1'h0)];
              reg354 = (|({$unsigned((|(8'ha3))),
                  ((!reg264) ?
                      $signed(reg270) : (forvar346 ?
                          reg328 : reg300))} > (reg300[(1'h0):(1'h0)] & ($unsigned(reg310) ?
                  $unsigned(reg345) : (reg287 ? (8'hb9) : reg278)))));
              reg355 <= $unsigned(reg354[(1'h1):(1'h0)]);
              reg356 <= (^~wire342[(4'hc):(2'h3)]);
              reg357 <= reg341[(4'h8):(3'h6)];
            end
          reg358 = $unsigned(reg356);
          if ($signed(wire257[(4'ha):(2'h2)]))
            begin
              reg359 = reg270;
              reg360 = {(^~$unsigned({$unsigned(reg343), (reg334 || reg297)}))};
              reg361 = $unsigned({$unsigned(((~|reg327) ?
                      (-reg291) : reg347[(5'h16):(5'h14)])),
                  (&(8'hbb))});
              reg362 <= $signed(reg357[(4'hc):(1'h0)]);
              reg363 <= (reg341 > reg325[(3'h4):(1'h1)]);
            end
          else
            begin
              reg359 = (~&(!({reg270[(2'h3):(1'h1)], (&reg348)} ?
                  ($signed(reg332) <<< {reg344}) : reg266)));
            end
          reg364 <= reg314[(2'h3):(2'h3)];
          if ((~$unsigned((~^(!{(7'h46), reg313})))))
            begin
              reg365 = ($signed($signed(($signed(reg270) ?
                      (reg270 ? reg263 : reg349) : wire257))) ?
                  ($signed(reg327) ?
                      (reg270[(3'h4):(1'h1)] ?
                          ($signed(reg345) ?
                              (reg315 < reg322) : reg285) : (!(wire342 ?
                              reg354 : reg356))) : (8'ha6)) : {$unsigned(({reg361} << (^~(7'h42)))),
                      ((reg289[(3'h5):(2'h2)] != reg329[(3'h4):(3'h4)]) != $unsigned(((7'h47) ?
                          (8'h9c) : reg330)))});
              reg366 <= ({$signed((-{(8'hbb)}))} ?
                  $signed((!$unsigned(reg329))) : reg325);
              reg367 <= (+($signed(reg325) | {($unsigned((8'h9e)) ?
                      (forvar352 == reg348) : reg282[(3'h4):(1'h0)])}));
              reg368 <= $unsigned(($signed((^~((8'ha0) ?
                  reg339 : wire259))) + (^($unsigned(reg353) ?
                  (8'ha3) : $unsigned(reg270)))));
              reg369 <= $unsigned({wire258});
            end
          else
            begin
              reg366 <= (reg348 - $unsigned(($signed(wire259[(4'hc):(2'h2)]) ?
                  $signed((reg349 ? reg366 : reg362)) : reg311)));
              reg367 <= (~$signed(($signed(reg361) >>> {reg358[(3'h4):(3'h4)]})));
            end
        end
    end
  assign wire370 = (reg264 - (^(+({reg319} ?
                       $signed((8'haa)) : reg310[(3'h5):(3'h4)]))));
  always
    @(posedge clk) begin
      reg371 = ((($signed($signed(reg273)) <<< ($signed(reg369) || (reg300 ?
              reg313 : reg328))) != $signed({(reg297 ? reg289 : reg314),
              (reg327 >>> (7'h48))})) ?
          reg363[(2'h2):(2'h2)] : reg275);
      for (forvar372 = (1'h0); (forvar372 < (1'h1)); forvar372 = (forvar372 + (1'h1)))
        begin
          reg373 <= (wire257[(1'h0):(1'h0)] ?
              $signed(reg290[(5'h11):(3'h6)]) : reg355[(1'h0):(1'h0)]);
          reg374 <= reg311;
          if (reg264)
            begin
              reg375 = ((^~(~&{reg368[(1'h1):(1'h0)], $unsigned((8'hb0))})) ?
                  ($unsigned(((reg278 ^ reg343) == (reg290 ?
                      wire342 : wire259))) * {reg270[(2'h3):(1'h0)],
                      $unsigned(reg266[(2'h3):(1'h1)])}) : $unsigned(reg343[(1'h0):(1'h0)]));
              reg376 = (^reg285);
              reg377 = (((~reg313) ?
                  (~^reg266) : (reg357 >> (8'hae))) != wire259);
              reg378 = ($signed(({((8'h9c) ? reg285 : (8'ha5))} + (~^(reg345 ?
                  reg275 : wire258)))) <<< reg373);
            end
          else
            begin
              reg375 = (^~$signed(reg373[(3'h4):(2'h3)]));
              reg376 = reg292;
              reg379 <= $signed(reg307[(3'h6):(3'h6)]);
            end
          for (forvar380 = (1'h0); (forvar380 < (2'h2)); forvar380 = (forvar380 + (1'h1)))
            begin
              reg381 = ($unsigned($signed(reg317)) ?
                  $signed((~&$signed((reg357 ~^ wire256)))) : (((~^reg317[(5'h12):(5'h12)]) ?
                      ($unsigned(reg299) ?
                          $signed(reg285) : (~wire256)) : $signed((reg377 && (8'haa)))) - (reg362 <<< reg364[(3'h7):(2'h3)])));
              reg382 = reg273[(2'h3):(2'h2)];
              reg383 = reg332;
              reg384 <= ($unsigned((reg377[(1'h0):(1'h0)] ?
                  ($signed((7'h48)) ?
                      {(7'h48),
                          wire259} : (reg319 ^~ reg270)) : reg298)) || (^~($signed(((7'h44) ?
                  reg327 : (8'hae))) - reg362)));
              reg385 <= (reg317[(3'h4):(1'h1)] + reg310);
            end
        end
      if (reg332[(4'he):(3'h7)])
        begin
          for (forvar386 = (1'h0); (forvar386 < (1'h0)); forvar386 = (forvar386 + (1'h1)))
            begin
              reg387 = $unsigned($unsigned($unsigned($unsigned((^reg367)))));
              reg388 <= $unsigned((~|reg343[(3'h4):(1'h0)]));
            end
          reg389 <= (+{$signed($unsigned((wire258 > reg305))),
              (-$unsigned(((8'hbc) ? wire342 : reg301)))});
          reg390 = $unsigned(($unsigned((-reg348)) + (reg319[(2'h3):(2'h3)] <= reg264[(1'h0):(1'h0)])));
          if ((!$signed(({$unsigned(reg329)} ?
              reg369[(4'hc):(3'h5)] : reg343[(3'h5):(3'h5)]))))
            begin
              reg391 = reg344[(3'h5):(1'h0)];
              reg392 <= reg319;
              reg393 = ($unsigned(reg379) ?
                  (8'hae) : (reg300[(1'h1):(1'h1)] < $unsigned(reg357[(5'h10):(3'h6)])));
            end
          else
            begin
              reg392 <= $signed(reg373);
              reg393 = ($signed($signed((((8'ha5) ^ reg377) > $signed((7'h40))))) ?
                  ((reg385[(3'h4):(2'h2)] ?
                      ($signed(reg327) ?
                          ((8'hbb) ?
                              reg369 : reg310) : $unsigned((8'ha7))) : (!$unsigned(reg341))) & reg270[(2'h3):(2'h3)]) : ($signed(reg301) < $unsigned($signed($unsigned(reg373)))));
              reg394 = {$unsigned($unsigned(reg299[(1'h0):(1'h0)])),
                  $unsigned($unsigned($signed((+reg290))))};
              reg395 = reg381[(1'h1):(1'h1)];
              reg396 = (wire257[(3'h4):(2'h2)] - (forvar386[(4'he):(4'ha)] >>> $signed(reg387[(4'hd):(3'h6)])));
            end
        end
      else
        begin
          for (forvar386 = (1'h0); (forvar386 < (2'h2)); forvar386 = (forvar386 + (1'h1)))
            begin
              reg388 <= (((~reg385) * reg332) ?
                  reg364[(3'h7):(3'h4)] : (~^reg317[(4'he):(1'h0)]));
              reg389 <= reg389[(2'h2):(1'h1)];
              reg392 <= $unsigned($signed(reg344[(2'h2):(1'h0)]));
              reg393 = $signed((!reg318));
            end
          reg394 = (+wire256);
          reg397 <= reg367[(2'h3):(1'h1)];
          reg398 = {$unsigned(($unsigned(reg348[(4'he):(2'h3)]) ?
                  reg379[(3'h4):(2'h3)] : (reg339[(1'h0):(1'h0)] > (+reg301)))),
              reg385};
        end
      if ({($unsigned((-(reg322 & reg355))) & (({reg394} ?
                  reg297[(2'h3):(1'h0)] : reg275[(3'h5):(2'h3)]) ?
              (~reg301[(1'h1):(1'h1)]) : reg389[(1'h1):(1'h0)])),
          reg379})
        begin
          reg399 <= $signed($unsigned((reg322 & reg385[(3'h4):(2'h3)])));
          if (reg379)
            begin
              reg400 = reg314[(4'hd):(4'hb)];
              reg401 = reg356;
              reg402 = (8'hbe);
              reg403 = (((reg379[(2'h2):(1'h0)] + reg389[(1'h0):(1'h0)]) >> $unsigned($unsigned(reg334))) ?
                  $unsigned($signed(((wire370 ? wire342 : reg348) ?
                      (forvar380 >= reg287) : {reg270,
                          reg327}))) : ((!reg348) ~^ $unsigned({$signed(reg314),
                      {reg383}})));
              reg404 = $signed(((($signed(reg398) ?
                          (reg298 ? wire256 : reg397) : {reg318, reg385}) ?
                      reg387[(4'he):(1'h1)] : (reg328[(5'h10):(4'he)] ?
                          $signed(reg355) : (8'hb2))) ?
                  $unsigned(reg273) : ($unsigned(((8'hb7) ?
                      reg356 : reg390)) || (~|reg322))));
            end
          else
            begin
              reg405 <= $unsigned(reg390);
              reg406 <= (~^reg329);
              reg407 = reg356;
              reg408 <= (reg315 ?
                  (reg311[(4'hc):(4'ha)] & reg345) : reg406[(3'h6):(1'h1)]);
              reg409 <= reg388[(1'h1):(1'h1)];
            end
        end
      else
        begin
          for (forvar399 = (1'h0); (forvar399 < (1'h0)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg405 <= $signed((!(reg311 ^ ((reg298 ?
                  wire256 : reg397) + (reg403 ? reg404 : reg367)))));
            end
          reg407 = ($unsigned($unsigned($unsigned((reg391 & (8'h9d))))) ?
              $unsigned(reg292) : reg318);
        end
    end
  always
    @(posedge clk) begin
      reg410 = ((wire258 ?
          {($signed((8'hb2)) ? (reg374 ? reg318 : (7'h45)) : $unsigned(reg379)),
              reg379} : {($signed((8'hb6)) ?
                  (reg299 ? wire370 : reg339) : reg305),
              reg357[(3'h5):(3'h4)]}) || {(^$signed(reg311))});
      if ((&$signed(reg273[(3'h5):(1'h1)])))
        begin
          reg411 = {((($unsigned(reg366) ?
                  (reg410 + (7'h43)) : (reg392 <<< reg363)) & $signed(wire256)) * (((reg334 ?
                      reg397 : reg368) ^~ (reg408 ? reg325 : reg291)) ?
                  ((reg364 ? reg275 : (7'h48)) ?
                      (reg266 ?
                          reg348 : (8'hae)) : $signed(reg345)) : $unsigned(((8'hb8) ?
                      (8'ha7) : reg317)))),
              (8'hbb)};
          if ({reg363})
            begin
              reg412 = {$signed(reg269[(4'hc):(3'h7)]), reg317[(4'hb):(4'ha)]};
              reg413 = $signed($signed($unsigned((|$signed((7'h47))))));
              reg414 <= $signed((((&reg269) ~^ (8'hbe)) ?
                  (reg364[(4'h8):(4'h8)] < $unsigned($unsigned((7'h41)))) : (reg270[(3'h4):(1'h1)] ?
                      (reg384[(4'he):(4'hc)] ?
                          $signed((7'h45)) : ((8'ha1) || reg292)) : wire342)));
              reg415 <= reg318[(2'h3):(2'h2)];
              reg416 <= $unsigned((^~(~&$signed((wire370 ?
                  reg367 : (8'hb0))))));
            end
          else
            begin
              reg412 = reg309;
              reg414 <= ((+((&$signed((8'hb8))) | (8'hba))) ?
                  (({(reg292 + reg416)} & reg392[(2'h3):(1'h1)]) - ($unsigned($unsigned((8'h9c))) ?
                      ((reg291 | reg343) == (reg356 ?
                          reg297 : reg305)) : ((^reg285) ?
                          (reg290 ? reg287 : reg319) : (reg319 ?
                              reg373 : reg327)))) : $signed(reg270));
            end
        end
      else
        begin
          if ($unsigned((|$signed((reg273[(3'h4):(1'h1)] * {reg314})))))
            begin
              reg411 = ($signed({reg348,
                  $unsigned($signed(reg414))}) ^~ ((($unsigned(reg301) ?
                      reg317 : $unsigned(reg416)) ?
                  ($signed(reg362) ?
                      (reg289 ?
                          reg320 : reg385) : (reg327 ~^ reg315)) : $unsigned((reg362 << reg392))) < $signed(((reg318 > reg414) ?
                  wire256[(1'h1):(1'h0)] : $unsigned(reg314)))));
              reg414 <= reg413[(4'hd):(3'h7)];
              reg417 = reg285[(4'he):(4'hc)];
            end
          else
            begin
              reg411 = $signed((wire259 ?
                  $signed(reg300) : $unsigned(($signed(reg417) ?
                      reg348 : $signed(reg289)))));
              reg412 = (8'h9d);
              reg414 <= (&((wire257[(2'h3):(1'h1)] ?
                      $signed($unsigned(reg332)) : (reg320[(5'h10):(4'he)] & (reg332 & (8'hb9)))) ?
                  $signed({(~^reg332)}) : $signed(({reg414} ?
                      $signed(reg309) : $signed(reg299)))));
              reg417 = {reg285[(4'h8):(3'h5)]};
              reg418 <= $unsigned(($unsigned(($signed(reg289) ?
                  (~reg392) : $unsigned((7'h42)))) & reg373));
            end
        end
      for (forvar419 = (1'h0); (forvar419 < (2'h2)); forvar419 = (forvar419 + (1'h1)))
        begin
          reg420 <= $signed({$signed((8'hb1)), wire342});
          reg421 = $unsigned(({((reg297 && wire259) ? (~(8'hb2)) : (~reg315))} ?
              reg410 : reg290));
          for (forvar422 = (1'h0); (forvar422 < (1'h1)); forvar422 = (forvar422 + (1'h1)))
            begin
              reg423 <= $signed((reg415 ?
                  reg389[(2'h2):(1'h0)] : (($signed(reg325) ?
                          (^wire342) : reg301) ?
                      $unsigned(reg384) : reg318[(1'h1):(1'h0)])));
              reg424 = reg412[(5'h11):(3'h5)];
              reg425 = reg299[(1'h0):(1'h0)];
              reg426 <= $unsigned((reg412[(4'ha):(4'ha)] ?
                  $signed((reg291 <= ((8'hbd) << (8'hb5)))) : $signed($unsigned($unsigned((8'hac))))));
            end
          reg427 <= reg423;
        end
      if ((~(($unsigned((reg322 >= reg385)) ?
              $signed($signed(reg285)) : (~^$signed(reg314))) ?
          (~|$signed($unsigned(reg264))) : reg330)))
        begin
          reg428 = {$signed(($unsigned((~&reg270)) >>> reg263))};
        end
      else
        begin
          reg429 <= {(reg408[(1'h0):(1'h0)] | reg329)};
        end
      if ((^$unsigned((~{reg341[(2'h2):(1'h0)], reg322}))))
        begin
          reg430 = $unsigned($unsigned((reg429[(2'h2):(1'h1)] ~^ reg311[(4'hc):(1'h0)])));
          for (forvar431 = (1'h0); (forvar431 < (1'h0)); forvar431 = (forvar431 + (1'h1)))
            begin
              reg432 = (reg416[(2'h2):(1'h1)] ?
                  $unsigned((~^reg344)) : (wire342 ?
                      $unsigned(reg410) : $signed(((reg311 ? reg341 : reg355) ?
                          (reg298 ? reg345 : reg282) : (reg334 ?
                              reg348 : (7'h42))))));
            end
          reg433 <= ((reg388[(1'h1):(1'h1)] ?
                  reg314[(4'h8):(1'h1)] : $unsigned((8'hb6))) ?
              reg388[(3'h5):(1'h0)] : (({$signed(reg412),
                  (-wire370)} >> ((8'ha6) <= {reg423, (8'ha7)})) || (~reg409)));
        end
      else
        begin
          reg431 <= (reg412[(4'he):(1'h1)] ?
              {(reg313[(3'h4):(1'h0)] ?
                      $signed((reg421 & reg317)) : reg415[(2'h3):(1'h0)])} : {$signed(reg405)});
          reg432 = $signed($signed($unsigned($unsigned((reg325 ^~ reg364)))));
          reg434 = (^reg428[(5'h10):(2'h3)]);
        end
    end
  assign wire435 = $signed(reg322);
  assign wire436 = reg282;
  always
    @(posedge clk) begin
      reg437 <= reg384;
      for (forvar438 = (1'h0); (forvar438 < (1'h0)); forvar438 = (forvar438 + (1'h1)))
        begin
          if (reg356[(3'h6):(3'h4)])
            begin
              reg439 = reg319[(3'h4):(2'h3)];
              reg440 <= $unsigned($signed((~^$signed({reg345}))));
              reg441 <= reg300[(2'h2):(1'h1)];
            end
          else
            begin
              reg439 = (+reg343[(4'h8):(3'h7)]);
              reg442 = reg285[(2'h2):(2'h2)];
              reg443 = ($signed($signed(reg364[(1'h1):(1'h0)])) <= (8'ha7));
            end
          reg444 <= ($unsigned($signed(($signed(reg416) <<< ((8'h9e) <<< reg332)))) ^~ $signed((reg291 ?
              reg285[(2'h2):(1'h0)] : (+(-reg418)))));
          reg445 = {$unsigned(reg317),
              ((reg388[(2'h2):(2'h2)] ?
                  $signed((reg343 ?
                      reg368 : reg406)) : (8'hbe)) < $signed($signed((reg366 ?
                  (8'hb7) : reg341))))};
          for (forvar446 = (1'h0); (forvar446 < (1'h0)); forvar446 = (forvar446 + (1'h1)))
            begin
              reg447 = (~$unsigned($signed(((^~reg345) ?
                  ((8'hb3) & (8'hb6)) : (reg273 <= reg443)))));
              reg448 = ((((reg433[(1'h1):(1'h1)] ?
                          reg431[(2'h2):(2'h2)] : reg320[(3'h6):(2'h2)]) ?
                      ($signed(reg420) ?
                          (reg322 ? reg327 : reg322) : {reg431,
                              reg300}) : reg373[(4'hd):(4'hb)]) & $unsigned(($signed((8'haa)) ?
                      reg344 : $signed(reg427)))) ?
                  (((&(^~(8'hab))) ?
                      reg307 : ($unsigned(reg416) | (!reg364))) << $unsigned(((7'h41) | $signed(reg299)))) : ((8'ha5) <= (|$signed(reg373[(1'h1):(1'h1)]))));
              reg449 <= reg366[(2'h2):(2'h2)];
              reg450 <= reg325[(3'h7):(1'h1)];
            end
          if (((|$unsigned((~$signed(reg385)))) ^ reg339[(4'h8):(3'h4)]))
            begin
              reg451 = ($unsigned((((reg392 >= reg309) ?
                      (reg433 ?
                          reg388 : reg405) : (reg414 < reg437)) - ($unsigned(reg285) ?
                      {reg427} : reg440))) ?
                  $unsigned(reg299[(1'h0):(1'h0)]) : (reg389[(1'h1):(1'h1)] & $signed($unsigned($signed(reg290)))));
              reg452 <= reg368;
              reg453 = $signed(reg329[(5'h16):(5'h16)]);
            end
          else
            begin
              reg451 = reg364;
              reg453 = $signed(reg313);
              reg454 <= (~(~&reg451[(4'h9):(4'h9)]));
              reg455 <= (~^(|(~|((reg330 < (8'had)) ?
                  (wire256 > reg297) : reg350))));
              reg456 = (8'ha8);
            end
        end
    end
  assign wire457 = $unsigned((($signed((reg313 ^~ reg289)) ~^ $signed((reg278 ?
                       reg287 : reg415))) ^ $unsigned((reg355[(2'h2):(2'h2)] & reg363))));
  always
    @(posedge clk) begin
      reg458 = $signed(reg373[(3'h5):(1'h1)]);
      if ((&wire370))
        begin
          reg459 <= reg416[(2'h3):(2'h3)];
          for (forvar460 = (1'h0); (forvar460 < (1'h0)); forvar460 = (forvar460 + (1'h1)))
            begin
              reg461 <= $signed($signed($signed(($unsigned(reg423) ?
                  $unsigned((8'hb9)) : {reg356, reg350}))));
            end
          reg462 = reg313;
          for (forvar463 = (1'h0); (forvar463 < (2'h3)); forvar463 = (forvar463 + (1'h1)))
            begin
              reg464 = reg367[(4'h9):(3'h7)];
              reg465 <= reg429[(2'h3):(1'h1)];
              reg466 = ((^{$unsigned(reg364[(4'h8):(2'h3)]), reg341}) ?
                  reg431 : {$signed((8'hb5)),
                      (reg317[(3'h4):(1'h1)] ?
                          (reg305 > $signed(reg348)) : (+reg379[(4'h9):(4'h9)]))});
              reg467 = reg462;
              reg468 = ((-{({reg431, reg392} & ((8'h9e) ^ reg348)),
                      $signed($signed((8'hb4)))}) ?
                  {(reg389[(2'h2):(1'h1)] ?
                          $unsigned($signed(reg325)) : wire457),
                      ((reg449 <= reg431) ?
                          $signed(reg315) : $unsigned(reg282[(2'h2):(1'h0)]))} : $unsigned($signed(wire457[(1'h1):(1'h1)])));
            end
        end
      else
        begin
          reg460 = reg452[(2'h2):(1'h1)];
          if (reg301[(4'h8):(3'h6)])
            begin
              reg461 <= (~^$signed(reg329[(4'hc):(2'h2)]));
              reg462 = (^~((^~(~^(reg339 < reg367))) * (|(^~(reg273 >>> wire259)))));
            end
          else
            begin
              reg461 <= $signed(((reg285 ?
                      ((8'hb9) ?
                          reg455 : reg369[(5'h10):(3'h6)]) : reg275[(3'h4):(3'h4)]) ?
                  reg467[(4'he):(4'h9)] : $signed($signed((reg310 ?
                      reg314 : reg392)))));
              reg463 <= reg345[(3'h4):(1'h0)];
              reg465 <= reg325[(1'h0):(1'h0)];
              reg469 <= reg334[(3'h5):(2'h2)];
            end
          for (forvar470 = (1'h0); (forvar470 < (2'h3)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 = ((((8'haf) ?
                  reg322[(3'h7):(3'h5)] : $signed($signed(reg374))) >= $unsigned((reg322[(5'h10):(3'h5)] + (reg367 ^ reg374)))) >= reg273[(4'ha):(3'h7)]);
            end
        end
      reg472 <= reg469[(4'hc):(3'h4)];
      for (forvar473 = (1'h0); (forvar473 < (3'h4)); forvar473 = (forvar473 + (1'h1)))
        begin
          reg474 = forvar473;
          for (forvar475 = (1'h0); (forvar475 < (2'h2)); forvar475 = (forvar475 + (1'h1)))
            begin
              reg476 <= reg465[(2'h2):(1'h0)];
            end
          for (forvar477 = (1'h0); (forvar477 < (2'h2)); forvar477 = (forvar477 + (1'h1)))
            begin
              reg478 <= (reg307 ?
                  ((reg409 * ((+reg472) ?
                          ((8'hb2) ? reg317 : (8'ha0)) : $unsigned(reg270))) ?
                      reg325[(1'h1):(1'h0)] : (~(~|$signed((8'hb7))))) : (&(-$signed(((7'h45) & reg317)))));
              reg479 = (~{($unsigned(reg357) & $unsigned(reg474[(4'h9):(3'h7)]))});
              reg480 = ((~|({(^reg314), $unsigned(reg273)} ?
                  (^~reg418[(2'h3):(2'h3)]) : (reg464 >>> (&reg420)))) >>> $unsigned($signed((reg356 ?
                  (reg467 ? (7'h48) : (7'h42)) : (~|reg356)))));
            end
          if ((|forvar475[(2'h3):(1'h1)]))
            begin
              reg481 <= (~&wire257[(4'hb):(3'h4)]);
              reg482 = ((8'hae) != wire258[(2'h2):(1'h1)]);
              reg483 = {$signed($unsigned($unsigned($unsigned(reg343))))};
              reg484 = $signed($signed(reg399[(4'hc):(4'hc)]));
              reg485 <= $signed((8'hb9));
            end
          else
            begin
              reg482 = (8'hb4);
              reg483 = ((((reg384 - (8'hae)) > (~^reg356[(4'ha):(1'h1)])) & $unsigned(reg384)) ?
                  reg478 : (({{reg367},
                      $signed(reg463)} || (~$signed(reg299))) & (!(8'hba))));
              reg484 = ((~^reg416[(3'h5):(3'h5)]) ?
                  reg350 : ($unsigned((^~((8'ha7) ? reg313 : reg325))) ?
                      reg362 : ($signed($unsigned(reg273)) | reg330[(3'h4):(1'h0)])));
              reg485 <= (&$signed($signed(((&(8'hb7)) ?
                  reg455[(4'hd):(4'ha)] : reg310))));
            end
        end
      for (forvar486 = (1'h0); (forvar486 < (1'h1)); forvar486 = (forvar486 + (1'h1)))
        begin
          if (reg467)
            begin
              reg487 = reg325[(3'h5):(2'h2)];
            end
          else
            begin
              reg487 = (($unsigned($signed(((8'haa) <<< wire257))) <<< ($signed(wire259[(5'h14):(3'h5)]) & (7'h47))) ?
                  $signed(reg433) : reg420);
              reg488 = reg460;
              reg489 <= (~((-reg485[(4'hd):(1'h1)]) ?
                  $unsigned(wire435) : wire370[(2'h3):(1'h0)]));
              reg490 = reg397[(4'hc):(4'hc)];
              reg491 = ((reg478 ? reg291 : {reg478}) ?
                  $unsigned(forvar477[(2'h2):(1'h0)]) : reg471);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar492 = (1'h0); (forvar492 < (1'h0)); forvar492 = (forvar492 + (1'h1)))
        begin
          if ((-(+(~^wire258[(3'h5):(1'h0)]))))
            begin
              reg493 = (reg264[(1'h1):(1'h1)] ?
                  (~|{forvar492[(3'h5):(3'h4)]}) : {((8'hb9) * (~|$signed(reg332)))});
              reg494 <= reg328;
              reg495 = reg455;
            end
          else
            begin
              reg494 <= (~(~^$signed({reg287[(1'h1):(1'h0)]})));
              reg495 = ($unsigned($unsigned((8'ha1))) >> (^~(reg379 && reg374)));
              reg496 <= (8'hbf);
            end
          for (forvar497 = (1'h0); (forvar497 < (3'h4)); forvar497 = (forvar497 + (1'h1)))
            begin
              reg498 = reg297;
              reg499 = reg270;
              reg500 <= (~(^~(8'haa)));
            end
          reg501 <= $signed(reg440);
          reg502 <= {reg431[(2'h2):(1'h1)],
              ((reg290[(5'h12):(4'hd)] ?
                  (7'h41) : ((reg263 ? reg493 : reg499) * (7'h43))) + reg472)};
          reg503 <= ($signed($unsigned(reg373[(3'h7):(3'h4)])) ?
              ((7'h45) - (^(reg499[(4'h9):(3'h5)] ?
                  ((8'ha2) ?
                      reg314 : wire457) : ((7'h46) | reg472)))) : {$unsigned((reg287[(1'h0):(1'h0)] ?
                      (reg452 ? reg493 : reg330) : reg379))});
        end
    end
  always
    @(posedge clk) begin
      reg504 <= $unsigned($unsigned((reg292 ?
          $unsigned((^~reg264)) : ($unsigned(reg264) ~^ $unsigned((8'had))))));
      reg505 = (~|(reg270 < {$signed((-reg300)),
          ({wire436, reg418} == (!reg329))}));
      for (forvar506 = (1'h0); (forvar506 < (1'h0)); forvar506 = (forvar506 + (1'h1)))
        begin
          if (($signed((^reg309[(3'h6):(1'h0)])) > ({(+$signed(reg269)),
              ((^~(8'hbd)) ~^ (7'h48))} + reg478)))
            begin
              reg507 = {reg389};
              reg508 <= (8'ha8);
              reg509 = {(8'haa)};
              reg510 <= ($unsigned(((wire435[(1'h1):(1'h0)] >= $unsigned(reg374)) ?
                  $signed((reg508 && reg469)) : reg322[(2'h2):(1'h1)])) - reg290[(5'h12):(5'h10)]);
              reg511 = $unsigned(reg431);
            end
          else
            begin
              reg508 <= {reg423[(5'h14):(1'h1)]};
            end
          reg512 <= ((~|$signed((reg469[(5'h13):(3'h7)] ?
                  {reg489} : (8'hbe)))) ?
              reg399 : reg463);
          for (forvar513 = (1'h0); (forvar513 < (2'h2)); forvar513 = (forvar513 + (1'h1)))
            begin
              reg514 <= reg384;
            end
        end
      reg515 = ((reg373 ? {(-(^(8'hb4)))} : (reg504 ^~ {{(8'h9e), reg489}})) ?
          $unsigned($unsigned($unsigned($signed(reg504)))) : reg388);
      if (reg320[(4'h9):(4'h8)])
        begin
          if ({$unsigned(($unsigned($signed(reg291)) >>> ((reg504 ?
                      (8'ha2) : reg461) ?
                  $unsigned(reg441) : reg345[(3'h4):(2'h2)])))})
            begin
              reg516 <= reg406;
              reg517 <= $unsigned((~((reg472[(3'h7):(3'h6)] >> (reg366 ?
                      reg507 : reg379)) ?
                  reg397 : ($unsigned(reg330) ? (8'h9d) : $signed(reg440)))));
              reg518 = (^~(wire259 && $signed($signed((!reg282)))));
              reg519 = (((+(~&(&(8'ha8)))) ^ (wire259[(5'h16):(4'hd)] << $unsigned($unsigned((7'h44))))) ?
                  reg278[(3'h4):(1'h0)] : reg508);
            end
          else
            begin
              reg518 = $unsigned(reg299[(1'h1):(1'h1)]);
              reg519 = (~|$unsigned($unsigned(((reg374 ? (8'ha5) : reg489) ?
                  reg469[(4'hf):(2'h2)] : $unsigned(reg476)))));
            end
          for (forvar520 = (1'h0); (forvar520 < (2'h3)); forvar520 = (forvar520 + (1'h1)))
            begin
              reg521 = $unsigned((~|reg364[(3'h5):(1'h1)]));
              reg522 = (reg287 + ((($unsigned(wire257) << $signed(reg329)) ?
                  (&(reg444 || reg469)) : forvar513[(1'h1):(1'h0)]) ~^ $unsigned($unsigned((~&reg502)))));
              reg523 = reg325;
              reg524 = reg433[(3'h7):(2'h3)];
              reg525 = ({$unsigned(((reg366 ? reg317 : reg501) ?
                          $signed(reg426) : (reg364 ? reg329 : wire257)))} ?
                  reg310[(3'h5):(1'h0)] : reg494);
            end
          for (forvar526 = (1'h0); (forvar526 < (1'h1)); forvar526 = (forvar526 + (1'h1)))
            begin
              reg527 = $unsigned(reg423);
              reg528 <= reg507;
              reg529 <= reg379;
            end
        end
      else
        begin
          for (forvar516 = (1'h0); (forvar516 < (1'h0)); forvar516 = (forvar516 + (1'h1)))
            begin
              reg518 = reg504[(1'h1):(1'h0)];
              reg519 = (reg406[(4'ha):(4'ha)] >>> reg285);
              reg520 <= (reg385 >= ((reg502[(1'h0):(1'h0)] ?
                  ((reg485 ?
                      reg503 : reg444) || forvar526[(4'h9):(1'h1)]) : (8'hab)) != $unsigned(($signed(reg385) ?
                  $unsigned((8'hb2)) : $signed(reg298)))));
            end
          if (((&$signed($signed((|reg339)))) ?
              ((^~wire259) > (-(reg478[(3'h4):(2'h2)] < $signed(reg334)))) : $unsigned(($signed(reg362) ?
                  reg318 : ((wire257 == reg369) == $signed(reg524))))))
            begin
              reg526 <= $signed($signed($unsigned($unsigned($signed(reg350)))));
              reg528 <= ($unsigned(reg522) ?
                  $unsigned({(~&(|reg285)), reg450}) : reg389[(1'h0):(1'h0)]);
              reg530 = $signed((+$signed(((~reg469) << $unsigned(reg525)))));
              reg531 <= reg334;
              reg532 = $signed(reg273);
            end
          else
            begin
              reg526 <= {$unsigned({$unsigned(reg345)}), reg397};
              reg527 = (((8'had) >>> (!({reg291, reg392} ?
                      (^~reg415) : (-reg379)))) ?
                  ((8'h9e) ?
                      (7'h4a) : ((!reg298) ^ ((~|reg415) ?
                          $unsigned(reg379) : reg524))) : (^($signed(reg363) ?
                      ({(7'h48), forvar513} < (reg505 == reg355)) : reg440)));
              reg528 <= reg318[(1'h0):(1'h0)];
              reg529 <= reg528;
            end
          for (forvar533 = (1'h0); (forvar533 < (1'h0)); forvar533 = (forvar533 + (1'h1)))
            begin
              reg534 = $signed(($signed(((reg350 >= reg522) ^ {reg469,
                      (8'ha7)})) ?
                  reg440 : reg459[(4'hb):(4'h8)]));
              reg535 = $unsigned($signed((((^~reg388) + $unsigned(reg516)) ?
                  ({(8'ha8)} ?
                      (~&reg508) : reg527[(2'h3):(2'h3)]) : ($signed((8'hbd)) < {reg472,
                      reg427}))));
              reg536 <= (((reg463[(4'h9):(4'h9)] ?
                          (8'hbb) : ((reg363 + reg444) * (reg459 ?
                              reg373 : reg269))) ?
                      reg298 : ((-reg459) * ({reg515} ?
                          $signed(wire342) : (8'hac)))) ?
                  (-($signed((wire342 ? reg266 : reg362)) ?
                      ($unsigned(reg450) ?
                          reg405 : $signed(reg496)) : reg278)) : $unsigned(reg330[(1'h0):(1'h0)]));
              reg537 <= ($signed($unsigned(forvar513)) ?
                  reg368[(1'h1):(1'h1)] : reg357[(3'h6):(3'h4)]);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar538 = (1'h0); (forvar538 < (3'h4)); forvar538 = (forvar538 + (1'h1)))
        begin
          reg539 <= $signed((({$unsigned(reg275),
              (reg516 ?
                  (7'h42) : reg418)} && reg420[(2'h2):(2'h2)]) & $signed(reg494[(2'h2):(2'h2)])));
        end
      reg540 = (reg397[(5'h15):(4'hb)] | reg305[(5'h11):(5'h10)]);
    end
  assign wire541 = (7'h43);
  assign wire542 = {reg309};
  always
    @(posedge clk) begin
      if (((~|({{reg478, (8'ha5)}, (8'h9f)} ?
              wire256[(1'h1):(1'h0)] : reg429[(4'h8):(3'h4)])) ?
          reg320[(3'h6):(3'h5)] : $signed((({reg500} ?
              (+(7'h47)) : ((8'hb4) >= reg341)) < (~reg385)))))
        begin
          reg543 <= reg489;
          for (forvar544 = (1'h0); (forvar544 < (2'h2)); forvar544 = (forvar544 + (1'h1)))
            begin
              reg545 <= $unsigned(((($signed((8'hb3)) ?
                      $signed(reg408) : (reg311 ^~ reg330)) ?
                  (-(!reg539)) : $signed((-(7'h49)))) != ((reg289[(2'h3):(2'h3)] + (^reg263)) ?
                  $signed($unsigned(reg315)) : $signed(reg341[(3'h6):(2'h3)]))));
              reg546 <= $unsigned($signed($signed(reg287[(1'h0):(1'h0)])));
              reg547 = $signed(($unsigned((-(8'ha2))) ?
                  ($signed((+reg367)) ?
                      (8'h9c) : reg282[(2'h3):(1'h1)]) : $unsigned(reg368[(1'h1):(1'h0)])));
            end
          for (forvar548 = (1'h0); (forvar548 < (2'h3)); forvar548 = (forvar548 + (1'h1)))
            begin
              reg549 <= $unsigned({reg459[(4'hf):(1'h0)]});
              reg550 = ((reg297[(1'h1):(1'h1)] ?
                      $signed({(reg264 ^ (8'h9d)),
                          ((8'hb7) <<< wire259)}) : reg494[(3'h4):(2'h2)]) ?
                  $unsigned($unsigned(reg269)) : $signed($signed((-(^reg399)))));
              reg551 <= (reg362 <<< (reg441 || $signed($signed((reg317 ?
                  reg528 : reg374)))));
            end
        end
      else
        begin
          reg543 <= $unsigned(reg368[(2'h3):(2'h3)]);
          if ($unsigned((!reg500)))
            begin
              reg544 <= $unsigned(reg269);
            end
          else
            begin
              reg544 <= forvar548;
              reg545 <= ({((((8'hb1) ? reg368 : wire258) ?
                          (-reg292) : $signed(reg313)) ^ reg373),
                      $signed((reg266 ^ (~|(8'ha7))))} ?
                  reg301 : (|(reg356[(3'h7):(3'h7)] && ({reg298} > reg517))));
              reg546 <= reg405;
              reg547 = $unsigned($signed((~&reg547)));
              reg548 = ((~&($unsigned((8'hba)) >>> $unsigned(reg423[(5'h12):(3'h5)]))) || reg429);
            end
          reg549 <= reg334;
        end
      for (forvar552 = (1'h0); (forvar552 < (2'h3)); forvar552 = (forvar552 + (1'h1)))
        begin
          if ({(~^$signed(((reg266 && reg504) || reg325))),
              ({(~^$unsigned((7'h44)))} <<< forvar544[(1'h1):(1'h0)])})
            begin
              reg553 <= $signed((&(8'h9d)));
              reg554 = reg452;
              reg555 = $signed($signed((($signed((8'hb1)) == {reg368, reg454}) ?
                  reg549[(4'hd):(3'h4)] : (7'h46))));
              reg556 = $unsigned(reg420);
              reg557 = wire342[(4'he):(1'h0)];
            end
          else
            begin
              reg553 <= $signed(($unsigned($signed($signed(reg332))) ?
                  reg289 : wire435[(3'h4):(1'h0)]));
            end
          if (((^~reg313[(4'h8):(1'h0)]) ~^ $unsigned($signed($unsigned(reg379[(4'h8):(2'h2)])))))
            begin
              reg558 <= ((!($signed(reg469) == ({reg548, reg537} ?
                      reg307[(2'h3):(2'h2)] : {wire457}))) ?
                  wire256 : (^~(&(~&$unsigned(reg341)))));
              reg559 = ((|reg356[(3'h5):(3'h5)]) ^ (!({(reg299 ~^ reg452),
                      reg472} ?
                  ($signed(reg357) ?
                      ((8'ha4) ? reg325 : wire256) : ((8'had) ?
                          reg332 : wire257)) : ({(8'h9c)} || $unsigned(reg528)))));
              reg560 <= $unsigned(reg290);
              reg561 = (((~&reg263) ?
                  ((^$unsigned((8'hac))) ?
                      ((reg514 ? reg367 : reg560) ?
                          reg389[(1'h0):(1'h0)] : $signed(reg313)) : reg478) : reg392[(2'h3):(1'h1)]) << $unsigned({reg291[(2'h2):(1'h1)],
                  ({reg469, (8'ha2)} ?
                      reg373[(4'hd):(1'h1)] : (reg452 < (8'hbc)))}));
            end
          else
            begin
              reg558 <= (reg543[(3'h4):(1'h1)] ?
                  $signed(({$signed(reg548)} ?
                      ($unsigned((8'hb7)) * reg418) : $signed(((8'h9c) ?
                          reg496 : reg309)))) : (^reg364[(3'h6):(2'h2)]));
            end
          reg562 <= {reg423[(4'ha):(3'h4)]};
          reg563 <= $unsigned((reg514[(1'h1):(1'h1)] ?
              reg463 : {((reg278 ? (8'hb8) : reg408) < ((8'hb3) ?
                      reg561 : reg539)),
                  $signed($signed((7'h4a)))}));
          for (forvar564 = (1'h0); (forvar564 < (2'h2)); forvar564 = (forvar564 + (1'h1)))
            begin
              reg565 <= (~^reg319[(4'ha):(3'h7)]);
              reg566 <= $unsigned(reg537[(5'h15):(4'hb)]);
              reg567 <= (!($unsigned((&$unsigned(reg298))) ^~ $signed($signed($signed((8'h9d))))));
              reg568 = (^(^~$signed(reg501)));
            end
        end
      reg569 <= $unsigned(reg366[(1'h0):(1'h0)]);
      if (reg550[(2'h2):(1'h1)])
        begin
          reg570 <= (^(~&(8'ha5)));
          reg571 = $signed(reg379[(2'h3):(2'h2)]);
        end
      else
        begin
          if (((reg332 ?
                  ((~(reg269 + reg314)) ?
                      (reg415 ?
                          ((8'hb8) < reg374) : $unsigned((8'hac))) : (|(reg282 ~^ reg385))) : reg547[(3'h5):(1'h0)]) ?
              reg320[(1'h1):(1'h0)] : ((&$unsigned({reg339})) >> reg571)))
            begin
              reg570 <= reg500[(1'h0):(1'h0)];
              reg572 <= reg567;
              reg573 <= ($signed((reg543[(4'hb):(3'h5)] ?
                      $signed(reg570[(3'h5):(3'h5)]) : ($unsigned((8'ha5)) >>> reg357[(2'h3):(1'h1)]))) ?
                  ($signed($signed($signed((8'ha0)))) ?
                      $unsigned(($unsigned((8'haa)) || {reg314,
                          reg452})) : reg444[(4'hd):(3'h6)]) : (-$signed(((reg266 * reg389) << (~|wire370)))));
              reg574 <= reg514;
              reg575 = ($signed((forvar552 * $unsigned((reg363 > (7'h4a))))) <<< reg503[(2'h2):(2'h2)]);
            end
          else
            begin
              reg571 = reg319[(1'h1):(1'h0)];
              reg575 = $unsigned(reg549);
              reg576 <= (~reg275);
            end
        end
      for (forvar577 = (1'h0); (forvar577 < (2'h3)); forvar577 = (forvar577 + (1'h1)))
        begin
          if (((reg551 | ({$signed(reg547), (-reg328)} ?
              reg350 : reg566[(3'h4):(2'h2)])) >= reg556[(1'h1):(1'h1)]))
            begin
              reg578 <= reg344;
              reg579 <= $unsigned(reg554[(1'h0):(1'h0)]);
              reg580 = reg356;
            end
          else
            begin
              reg578 <= (wire259 != {(reg450 ?
                      (!$unsigned((8'hbb))) : ((^wire436) <<< (reg406 ?
                          reg463 : reg364))),
                  $unsigned($signed((reg560 * reg441)))});
              reg580 = $signed({reg452});
            end
          for (forvar581 = (1'h0); (forvar581 < (2'h3)); forvar581 = (forvar581 + (1'h1)))
            begin
              reg582 <= reg510;
            end
        end
    end
  assign wire583 = ({reg379} <= (reg320[(1'h0):(1'h0)] ?
                       $unsigned($unsigned($signed(reg389))) : (((reg348 ?
                                   reg266 : reg551) ?
                               {reg450, reg366} : (~^reg367)) ?
                           (~(8'ha5)) : reg416)));
  always
    @(posedge clk) begin
      reg584 <= reg364[(3'h4):(1'h1)];
      if ($unsigned(reg437))
        begin
          reg585 <= {(~|(reg563 ?
                  ($unsigned(reg301) != $unsigned(reg574)) : ($signed(reg287) <= {reg399,
                      (7'h4a)}))),
              reg508[(4'ha):(4'ha)]};
        end
      else
        begin
          if ((^reg313[(2'h3):(2'h3)]))
            begin
              reg585 <= (+reg287);
              reg586 = ((~($signed($unsigned((7'h44))) >> {reg344})) < ($signed((7'h4a)) >= $signed($signed((reg452 ?
                  (8'h9c) : reg531)))));
              reg587 = reg384[(3'h5):(3'h5)];
              reg588 = $unsigned(reg273[(4'h8):(3'h5)]);
              reg589 = $unsigned($unsigned($signed({(reg455 ? reg431 : reg444),
                  reg429})));
            end
          else
            begin
              reg585 <= (reg270[(2'h2):(1'h0)] | reg330[(1'h1):(1'h0)]);
              reg586 = reg569;
            end
          reg590 <= reg409;
        end
    end
  always
    @(posedge clk) begin
      reg591 <= $unsigned((!$signed($unsigned((wire541 | reg415)))));
    end
  always
    @(posedge clk) begin
      reg592 = ($unsigned((~&$signed(((8'haf) ?
          reg289 : reg405)))) & ((^(8'h9e)) ?
          ($unsigned({(8'hb4)}) && $unsigned($unsigned(reg463))) : (8'hbd)));
      if ((+((reg562[(2'h2):(1'h1)] ? (-reg364) : (-reg570)) ?
          (&reg526[(1'h0):(1'h0)]) : $signed(reg309))))
        begin
          reg593 <= ($signed($signed($unsigned((reg469 < reg514)))) + ((wire257 ?
              ($unsigned(reg399) * reg437[(4'h9):(4'h8)]) : (reg299 * reg290)) ^ $signed(($signed(reg309) || $unsigned(reg355)))));
          if (reg569)
            begin
              reg594 = (&reg399);
            end
          else
            begin
              reg594 = ((&($signed((reg341 ? reg508 : reg426)) ?
                  reg426[(1'h0):(1'h0)] : reg305)) <<< $signed($signed(((reg311 ?
                      wire370 : reg366) ?
                  (reg311 ? reg485 : reg291) : (8'hab)))));
              reg595 <= (($unsigned(reg429[(3'h6):(2'h2)]) ?
                      $signed($unsigned(((8'hbf) ?
                          reg501 : reg328))) : (reg563[(3'h5):(3'h4)] ?
                          ($signed(reg544) || (wire542 + reg545)) : ($signed(reg297) < {(8'hb3),
                              reg311}))) ?
                  ({reg319, (|$signed(reg291))} < ($unsigned((!reg441)) ?
                      (&(reg465 ?
                          reg500 : reg270)) : ((reg539 <<< reg339) >>> (reg574 ?
                          reg504 : reg344)))) : $unsigned($signed(reg565[(4'hb):(4'h9)])));
            end
        end
      else
        begin
          for (forvar593 = (1'h0); (forvar593 < (1'h1)); forvar593 = (forvar593 + (1'h1)))
            begin
              reg595 <= ((7'h46) ?
                  (8'h9c) : ((&(~&$unsigned(reg289))) ?
                      ($unsigned($unsigned(reg528)) && $unsigned(reg275)) : reg317));
              reg596 = reg585;
            end
          reg597 = reg405;
          reg598 <= reg318;
          reg599 = $unsigned({($unsigned((reg278 ?
                  wire258 : reg516)) ^ (8'hbc))});
        end
    end
  always
    @(posedge clk) begin
      reg600 <= wire256[(1'h0):(1'h0)];
      reg601 <= (($signed(reg369) ? (&reg408) : (~|reg344[(1'h0):(1'h0)])) ?
          (({(reg562 ^ reg423), (^reg285)} ?
              $signed(reg558[(3'h4):(2'h2)]) : $unsigned(reg551[(4'he):(4'h9)])) && (!reg368)) : {((^reg481[(5'h12):(4'ha)]) ?
                  (8'hae) : $unsigned($unsigned(reg600)))});
      reg602 = $signed({(&((reg494 ? (8'ha9) : (8'h9d)) ?
              $unsigned(reg573) : reg278[(3'h4):(3'h4)])),
          reg399});
      if ((($signed($unsigned(reg601[(5'h12):(4'hb)])) ?
              {(reg385[(3'h5):(3'h4)] <= reg485),
                  $unsigned($unsigned(reg585))} : $signed((!wire435[(3'h6):(2'h3)]))) ?
          (~(({reg317,
              (8'hbb)} ^ $unsigned(reg591)) & (-reg397[(3'h7):(3'h4)]))) : $unsigned($unsigned(reg287[(2'h2):(1'h1)]))))
        begin
          reg603 = (-$signed($signed(($unsigned(reg544) ~^ (^(8'ha0))))));
          if (((+reg328) + reg362[(4'hb):(4'ha)]))
            begin
              reg604 <= {{reg264[(3'h7):(3'h4)]},
                  (!{((reg543 * reg576) == $unsigned((8'haf)))})};
              reg605 = (reg569 + $signed(reg313[(3'h7):(3'h4)]));
              reg606 = $unsigned((7'h40));
              reg607 <= $unsigned(reg431[(1'h0):(1'h0)]);
            end
          else
            begin
              reg604 <= reg565;
              reg607 <= (-$signed((~^(~^(reg558 > reg408)))));
              reg608 = (reg368[(2'h3):(1'h1)] ?
                  $signed(reg408[(1'h0):(1'h0)]) : $signed((8'ha5)));
              reg609 <= reg397[(2'h2):(1'h0)];
              reg610 = (~&$signed($unsigned($signed(reg343))));
            end
          reg611 = (reg301 ?
              $unsigned((~&reg610[(4'h9):(2'h3)])) : $signed(reg314[(4'h9):(4'h8)]));
        end
      else
        begin
          reg604 <= (reg388[(2'h3):(1'h1)] && (~^((^(-reg469)) * (~|(8'ha1)))));
          for (forvar605 = (1'h0); (forvar605 < (1'h0)); forvar605 = (forvar605 + (1'h1)))
            begin
              reg606 = ({reg461,
                  {((reg574 ? reg278 : (8'h9e)) ?
                          (~(7'h4a)) : wire435[(4'h8):(1'h0)])}} != $unsigned(((+(!reg572)) ^ reg300)));
              reg607 <= $unsigned(reg465[(4'hb):(3'h6)]);
            end
          reg608 = $unsigned(reg459);
        end
    end
  assign wire612 = (reg501[(1'h1):(1'h1)] ?
                       {(8'hb1),
                           $signed(reg433[(3'h6):(3'h4)])} : ((reg367[(3'h7):(3'h6)] ?
                               (reg526 ?
                                   reg291[(4'hd):(1'h0)] : $unsigned(reg362)) : (7'h48)) ?
                           $signed(reg339[(3'h6):(3'h5)]) : reg330));
  assign wire613 = (8'haa);
  assign wire614 = reg600[(3'h7):(3'h7)];
endmodule